//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 41
  second input length: 5
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_41_5(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  input [40:0] IN1;
  input [4:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [4:0] P5;
  output [4:0] P6;
  output [4:0] P7;
  output [4:0] P8;
  output [4:0] P9;
  output [4:0] P10;
  output [4:0] P11;
  output [4:0] P12;
  output [4:0] P13;
  output [4:0] P14;
  output [4:0] P15;
  output [4:0] P16;
  output [4:0] P17;
  output [4:0] P18;
  output [4:0] P19;
  output [4:0] P20;
  output [4:0] P21;
  output [4:0] P22;
  output [4:0] P23;
  output [4:0] P24;
  output [4:0] P25;
  output [4:0] P26;
  output [4:0] P27;
  output [4:0] P28;
  output [4:0] P29;
  output [4:0] P30;
  output [4:0] P31;
  output [4:0] P32;
  output [4:0] P33;
  output [4:0] P34;
  output [4:0] P35;
  output [4:0] P36;
  output [4:0] P37;
  output [4:0] P38;
  output [4:0] P39;
  output [4:0] P40;
  output [3:0] P41;
  output [2:0] P42;
  output [1:0] P43;
  output [0:0] P44;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[0] = IN1[1]&IN2[4];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[1] = IN1[2]&IN2[3];
  assign P6[0] = IN1[2]&IN2[4];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[2] = IN1[3]&IN2[2];
  assign P6[1] = IN1[3]&IN2[3];
  assign P7[0] = IN1[3]&IN2[4];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[3] = IN1[4]&IN2[1];
  assign P6[2] = IN1[4]&IN2[2];
  assign P7[1] = IN1[4]&IN2[3];
  assign P8[0] = IN1[4]&IN2[4];
  assign P5[4] = IN1[5]&IN2[0];
  assign P6[3] = IN1[5]&IN2[1];
  assign P7[2] = IN1[5]&IN2[2];
  assign P8[1] = IN1[5]&IN2[3];
  assign P9[0] = IN1[5]&IN2[4];
  assign P6[4] = IN1[6]&IN2[0];
  assign P7[3] = IN1[6]&IN2[1];
  assign P8[2] = IN1[6]&IN2[2];
  assign P9[1] = IN1[6]&IN2[3];
  assign P10[0] = IN1[6]&IN2[4];
  assign P7[4] = IN1[7]&IN2[0];
  assign P8[3] = IN1[7]&IN2[1];
  assign P9[2] = IN1[7]&IN2[2];
  assign P10[1] = IN1[7]&IN2[3];
  assign P11[0] = IN1[7]&IN2[4];
  assign P8[4] = IN1[8]&IN2[0];
  assign P9[3] = IN1[8]&IN2[1];
  assign P10[2] = IN1[8]&IN2[2];
  assign P11[1] = IN1[8]&IN2[3];
  assign P12[0] = IN1[8]&IN2[4];
  assign P9[4] = IN1[9]&IN2[0];
  assign P10[3] = IN1[9]&IN2[1];
  assign P11[2] = IN1[9]&IN2[2];
  assign P12[1] = IN1[9]&IN2[3];
  assign P13[0] = IN1[9]&IN2[4];
  assign P10[4] = IN1[10]&IN2[0];
  assign P11[3] = IN1[10]&IN2[1];
  assign P12[2] = IN1[10]&IN2[2];
  assign P13[1] = IN1[10]&IN2[3];
  assign P14[0] = IN1[10]&IN2[4];
  assign P11[4] = IN1[11]&IN2[0];
  assign P12[3] = IN1[11]&IN2[1];
  assign P13[2] = IN1[11]&IN2[2];
  assign P14[1] = IN1[11]&IN2[3];
  assign P15[0] = IN1[11]&IN2[4];
  assign P12[4] = IN1[12]&IN2[0];
  assign P13[3] = IN1[12]&IN2[1];
  assign P14[2] = IN1[12]&IN2[2];
  assign P15[1] = IN1[12]&IN2[3];
  assign P16[0] = IN1[12]&IN2[4];
  assign P13[4] = IN1[13]&IN2[0];
  assign P14[3] = IN1[13]&IN2[1];
  assign P15[2] = IN1[13]&IN2[2];
  assign P16[1] = IN1[13]&IN2[3];
  assign P17[0] = IN1[13]&IN2[4];
  assign P14[4] = IN1[14]&IN2[0];
  assign P15[3] = IN1[14]&IN2[1];
  assign P16[2] = IN1[14]&IN2[2];
  assign P17[1] = IN1[14]&IN2[3];
  assign P18[0] = IN1[14]&IN2[4];
  assign P15[4] = IN1[15]&IN2[0];
  assign P16[3] = IN1[15]&IN2[1];
  assign P17[2] = IN1[15]&IN2[2];
  assign P18[1] = IN1[15]&IN2[3];
  assign P19[0] = IN1[15]&IN2[4];
  assign P16[4] = IN1[16]&IN2[0];
  assign P17[3] = IN1[16]&IN2[1];
  assign P18[2] = IN1[16]&IN2[2];
  assign P19[1] = IN1[16]&IN2[3];
  assign P20[0] = IN1[16]&IN2[4];
  assign P17[4] = IN1[17]&IN2[0];
  assign P18[3] = IN1[17]&IN2[1];
  assign P19[2] = IN1[17]&IN2[2];
  assign P20[1] = IN1[17]&IN2[3];
  assign P21[0] = IN1[17]&IN2[4];
  assign P18[4] = IN1[18]&IN2[0];
  assign P19[3] = IN1[18]&IN2[1];
  assign P20[2] = IN1[18]&IN2[2];
  assign P21[1] = IN1[18]&IN2[3];
  assign P22[0] = IN1[18]&IN2[4];
  assign P19[4] = IN1[19]&IN2[0];
  assign P20[3] = IN1[19]&IN2[1];
  assign P21[2] = IN1[19]&IN2[2];
  assign P22[1] = IN1[19]&IN2[3];
  assign P23[0] = IN1[19]&IN2[4];
  assign P20[4] = IN1[20]&IN2[0];
  assign P21[3] = IN1[20]&IN2[1];
  assign P22[2] = IN1[20]&IN2[2];
  assign P23[1] = IN1[20]&IN2[3];
  assign P24[0] = IN1[20]&IN2[4];
  assign P21[4] = IN1[21]&IN2[0];
  assign P22[3] = IN1[21]&IN2[1];
  assign P23[2] = IN1[21]&IN2[2];
  assign P24[1] = IN1[21]&IN2[3];
  assign P25[0] = IN1[21]&IN2[4];
  assign P22[4] = IN1[22]&IN2[0];
  assign P23[3] = IN1[22]&IN2[1];
  assign P24[2] = IN1[22]&IN2[2];
  assign P25[1] = IN1[22]&IN2[3];
  assign P26[0] = IN1[22]&IN2[4];
  assign P23[4] = IN1[23]&IN2[0];
  assign P24[3] = IN1[23]&IN2[1];
  assign P25[2] = IN1[23]&IN2[2];
  assign P26[1] = IN1[23]&IN2[3];
  assign P27[0] = IN1[23]&IN2[4];
  assign P24[4] = IN1[24]&IN2[0];
  assign P25[3] = IN1[24]&IN2[1];
  assign P26[2] = IN1[24]&IN2[2];
  assign P27[1] = IN1[24]&IN2[3];
  assign P28[0] = IN1[24]&IN2[4];
  assign P25[4] = IN1[25]&IN2[0];
  assign P26[3] = IN1[25]&IN2[1];
  assign P27[2] = IN1[25]&IN2[2];
  assign P28[1] = IN1[25]&IN2[3];
  assign P29[0] = IN1[25]&IN2[4];
  assign P26[4] = IN1[26]&IN2[0];
  assign P27[3] = IN1[26]&IN2[1];
  assign P28[2] = IN1[26]&IN2[2];
  assign P29[1] = IN1[26]&IN2[3];
  assign P30[0] = IN1[26]&IN2[4];
  assign P27[4] = IN1[27]&IN2[0];
  assign P28[3] = IN1[27]&IN2[1];
  assign P29[2] = IN1[27]&IN2[2];
  assign P30[1] = IN1[27]&IN2[3];
  assign P31[0] = IN1[27]&IN2[4];
  assign P28[4] = IN1[28]&IN2[0];
  assign P29[3] = IN1[28]&IN2[1];
  assign P30[2] = IN1[28]&IN2[2];
  assign P31[1] = IN1[28]&IN2[3];
  assign P32[0] = IN1[28]&IN2[4];
  assign P29[4] = IN1[29]&IN2[0];
  assign P30[3] = IN1[29]&IN2[1];
  assign P31[2] = IN1[29]&IN2[2];
  assign P32[1] = IN1[29]&IN2[3];
  assign P33[0] = IN1[29]&IN2[4];
  assign P30[4] = IN1[30]&IN2[0];
  assign P31[3] = IN1[30]&IN2[1];
  assign P32[2] = IN1[30]&IN2[2];
  assign P33[1] = IN1[30]&IN2[3];
  assign P34[0] = IN1[30]&IN2[4];
  assign P31[4] = IN1[31]&IN2[0];
  assign P32[3] = IN1[31]&IN2[1];
  assign P33[2] = IN1[31]&IN2[2];
  assign P34[1] = IN1[31]&IN2[3];
  assign P35[0] = IN1[31]&IN2[4];
  assign P32[4] = IN1[32]&IN2[0];
  assign P33[3] = IN1[32]&IN2[1];
  assign P34[2] = IN1[32]&IN2[2];
  assign P35[1] = IN1[32]&IN2[3];
  assign P36[0] = IN1[32]&IN2[4];
  assign P33[4] = IN1[33]&IN2[0];
  assign P34[3] = IN1[33]&IN2[1];
  assign P35[2] = IN1[33]&IN2[2];
  assign P36[1] = IN1[33]&IN2[3];
  assign P37[0] = IN1[33]&IN2[4];
  assign P34[4] = IN1[34]&IN2[0];
  assign P35[3] = IN1[34]&IN2[1];
  assign P36[2] = IN1[34]&IN2[2];
  assign P37[1] = IN1[34]&IN2[3];
  assign P38[0] = IN1[34]&IN2[4];
  assign P35[4] = IN1[35]&IN2[0];
  assign P36[3] = IN1[35]&IN2[1];
  assign P37[2] = IN1[35]&IN2[2];
  assign P38[1] = IN1[35]&IN2[3];
  assign P39[0] = IN1[35]&IN2[4];
  assign P36[4] = IN1[36]&IN2[0];
  assign P37[3] = IN1[36]&IN2[1];
  assign P38[2] = IN1[36]&IN2[2];
  assign P39[1] = IN1[36]&IN2[3];
  assign P40[0] = IN1[36]&IN2[4];
  assign P37[4] = IN1[37]&IN2[0];
  assign P38[3] = IN1[37]&IN2[1];
  assign P39[2] = IN1[37]&IN2[2];
  assign P40[1] = IN1[37]&IN2[3];
  assign P41[0] = IN1[37]&IN2[4];
  assign P38[4] = IN1[38]&IN2[0];
  assign P39[3] = IN1[38]&IN2[1];
  assign P40[2] = IN1[38]&IN2[2];
  assign P41[1] = IN1[38]&IN2[3];
  assign P42[0] = IN1[38]&IN2[4];
  assign P39[4] = IN1[39]&IN2[0];
  assign P40[3] = IN1[39]&IN2[1];
  assign P41[2] = IN1[39]&IN2[2];
  assign P42[1] = IN1[39]&IN2[3];
  assign P43[0] = IN1[39]&IN2[4];
  assign P40[4] = IN1[40]&IN2[0];
  assign P41[3] = IN1[40]&IN2[1];
  assign P42[2] = IN1[40]&IN2[2];
  assign P43[1] = IN1[40]&IN2[3];
  assign P44[0] = IN1[40]&IN2[4];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [4:0] IN5;
  input [4:0] IN6;
  input [4:0] IN7;
  input [4:0] IN8;
  input [4:0] IN9;
  input [4:0] IN10;
  input [4:0] IN11;
  input [4:0] IN12;
  input [4:0] IN13;
  input [4:0] IN14;
  input [4:0] IN15;
  input [4:0] IN16;
  input [4:0] IN17;
  input [4:0] IN18;
  input [4:0] IN19;
  input [4:0] IN20;
  input [4:0] IN21;
  input [4:0] IN22;
  input [4:0] IN23;
  input [4:0] IN24;
  input [4:0] IN25;
  input [4:0] IN26;
  input [4:0] IN27;
  input [4:0] IN28;
  input [4:0] IN29;
  input [4:0] IN30;
  input [4:0] IN31;
  input [4:0] IN32;
  input [4:0] IN33;
  input [4:0] IN34;
  input [4:0] IN35;
  input [4:0] IN36;
  input [4:0] IN37;
  input [4:0] IN38;
  input [4:0] IN39;
  input [4:0] IN40;
  input [3:0] IN41;
  input [2:0] IN42;
  input [1:0] IN43;
  input [0:0] IN44;
  output [44:0] Out1;
  output [3:0] Out2;
  wire w206;
  wire w207;
  wire w208;
  wire w209;
  wire w210;
  wire w211;
  wire w212;
  wire w213;
  wire w214;
  wire w215;
  wire w216;
  wire w217;
  wire w218;
  wire w219;
  wire w220;
  wire w221;
  wire w222;
  wire w223;
  wire w224;
  wire w225;
  wire w226;
  wire w227;
  wire w228;
  wire w229;
  wire w230;
  wire w231;
  wire w232;
  wire w233;
  wire w234;
  wire w235;
  wire w236;
  wire w237;
  wire w238;
  wire w239;
  wire w240;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w246;
  wire w247;
  wire w248;
  wire w249;
  wire w250;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w446;
  wire w448;
  wire w450;
  wire w452;
  wire w454;
  wire w456;
  wire w458;
  wire w460;
  wire w462;
  wire w464;
  wire w466;
  wire w468;
  wire w470;
  wire w472;
  wire w474;
  wire w476;
  wire w478;
  wire w480;
  wire w482;
  wire w484;
  wire w486;
  wire w488;
  wire w490;
  wire w492;
  wire w494;
  wire w496;
  wire w498;
  wire w500;
  wire w502;
  wire w504;
  wire w506;
  wire w508;
  wire w510;
  wire w512;
  wire w514;
  wire w516;
  wire w518;
  wire w520;
  wire w522;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w206);
  FullAdder U1 (w206, IN2[0], IN2[1], w207, w208);
  FullAdder U2 (w208, IN3[0], IN3[1], w209, w210);
  FullAdder U3 (w210, IN4[0], IN4[1], w211, w212);
  FullAdder U4 (w212, IN5[0], IN5[1], w213, w214);
  FullAdder U5 (w214, IN6[0], IN6[1], w215, w216);
  FullAdder U6 (w216, IN7[0], IN7[1], w217, w218);
  FullAdder U7 (w218, IN8[0], IN8[1], w219, w220);
  FullAdder U8 (w220, IN9[0], IN9[1], w221, w222);
  FullAdder U9 (w222, IN10[0], IN10[1], w223, w224);
  FullAdder U10 (w224, IN11[0], IN11[1], w225, w226);
  FullAdder U11 (w226, IN12[0], IN12[1], w227, w228);
  FullAdder U12 (w228, IN13[0], IN13[1], w229, w230);
  FullAdder U13 (w230, IN14[0], IN14[1], w231, w232);
  FullAdder U14 (w232, IN15[0], IN15[1], w233, w234);
  FullAdder U15 (w234, IN16[0], IN16[1], w235, w236);
  FullAdder U16 (w236, IN17[0], IN17[1], w237, w238);
  FullAdder U17 (w238, IN18[0], IN18[1], w239, w240);
  FullAdder U18 (w240, IN19[0], IN19[1], w241, w242);
  FullAdder U19 (w242, IN20[0], IN20[1], w243, w244);
  FullAdder U20 (w244, IN21[0], IN21[1], w245, w246);
  FullAdder U21 (w246, IN22[0], IN22[1], w247, w248);
  FullAdder U22 (w248, IN23[0], IN23[1], w249, w250);
  FullAdder U23 (w250, IN24[0], IN24[1], w251, w252);
  FullAdder U24 (w252, IN25[0], IN25[1], w253, w254);
  FullAdder U25 (w254, IN26[0], IN26[1], w255, w256);
  FullAdder U26 (w256, IN27[0], IN27[1], w257, w258);
  FullAdder U27 (w258, IN28[0], IN28[1], w259, w260);
  FullAdder U28 (w260, IN29[0], IN29[1], w261, w262);
  FullAdder U29 (w262, IN30[0], IN30[1], w263, w264);
  FullAdder U30 (w264, IN31[0], IN31[1], w265, w266);
  FullAdder U31 (w266, IN32[0], IN32[1], w267, w268);
  FullAdder U32 (w268, IN33[0], IN33[1], w269, w270);
  FullAdder U33 (w270, IN34[0], IN34[1], w271, w272);
  FullAdder U34 (w272, IN35[0], IN35[1], w273, w274);
  FullAdder U35 (w274, IN36[0], IN36[1], w275, w276);
  FullAdder U36 (w276, IN37[0], IN37[1], w277, w278);
  FullAdder U37 (w278, IN38[0], IN38[1], w279, w280);
  FullAdder U38 (w280, IN39[0], IN39[1], w281, w282);
  FullAdder U39 (w282, IN40[0], IN40[1], w283, w284);
  HalfAdder U40 (w207, IN2[2], Out1[2], w286);
  FullAdder U41 (w286, w209, IN3[2], w287, w288);
  FullAdder U42 (w288, w211, IN4[2], w289, w290);
  FullAdder U43 (w290, w213, IN5[2], w291, w292);
  FullAdder U44 (w292, w215, IN6[2], w293, w294);
  FullAdder U45 (w294, w217, IN7[2], w295, w296);
  FullAdder U46 (w296, w219, IN8[2], w297, w298);
  FullAdder U47 (w298, w221, IN9[2], w299, w300);
  FullAdder U48 (w300, w223, IN10[2], w301, w302);
  FullAdder U49 (w302, w225, IN11[2], w303, w304);
  FullAdder U50 (w304, w227, IN12[2], w305, w306);
  FullAdder U51 (w306, w229, IN13[2], w307, w308);
  FullAdder U52 (w308, w231, IN14[2], w309, w310);
  FullAdder U53 (w310, w233, IN15[2], w311, w312);
  FullAdder U54 (w312, w235, IN16[2], w313, w314);
  FullAdder U55 (w314, w237, IN17[2], w315, w316);
  FullAdder U56 (w316, w239, IN18[2], w317, w318);
  FullAdder U57 (w318, w241, IN19[2], w319, w320);
  FullAdder U58 (w320, w243, IN20[2], w321, w322);
  FullAdder U59 (w322, w245, IN21[2], w323, w324);
  FullAdder U60 (w324, w247, IN22[2], w325, w326);
  FullAdder U61 (w326, w249, IN23[2], w327, w328);
  FullAdder U62 (w328, w251, IN24[2], w329, w330);
  FullAdder U63 (w330, w253, IN25[2], w331, w332);
  FullAdder U64 (w332, w255, IN26[2], w333, w334);
  FullAdder U65 (w334, w257, IN27[2], w335, w336);
  FullAdder U66 (w336, w259, IN28[2], w337, w338);
  FullAdder U67 (w338, w261, IN29[2], w339, w340);
  FullAdder U68 (w340, w263, IN30[2], w341, w342);
  FullAdder U69 (w342, w265, IN31[2], w343, w344);
  FullAdder U70 (w344, w267, IN32[2], w345, w346);
  FullAdder U71 (w346, w269, IN33[2], w347, w348);
  FullAdder U72 (w348, w271, IN34[2], w349, w350);
  FullAdder U73 (w350, w273, IN35[2], w351, w352);
  FullAdder U74 (w352, w275, IN36[2], w353, w354);
  FullAdder U75 (w354, w277, IN37[2], w355, w356);
  FullAdder U76 (w356, w279, IN38[2], w357, w358);
  FullAdder U77 (w358, w281, IN39[2], w359, w360);
  FullAdder U78 (w360, w283, IN40[2], w361, w362);
  FullAdder U79 (w362, w284, IN41[0], w363, w364);
  HalfAdder U80 (w287, IN3[3], Out1[3], w366);
  FullAdder U81 (w366, w289, IN4[3], w367, w368);
  FullAdder U82 (w368, w291, IN5[3], w369, w370);
  FullAdder U83 (w370, w293, IN6[3], w371, w372);
  FullAdder U84 (w372, w295, IN7[3], w373, w374);
  FullAdder U85 (w374, w297, IN8[3], w375, w376);
  FullAdder U86 (w376, w299, IN9[3], w377, w378);
  FullAdder U87 (w378, w301, IN10[3], w379, w380);
  FullAdder U88 (w380, w303, IN11[3], w381, w382);
  FullAdder U89 (w382, w305, IN12[3], w383, w384);
  FullAdder U90 (w384, w307, IN13[3], w385, w386);
  FullAdder U91 (w386, w309, IN14[3], w387, w388);
  FullAdder U92 (w388, w311, IN15[3], w389, w390);
  FullAdder U93 (w390, w313, IN16[3], w391, w392);
  FullAdder U94 (w392, w315, IN17[3], w393, w394);
  FullAdder U95 (w394, w317, IN18[3], w395, w396);
  FullAdder U96 (w396, w319, IN19[3], w397, w398);
  FullAdder U97 (w398, w321, IN20[3], w399, w400);
  FullAdder U98 (w400, w323, IN21[3], w401, w402);
  FullAdder U99 (w402, w325, IN22[3], w403, w404);
  FullAdder U100 (w404, w327, IN23[3], w405, w406);
  FullAdder U101 (w406, w329, IN24[3], w407, w408);
  FullAdder U102 (w408, w331, IN25[3], w409, w410);
  FullAdder U103 (w410, w333, IN26[3], w411, w412);
  FullAdder U104 (w412, w335, IN27[3], w413, w414);
  FullAdder U105 (w414, w337, IN28[3], w415, w416);
  FullAdder U106 (w416, w339, IN29[3], w417, w418);
  FullAdder U107 (w418, w341, IN30[3], w419, w420);
  FullAdder U108 (w420, w343, IN31[3], w421, w422);
  FullAdder U109 (w422, w345, IN32[3], w423, w424);
  FullAdder U110 (w424, w347, IN33[3], w425, w426);
  FullAdder U111 (w426, w349, IN34[3], w427, w428);
  FullAdder U112 (w428, w351, IN35[3], w429, w430);
  FullAdder U113 (w430, w353, IN36[3], w431, w432);
  FullAdder U114 (w432, w355, IN37[3], w433, w434);
  FullAdder U115 (w434, w357, IN38[3], w435, w436);
  FullAdder U116 (w436, w359, IN39[3], w437, w438);
  FullAdder U117 (w438, w361, IN40[3], w439, w440);
  FullAdder U118 (w440, w363, IN41[1], w441, w442);
  FullAdder U119 (w442, w364, IN42[0], w443, w444);
  HalfAdder U120 (w367, IN4[4], Out1[4], w446);
  FullAdder U121 (w446, w369, IN5[4], Out1[5], w448);
  FullAdder U122 (w448, w371, IN6[4], Out1[6], w450);
  FullAdder U123 (w450, w373, IN7[4], Out1[7], w452);
  FullAdder U124 (w452, w375, IN8[4], Out1[8], w454);
  FullAdder U125 (w454, w377, IN9[4], Out1[9], w456);
  FullAdder U126 (w456, w379, IN10[4], Out1[10], w458);
  FullAdder U127 (w458, w381, IN11[4], Out1[11], w460);
  FullAdder U128 (w460, w383, IN12[4], Out1[12], w462);
  FullAdder U129 (w462, w385, IN13[4], Out1[13], w464);
  FullAdder U130 (w464, w387, IN14[4], Out1[14], w466);
  FullAdder U131 (w466, w389, IN15[4], Out1[15], w468);
  FullAdder U132 (w468, w391, IN16[4], Out1[16], w470);
  FullAdder U133 (w470, w393, IN17[4], Out1[17], w472);
  FullAdder U134 (w472, w395, IN18[4], Out1[18], w474);
  FullAdder U135 (w474, w397, IN19[4], Out1[19], w476);
  FullAdder U136 (w476, w399, IN20[4], Out1[20], w478);
  FullAdder U137 (w478, w401, IN21[4], Out1[21], w480);
  FullAdder U138 (w480, w403, IN22[4], Out1[22], w482);
  FullAdder U139 (w482, w405, IN23[4], Out1[23], w484);
  FullAdder U140 (w484, w407, IN24[4], Out1[24], w486);
  FullAdder U141 (w486, w409, IN25[4], Out1[25], w488);
  FullAdder U142 (w488, w411, IN26[4], Out1[26], w490);
  FullAdder U143 (w490, w413, IN27[4], Out1[27], w492);
  FullAdder U144 (w492, w415, IN28[4], Out1[28], w494);
  FullAdder U145 (w494, w417, IN29[4], Out1[29], w496);
  FullAdder U146 (w496, w419, IN30[4], Out1[30], w498);
  FullAdder U147 (w498, w421, IN31[4], Out1[31], w500);
  FullAdder U148 (w500, w423, IN32[4], Out1[32], w502);
  FullAdder U149 (w502, w425, IN33[4], Out1[33], w504);
  FullAdder U150 (w504, w427, IN34[4], Out1[34], w506);
  FullAdder U151 (w506, w429, IN35[4], Out1[35], w508);
  FullAdder U152 (w508, w431, IN36[4], Out1[36], w510);
  FullAdder U153 (w510, w433, IN37[4], Out1[37], w512);
  FullAdder U154 (w512, w435, IN38[4], Out1[38], w514);
  FullAdder U155 (w514, w437, IN39[4], Out1[39], w516);
  FullAdder U156 (w516, w439, IN40[4], Out1[40], w518);
  FullAdder U157 (w518, w441, IN41[2], Out1[41], w520);
  FullAdder U158 (w520, w443, IN42[1], Out1[42], w522);
  FullAdder U159 (w522, w444, IN43[0], Out1[43], Out1[44]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN41[3];
  assign Out2[1] = IN42[2];
  assign Out2[2] = IN43[1];
  assign Out2[3] = IN44[0];

endmodule
module RC_4_4(IN1, IN2, Out);
  input [3:0] IN1;
  input [3:0] IN2;
  output [4:0] Out;
  wire w9;
  wire w11;
  wire w13;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w9);
  FullAdder U1 (IN1[1], IN2[1], w9, Out[1], w11);
  FullAdder U2 (IN1[2], IN2[2], w11, Out[2], w13);
  FullAdder U3 (IN1[3], IN2[3], w13, Out[3], Out[4]);

endmodule
module NR_41_5(IN1, IN2, Out);
  input [40:0] IN1;
  input [4:0] IN2;
  output [45:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [4:0] P5;
  wire [4:0] P6;
  wire [4:0] P7;
  wire [4:0] P8;
  wire [4:0] P9;
  wire [4:0] P10;
  wire [4:0] P11;
  wire [4:0] P12;
  wire [4:0] P13;
  wire [4:0] P14;
  wire [4:0] P15;
  wire [4:0] P16;
  wire [4:0] P17;
  wire [4:0] P18;
  wire [4:0] P19;
  wire [4:0] P20;
  wire [4:0] P21;
  wire [4:0] P22;
  wire [4:0] P23;
  wire [4:0] P24;
  wire [4:0] P25;
  wire [4:0] P26;
  wire [4:0] P27;
  wire [4:0] P28;
  wire [4:0] P29;
  wire [4:0] P30;
  wire [4:0] P31;
  wire [4:0] P32;
  wire [4:0] P33;
  wire [4:0] P34;
  wire [4:0] P35;
  wire [4:0] P36;
  wire [4:0] P37;
  wire [4:0] P38;
  wire [4:0] P39;
  wire [4:0] P40;
  wire [3:0] P41;
  wire [2:0] P42;
  wire [1:0] P43;
  wire [0:0] P44;
  wire [44:0] R1;
  wire [3:0] R2;
  wire [45:0] aOut;
  U_SP_41_5 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, R1, R2);
  RC_4_4 S2 (R1[44:41], R2, aOut[45:41]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign Out = aOut[45:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
