//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 57
  second input length: 7
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_57_7(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  input [56:0] IN1;
  input [6:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [6:0] P37;
  output [6:0] P38;
  output [6:0] P39;
  output [6:0] P40;
  output [6:0] P41;
  output [6:0] P42;
  output [6:0] P43;
  output [6:0] P44;
  output [6:0] P45;
  output [6:0] P46;
  output [6:0] P47;
  output [6:0] P48;
  output [6:0] P49;
  output [6:0] P50;
  output [6:0] P51;
  output [6:0] P52;
  output [6:0] P53;
  output [6:0] P54;
  output [6:0] P55;
  output [6:0] P56;
  output [5:0] P57;
  output [4:0] P58;
  output [3:0] P59;
  output [2:0] P60;
  output [1:0] P61;
  output [0:0] P62;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[0] = IN1[1]&IN2[6];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[1] = IN1[2]&IN2[5];
  assign P8[0] = IN1[2]&IN2[6];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[2] = IN1[3]&IN2[4];
  assign P8[1] = IN1[3]&IN2[5];
  assign P9[0] = IN1[3]&IN2[6];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[3] = IN1[4]&IN2[3];
  assign P8[2] = IN1[4]&IN2[4];
  assign P9[1] = IN1[4]&IN2[5];
  assign P10[0] = IN1[4]&IN2[6];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[4] = IN1[5]&IN2[2];
  assign P8[3] = IN1[5]&IN2[3];
  assign P9[2] = IN1[5]&IN2[4];
  assign P10[1] = IN1[5]&IN2[5];
  assign P11[0] = IN1[5]&IN2[6];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[5] = IN1[6]&IN2[1];
  assign P8[4] = IN1[6]&IN2[2];
  assign P9[3] = IN1[6]&IN2[3];
  assign P10[2] = IN1[6]&IN2[4];
  assign P11[1] = IN1[6]&IN2[5];
  assign P12[0] = IN1[6]&IN2[6];
  assign P7[6] = IN1[7]&IN2[0];
  assign P8[5] = IN1[7]&IN2[1];
  assign P9[4] = IN1[7]&IN2[2];
  assign P10[3] = IN1[7]&IN2[3];
  assign P11[2] = IN1[7]&IN2[4];
  assign P12[1] = IN1[7]&IN2[5];
  assign P13[0] = IN1[7]&IN2[6];
  assign P8[6] = IN1[8]&IN2[0];
  assign P9[5] = IN1[8]&IN2[1];
  assign P10[4] = IN1[8]&IN2[2];
  assign P11[3] = IN1[8]&IN2[3];
  assign P12[2] = IN1[8]&IN2[4];
  assign P13[1] = IN1[8]&IN2[5];
  assign P14[0] = IN1[8]&IN2[6];
  assign P9[6] = IN1[9]&IN2[0];
  assign P10[5] = IN1[9]&IN2[1];
  assign P11[4] = IN1[9]&IN2[2];
  assign P12[3] = IN1[9]&IN2[3];
  assign P13[2] = IN1[9]&IN2[4];
  assign P14[1] = IN1[9]&IN2[5];
  assign P15[0] = IN1[9]&IN2[6];
  assign P10[6] = IN1[10]&IN2[0];
  assign P11[5] = IN1[10]&IN2[1];
  assign P12[4] = IN1[10]&IN2[2];
  assign P13[3] = IN1[10]&IN2[3];
  assign P14[2] = IN1[10]&IN2[4];
  assign P15[1] = IN1[10]&IN2[5];
  assign P16[0] = IN1[10]&IN2[6];
  assign P11[6] = IN1[11]&IN2[0];
  assign P12[5] = IN1[11]&IN2[1];
  assign P13[4] = IN1[11]&IN2[2];
  assign P14[3] = IN1[11]&IN2[3];
  assign P15[2] = IN1[11]&IN2[4];
  assign P16[1] = IN1[11]&IN2[5];
  assign P17[0] = IN1[11]&IN2[6];
  assign P12[6] = IN1[12]&IN2[0];
  assign P13[5] = IN1[12]&IN2[1];
  assign P14[4] = IN1[12]&IN2[2];
  assign P15[3] = IN1[12]&IN2[3];
  assign P16[2] = IN1[12]&IN2[4];
  assign P17[1] = IN1[12]&IN2[5];
  assign P18[0] = IN1[12]&IN2[6];
  assign P13[6] = IN1[13]&IN2[0];
  assign P14[5] = IN1[13]&IN2[1];
  assign P15[4] = IN1[13]&IN2[2];
  assign P16[3] = IN1[13]&IN2[3];
  assign P17[2] = IN1[13]&IN2[4];
  assign P18[1] = IN1[13]&IN2[5];
  assign P19[0] = IN1[13]&IN2[6];
  assign P14[6] = IN1[14]&IN2[0];
  assign P15[5] = IN1[14]&IN2[1];
  assign P16[4] = IN1[14]&IN2[2];
  assign P17[3] = IN1[14]&IN2[3];
  assign P18[2] = IN1[14]&IN2[4];
  assign P19[1] = IN1[14]&IN2[5];
  assign P20[0] = IN1[14]&IN2[6];
  assign P15[6] = IN1[15]&IN2[0];
  assign P16[5] = IN1[15]&IN2[1];
  assign P17[4] = IN1[15]&IN2[2];
  assign P18[3] = IN1[15]&IN2[3];
  assign P19[2] = IN1[15]&IN2[4];
  assign P20[1] = IN1[15]&IN2[5];
  assign P21[0] = IN1[15]&IN2[6];
  assign P16[6] = IN1[16]&IN2[0];
  assign P17[5] = IN1[16]&IN2[1];
  assign P18[4] = IN1[16]&IN2[2];
  assign P19[3] = IN1[16]&IN2[3];
  assign P20[2] = IN1[16]&IN2[4];
  assign P21[1] = IN1[16]&IN2[5];
  assign P22[0] = IN1[16]&IN2[6];
  assign P17[6] = IN1[17]&IN2[0];
  assign P18[5] = IN1[17]&IN2[1];
  assign P19[4] = IN1[17]&IN2[2];
  assign P20[3] = IN1[17]&IN2[3];
  assign P21[2] = IN1[17]&IN2[4];
  assign P22[1] = IN1[17]&IN2[5];
  assign P23[0] = IN1[17]&IN2[6];
  assign P18[6] = IN1[18]&IN2[0];
  assign P19[5] = IN1[18]&IN2[1];
  assign P20[4] = IN1[18]&IN2[2];
  assign P21[3] = IN1[18]&IN2[3];
  assign P22[2] = IN1[18]&IN2[4];
  assign P23[1] = IN1[18]&IN2[5];
  assign P24[0] = IN1[18]&IN2[6];
  assign P19[6] = IN1[19]&IN2[0];
  assign P20[5] = IN1[19]&IN2[1];
  assign P21[4] = IN1[19]&IN2[2];
  assign P22[3] = IN1[19]&IN2[3];
  assign P23[2] = IN1[19]&IN2[4];
  assign P24[1] = IN1[19]&IN2[5];
  assign P25[0] = IN1[19]&IN2[6];
  assign P20[6] = IN1[20]&IN2[0];
  assign P21[5] = IN1[20]&IN2[1];
  assign P22[4] = IN1[20]&IN2[2];
  assign P23[3] = IN1[20]&IN2[3];
  assign P24[2] = IN1[20]&IN2[4];
  assign P25[1] = IN1[20]&IN2[5];
  assign P26[0] = IN1[20]&IN2[6];
  assign P21[6] = IN1[21]&IN2[0];
  assign P22[5] = IN1[21]&IN2[1];
  assign P23[4] = IN1[21]&IN2[2];
  assign P24[3] = IN1[21]&IN2[3];
  assign P25[2] = IN1[21]&IN2[4];
  assign P26[1] = IN1[21]&IN2[5];
  assign P27[0] = IN1[21]&IN2[6];
  assign P22[6] = IN1[22]&IN2[0];
  assign P23[5] = IN1[22]&IN2[1];
  assign P24[4] = IN1[22]&IN2[2];
  assign P25[3] = IN1[22]&IN2[3];
  assign P26[2] = IN1[22]&IN2[4];
  assign P27[1] = IN1[22]&IN2[5];
  assign P28[0] = IN1[22]&IN2[6];
  assign P23[6] = IN1[23]&IN2[0];
  assign P24[5] = IN1[23]&IN2[1];
  assign P25[4] = IN1[23]&IN2[2];
  assign P26[3] = IN1[23]&IN2[3];
  assign P27[2] = IN1[23]&IN2[4];
  assign P28[1] = IN1[23]&IN2[5];
  assign P29[0] = IN1[23]&IN2[6];
  assign P24[6] = IN1[24]&IN2[0];
  assign P25[5] = IN1[24]&IN2[1];
  assign P26[4] = IN1[24]&IN2[2];
  assign P27[3] = IN1[24]&IN2[3];
  assign P28[2] = IN1[24]&IN2[4];
  assign P29[1] = IN1[24]&IN2[5];
  assign P30[0] = IN1[24]&IN2[6];
  assign P25[6] = IN1[25]&IN2[0];
  assign P26[5] = IN1[25]&IN2[1];
  assign P27[4] = IN1[25]&IN2[2];
  assign P28[3] = IN1[25]&IN2[3];
  assign P29[2] = IN1[25]&IN2[4];
  assign P30[1] = IN1[25]&IN2[5];
  assign P31[0] = IN1[25]&IN2[6];
  assign P26[6] = IN1[26]&IN2[0];
  assign P27[5] = IN1[26]&IN2[1];
  assign P28[4] = IN1[26]&IN2[2];
  assign P29[3] = IN1[26]&IN2[3];
  assign P30[2] = IN1[26]&IN2[4];
  assign P31[1] = IN1[26]&IN2[5];
  assign P32[0] = IN1[26]&IN2[6];
  assign P27[6] = IN1[27]&IN2[0];
  assign P28[5] = IN1[27]&IN2[1];
  assign P29[4] = IN1[27]&IN2[2];
  assign P30[3] = IN1[27]&IN2[3];
  assign P31[2] = IN1[27]&IN2[4];
  assign P32[1] = IN1[27]&IN2[5];
  assign P33[0] = IN1[27]&IN2[6];
  assign P28[6] = IN1[28]&IN2[0];
  assign P29[5] = IN1[28]&IN2[1];
  assign P30[4] = IN1[28]&IN2[2];
  assign P31[3] = IN1[28]&IN2[3];
  assign P32[2] = IN1[28]&IN2[4];
  assign P33[1] = IN1[28]&IN2[5];
  assign P34[0] = IN1[28]&IN2[6];
  assign P29[6] = IN1[29]&IN2[0];
  assign P30[5] = IN1[29]&IN2[1];
  assign P31[4] = IN1[29]&IN2[2];
  assign P32[3] = IN1[29]&IN2[3];
  assign P33[2] = IN1[29]&IN2[4];
  assign P34[1] = IN1[29]&IN2[5];
  assign P35[0] = IN1[29]&IN2[6];
  assign P30[6] = IN1[30]&IN2[0];
  assign P31[5] = IN1[30]&IN2[1];
  assign P32[4] = IN1[30]&IN2[2];
  assign P33[3] = IN1[30]&IN2[3];
  assign P34[2] = IN1[30]&IN2[4];
  assign P35[1] = IN1[30]&IN2[5];
  assign P36[0] = IN1[30]&IN2[6];
  assign P31[6] = IN1[31]&IN2[0];
  assign P32[5] = IN1[31]&IN2[1];
  assign P33[4] = IN1[31]&IN2[2];
  assign P34[3] = IN1[31]&IN2[3];
  assign P35[2] = IN1[31]&IN2[4];
  assign P36[1] = IN1[31]&IN2[5];
  assign P37[0] = IN1[31]&IN2[6];
  assign P32[6] = IN1[32]&IN2[0];
  assign P33[5] = IN1[32]&IN2[1];
  assign P34[4] = IN1[32]&IN2[2];
  assign P35[3] = IN1[32]&IN2[3];
  assign P36[2] = IN1[32]&IN2[4];
  assign P37[1] = IN1[32]&IN2[5];
  assign P38[0] = IN1[32]&IN2[6];
  assign P33[6] = IN1[33]&IN2[0];
  assign P34[5] = IN1[33]&IN2[1];
  assign P35[4] = IN1[33]&IN2[2];
  assign P36[3] = IN1[33]&IN2[3];
  assign P37[2] = IN1[33]&IN2[4];
  assign P38[1] = IN1[33]&IN2[5];
  assign P39[0] = IN1[33]&IN2[6];
  assign P34[6] = IN1[34]&IN2[0];
  assign P35[5] = IN1[34]&IN2[1];
  assign P36[4] = IN1[34]&IN2[2];
  assign P37[3] = IN1[34]&IN2[3];
  assign P38[2] = IN1[34]&IN2[4];
  assign P39[1] = IN1[34]&IN2[5];
  assign P40[0] = IN1[34]&IN2[6];
  assign P35[6] = IN1[35]&IN2[0];
  assign P36[5] = IN1[35]&IN2[1];
  assign P37[4] = IN1[35]&IN2[2];
  assign P38[3] = IN1[35]&IN2[3];
  assign P39[2] = IN1[35]&IN2[4];
  assign P40[1] = IN1[35]&IN2[5];
  assign P41[0] = IN1[35]&IN2[6];
  assign P36[6] = IN1[36]&IN2[0];
  assign P37[5] = IN1[36]&IN2[1];
  assign P38[4] = IN1[36]&IN2[2];
  assign P39[3] = IN1[36]&IN2[3];
  assign P40[2] = IN1[36]&IN2[4];
  assign P41[1] = IN1[36]&IN2[5];
  assign P42[0] = IN1[36]&IN2[6];
  assign P37[6] = IN1[37]&IN2[0];
  assign P38[5] = IN1[37]&IN2[1];
  assign P39[4] = IN1[37]&IN2[2];
  assign P40[3] = IN1[37]&IN2[3];
  assign P41[2] = IN1[37]&IN2[4];
  assign P42[1] = IN1[37]&IN2[5];
  assign P43[0] = IN1[37]&IN2[6];
  assign P38[6] = IN1[38]&IN2[0];
  assign P39[5] = IN1[38]&IN2[1];
  assign P40[4] = IN1[38]&IN2[2];
  assign P41[3] = IN1[38]&IN2[3];
  assign P42[2] = IN1[38]&IN2[4];
  assign P43[1] = IN1[38]&IN2[5];
  assign P44[0] = IN1[38]&IN2[6];
  assign P39[6] = IN1[39]&IN2[0];
  assign P40[5] = IN1[39]&IN2[1];
  assign P41[4] = IN1[39]&IN2[2];
  assign P42[3] = IN1[39]&IN2[3];
  assign P43[2] = IN1[39]&IN2[4];
  assign P44[1] = IN1[39]&IN2[5];
  assign P45[0] = IN1[39]&IN2[6];
  assign P40[6] = IN1[40]&IN2[0];
  assign P41[5] = IN1[40]&IN2[1];
  assign P42[4] = IN1[40]&IN2[2];
  assign P43[3] = IN1[40]&IN2[3];
  assign P44[2] = IN1[40]&IN2[4];
  assign P45[1] = IN1[40]&IN2[5];
  assign P46[0] = IN1[40]&IN2[6];
  assign P41[6] = IN1[41]&IN2[0];
  assign P42[5] = IN1[41]&IN2[1];
  assign P43[4] = IN1[41]&IN2[2];
  assign P44[3] = IN1[41]&IN2[3];
  assign P45[2] = IN1[41]&IN2[4];
  assign P46[1] = IN1[41]&IN2[5];
  assign P47[0] = IN1[41]&IN2[6];
  assign P42[6] = IN1[42]&IN2[0];
  assign P43[5] = IN1[42]&IN2[1];
  assign P44[4] = IN1[42]&IN2[2];
  assign P45[3] = IN1[42]&IN2[3];
  assign P46[2] = IN1[42]&IN2[4];
  assign P47[1] = IN1[42]&IN2[5];
  assign P48[0] = IN1[42]&IN2[6];
  assign P43[6] = IN1[43]&IN2[0];
  assign P44[5] = IN1[43]&IN2[1];
  assign P45[4] = IN1[43]&IN2[2];
  assign P46[3] = IN1[43]&IN2[3];
  assign P47[2] = IN1[43]&IN2[4];
  assign P48[1] = IN1[43]&IN2[5];
  assign P49[0] = IN1[43]&IN2[6];
  assign P44[6] = IN1[44]&IN2[0];
  assign P45[5] = IN1[44]&IN2[1];
  assign P46[4] = IN1[44]&IN2[2];
  assign P47[3] = IN1[44]&IN2[3];
  assign P48[2] = IN1[44]&IN2[4];
  assign P49[1] = IN1[44]&IN2[5];
  assign P50[0] = IN1[44]&IN2[6];
  assign P45[6] = IN1[45]&IN2[0];
  assign P46[5] = IN1[45]&IN2[1];
  assign P47[4] = IN1[45]&IN2[2];
  assign P48[3] = IN1[45]&IN2[3];
  assign P49[2] = IN1[45]&IN2[4];
  assign P50[1] = IN1[45]&IN2[5];
  assign P51[0] = IN1[45]&IN2[6];
  assign P46[6] = IN1[46]&IN2[0];
  assign P47[5] = IN1[46]&IN2[1];
  assign P48[4] = IN1[46]&IN2[2];
  assign P49[3] = IN1[46]&IN2[3];
  assign P50[2] = IN1[46]&IN2[4];
  assign P51[1] = IN1[46]&IN2[5];
  assign P52[0] = IN1[46]&IN2[6];
  assign P47[6] = IN1[47]&IN2[0];
  assign P48[5] = IN1[47]&IN2[1];
  assign P49[4] = IN1[47]&IN2[2];
  assign P50[3] = IN1[47]&IN2[3];
  assign P51[2] = IN1[47]&IN2[4];
  assign P52[1] = IN1[47]&IN2[5];
  assign P53[0] = IN1[47]&IN2[6];
  assign P48[6] = IN1[48]&IN2[0];
  assign P49[5] = IN1[48]&IN2[1];
  assign P50[4] = IN1[48]&IN2[2];
  assign P51[3] = IN1[48]&IN2[3];
  assign P52[2] = IN1[48]&IN2[4];
  assign P53[1] = IN1[48]&IN2[5];
  assign P54[0] = IN1[48]&IN2[6];
  assign P49[6] = IN1[49]&IN2[0];
  assign P50[5] = IN1[49]&IN2[1];
  assign P51[4] = IN1[49]&IN2[2];
  assign P52[3] = IN1[49]&IN2[3];
  assign P53[2] = IN1[49]&IN2[4];
  assign P54[1] = IN1[49]&IN2[5];
  assign P55[0] = IN1[49]&IN2[6];
  assign P50[6] = IN1[50]&IN2[0];
  assign P51[5] = IN1[50]&IN2[1];
  assign P52[4] = IN1[50]&IN2[2];
  assign P53[3] = IN1[50]&IN2[3];
  assign P54[2] = IN1[50]&IN2[4];
  assign P55[1] = IN1[50]&IN2[5];
  assign P56[0] = IN1[50]&IN2[6];
  assign P51[6] = IN1[51]&IN2[0];
  assign P52[5] = IN1[51]&IN2[1];
  assign P53[4] = IN1[51]&IN2[2];
  assign P54[3] = IN1[51]&IN2[3];
  assign P55[2] = IN1[51]&IN2[4];
  assign P56[1] = IN1[51]&IN2[5];
  assign P57[0] = IN1[51]&IN2[6];
  assign P52[6] = IN1[52]&IN2[0];
  assign P53[5] = IN1[52]&IN2[1];
  assign P54[4] = IN1[52]&IN2[2];
  assign P55[3] = IN1[52]&IN2[3];
  assign P56[2] = IN1[52]&IN2[4];
  assign P57[1] = IN1[52]&IN2[5];
  assign P58[0] = IN1[52]&IN2[6];
  assign P53[6] = IN1[53]&IN2[0];
  assign P54[5] = IN1[53]&IN2[1];
  assign P55[4] = IN1[53]&IN2[2];
  assign P56[3] = IN1[53]&IN2[3];
  assign P57[2] = IN1[53]&IN2[4];
  assign P58[1] = IN1[53]&IN2[5];
  assign P59[0] = IN1[53]&IN2[6];
  assign P54[6] = IN1[54]&IN2[0];
  assign P55[5] = IN1[54]&IN2[1];
  assign P56[4] = IN1[54]&IN2[2];
  assign P57[3] = IN1[54]&IN2[3];
  assign P58[2] = IN1[54]&IN2[4];
  assign P59[1] = IN1[54]&IN2[5];
  assign P60[0] = IN1[54]&IN2[6];
  assign P55[6] = IN1[55]&IN2[0];
  assign P56[5] = IN1[55]&IN2[1];
  assign P57[4] = IN1[55]&IN2[2];
  assign P58[3] = IN1[55]&IN2[3];
  assign P59[2] = IN1[55]&IN2[4];
  assign P60[1] = IN1[55]&IN2[5];
  assign P61[0] = IN1[55]&IN2[6];
  assign P56[6] = IN1[56]&IN2[0];
  assign P57[5] = IN1[56]&IN2[1];
  assign P58[4] = IN1[56]&IN2[2];
  assign P59[3] = IN1[56]&IN2[3];
  assign P60[2] = IN1[56]&IN2[4];
  assign P61[1] = IN1[56]&IN2[5];
  assign P62[0] = IN1[56]&IN2[6];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [6:0] IN37;
  input [6:0] IN38;
  input [6:0] IN39;
  input [6:0] IN40;
  input [6:0] IN41;
  input [6:0] IN42;
  input [6:0] IN43;
  input [6:0] IN44;
  input [6:0] IN45;
  input [6:0] IN46;
  input [6:0] IN47;
  input [6:0] IN48;
  input [6:0] IN49;
  input [6:0] IN50;
  input [6:0] IN51;
  input [6:0] IN52;
  input [6:0] IN53;
  input [6:0] IN54;
  input [6:0] IN55;
  input [6:0] IN56;
  input [5:0] IN57;
  input [4:0] IN58;
  input [3:0] IN59;
  input [2:0] IN60;
  input [1:0] IN61;
  input [0:0] IN62;
  output [62:0] Out1;
  output [5:0] Out2;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w960;
  wire w962;
  wire w964;
  wire w966;
  wire w968;
  wire w970;
  wire w972;
  wire w974;
  wire w976;
  wire w978;
  wire w980;
  wire w982;
  wire w984;
  wire w986;
  wire w988;
  wire w990;
  wire w992;
  wire w994;
  wire w996;
  wire w998;
  wire w1000;
  wire w1002;
  wire w1004;
  wire w1006;
  wire w1008;
  wire w1010;
  wire w1012;
  wire w1014;
  wire w1016;
  wire w1018;
  wire w1020;
  wire w1022;
  wire w1024;
  wire w1026;
  wire w1028;
  wire w1030;
  wire w1032;
  wire w1034;
  wire w1036;
  wire w1038;
  wire w1040;
  wire w1042;
  wire w1044;
  wire w1046;
  wire w1048;
  wire w1050;
  wire w1052;
  wire w1054;
  wire w1056;
  wire w1058;
  wire w1060;
  wire w1062;
  wire w1064;
  wire w1066;
  wire w1068;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w400);
  FullAdder U1 (w400, IN2[0], IN2[1], w401, w402);
  FullAdder U2 (w402, IN3[0], IN3[1], w403, w404);
  FullAdder U3 (w404, IN4[0], IN4[1], w405, w406);
  FullAdder U4 (w406, IN5[0], IN5[1], w407, w408);
  FullAdder U5 (w408, IN6[0], IN6[1], w409, w410);
  FullAdder U6 (w410, IN7[0], IN7[1], w411, w412);
  FullAdder U7 (w412, IN8[0], IN8[1], w413, w414);
  FullAdder U8 (w414, IN9[0], IN9[1], w415, w416);
  FullAdder U9 (w416, IN10[0], IN10[1], w417, w418);
  FullAdder U10 (w418, IN11[0], IN11[1], w419, w420);
  FullAdder U11 (w420, IN12[0], IN12[1], w421, w422);
  FullAdder U12 (w422, IN13[0], IN13[1], w423, w424);
  FullAdder U13 (w424, IN14[0], IN14[1], w425, w426);
  FullAdder U14 (w426, IN15[0], IN15[1], w427, w428);
  FullAdder U15 (w428, IN16[0], IN16[1], w429, w430);
  FullAdder U16 (w430, IN17[0], IN17[1], w431, w432);
  FullAdder U17 (w432, IN18[0], IN18[1], w433, w434);
  FullAdder U18 (w434, IN19[0], IN19[1], w435, w436);
  FullAdder U19 (w436, IN20[0], IN20[1], w437, w438);
  FullAdder U20 (w438, IN21[0], IN21[1], w439, w440);
  FullAdder U21 (w440, IN22[0], IN22[1], w441, w442);
  FullAdder U22 (w442, IN23[0], IN23[1], w443, w444);
  FullAdder U23 (w444, IN24[0], IN24[1], w445, w446);
  FullAdder U24 (w446, IN25[0], IN25[1], w447, w448);
  FullAdder U25 (w448, IN26[0], IN26[1], w449, w450);
  FullAdder U26 (w450, IN27[0], IN27[1], w451, w452);
  FullAdder U27 (w452, IN28[0], IN28[1], w453, w454);
  FullAdder U28 (w454, IN29[0], IN29[1], w455, w456);
  FullAdder U29 (w456, IN30[0], IN30[1], w457, w458);
  FullAdder U30 (w458, IN31[0], IN31[1], w459, w460);
  FullAdder U31 (w460, IN32[0], IN32[1], w461, w462);
  FullAdder U32 (w462, IN33[0], IN33[1], w463, w464);
  FullAdder U33 (w464, IN34[0], IN34[1], w465, w466);
  FullAdder U34 (w466, IN35[0], IN35[1], w467, w468);
  FullAdder U35 (w468, IN36[0], IN36[1], w469, w470);
  FullAdder U36 (w470, IN37[0], IN37[1], w471, w472);
  FullAdder U37 (w472, IN38[0], IN38[1], w473, w474);
  FullAdder U38 (w474, IN39[0], IN39[1], w475, w476);
  FullAdder U39 (w476, IN40[0], IN40[1], w477, w478);
  FullAdder U40 (w478, IN41[0], IN41[1], w479, w480);
  FullAdder U41 (w480, IN42[0], IN42[1], w481, w482);
  FullAdder U42 (w482, IN43[0], IN43[1], w483, w484);
  FullAdder U43 (w484, IN44[0], IN44[1], w485, w486);
  FullAdder U44 (w486, IN45[0], IN45[1], w487, w488);
  FullAdder U45 (w488, IN46[0], IN46[1], w489, w490);
  FullAdder U46 (w490, IN47[0], IN47[1], w491, w492);
  FullAdder U47 (w492, IN48[0], IN48[1], w493, w494);
  FullAdder U48 (w494, IN49[0], IN49[1], w495, w496);
  FullAdder U49 (w496, IN50[0], IN50[1], w497, w498);
  FullAdder U50 (w498, IN51[0], IN51[1], w499, w500);
  FullAdder U51 (w500, IN52[0], IN52[1], w501, w502);
  FullAdder U52 (w502, IN53[0], IN53[1], w503, w504);
  FullAdder U53 (w504, IN54[0], IN54[1], w505, w506);
  FullAdder U54 (w506, IN55[0], IN55[1], w507, w508);
  FullAdder U55 (w508, IN56[0], IN56[1], w509, w510);
  HalfAdder U56 (w401, IN2[2], Out1[2], w512);
  FullAdder U57 (w512, w403, IN3[2], w513, w514);
  FullAdder U58 (w514, w405, IN4[2], w515, w516);
  FullAdder U59 (w516, w407, IN5[2], w517, w518);
  FullAdder U60 (w518, w409, IN6[2], w519, w520);
  FullAdder U61 (w520, w411, IN7[2], w521, w522);
  FullAdder U62 (w522, w413, IN8[2], w523, w524);
  FullAdder U63 (w524, w415, IN9[2], w525, w526);
  FullAdder U64 (w526, w417, IN10[2], w527, w528);
  FullAdder U65 (w528, w419, IN11[2], w529, w530);
  FullAdder U66 (w530, w421, IN12[2], w531, w532);
  FullAdder U67 (w532, w423, IN13[2], w533, w534);
  FullAdder U68 (w534, w425, IN14[2], w535, w536);
  FullAdder U69 (w536, w427, IN15[2], w537, w538);
  FullAdder U70 (w538, w429, IN16[2], w539, w540);
  FullAdder U71 (w540, w431, IN17[2], w541, w542);
  FullAdder U72 (w542, w433, IN18[2], w543, w544);
  FullAdder U73 (w544, w435, IN19[2], w545, w546);
  FullAdder U74 (w546, w437, IN20[2], w547, w548);
  FullAdder U75 (w548, w439, IN21[2], w549, w550);
  FullAdder U76 (w550, w441, IN22[2], w551, w552);
  FullAdder U77 (w552, w443, IN23[2], w553, w554);
  FullAdder U78 (w554, w445, IN24[2], w555, w556);
  FullAdder U79 (w556, w447, IN25[2], w557, w558);
  FullAdder U80 (w558, w449, IN26[2], w559, w560);
  FullAdder U81 (w560, w451, IN27[2], w561, w562);
  FullAdder U82 (w562, w453, IN28[2], w563, w564);
  FullAdder U83 (w564, w455, IN29[2], w565, w566);
  FullAdder U84 (w566, w457, IN30[2], w567, w568);
  FullAdder U85 (w568, w459, IN31[2], w569, w570);
  FullAdder U86 (w570, w461, IN32[2], w571, w572);
  FullAdder U87 (w572, w463, IN33[2], w573, w574);
  FullAdder U88 (w574, w465, IN34[2], w575, w576);
  FullAdder U89 (w576, w467, IN35[2], w577, w578);
  FullAdder U90 (w578, w469, IN36[2], w579, w580);
  FullAdder U91 (w580, w471, IN37[2], w581, w582);
  FullAdder U92 (w582, w473, IN38[2], w583, w584);
  FullAdder U93 (w584, w475, IN39[2], w585, w586);
  FullAdder U94 (w586, w477, IN40[2], w587, w588);
  FullAdder U95 (w588, w479, IN41[2], w589, w590);
  FullAdder U96 (w590, w481, IN42[2], w591, w592);
  FullAdder U97 (w592, w483, IN43[2], w593, w594);
  FullAdder U98 (w594, w485, IN44[2], w595, w596);
  FullAdder U99 (w596, w487, IN45[2], w597, w598);
  FullAdder U100 (w598, w489, IN46[2], w599, w600);
  FullAdder U101 (w600, w491, IN47[2], w601, w602);
  FullAdder U102 (w602, w493, IN48[2], w603, w604);
  FullAdder U103 (w604, w495, IN49[2], w605, w606);
  FullAdder U104 (w606, w497, IN50[2], w607, w608);
  FullAdder U105 (w608, w499, IN51[2], w609, w610);
  FullAdder U106 (w610, w501, IN52[2], w611, w612);
  FullAdder U107 (w612, w503, IN53[2], w613, w614);
  FullAdder U108 (w614, w505, IN54[2], w615, w616);
  FullAdder U109 (w616, w507, IN55[2], w617, w618);
  FullAdder U110 (w618, w509, IN56[2], w619, w620);
  FullAdder U111 (w620, w510, IN57[0], w621, w622);
  HalfAdder U112 (w513, IN3[3], Out1[3], w624);
  FullAdder U113 (w624, w515, IN4[3], w625, w626);
  FullAdder U114 (w626, w517, IN5[3], w627, w628);
  FullAdder U115 (w628, w519, IN6[3], w629, w630);
  FullAdder U116 (w630, w521, IN7[3], w631, w632);
  FullAdder U117 (w632, w523, IN8[3], w633, w634);
  FullAdder U118 (w634, w525, IN9[3], w635, w636);
  FullAdder U119 (w636, w527, IN10[3], w637, w638);
  FullAdder U120 (w638, w529, IN11[3], w639, w640);
  FullAdder U121 (w640, w531, IN12[3], w641, w642);
  FullAdder U122 (w642, w533, IN13[3], w643, w644);
  FullAdder U123 (w644, w535, IN14[3], w645, w646);
  FullAdder U124 (w646, w537, IN15[3], w647, w648);
  FullAdder U125 (w648, w539, IN16[3], w649, w650);
  FullAdder U126 (w650, w541, IN17[3], w651, w652);
  FullAdder U127 (w652, w543, IN18[3], w653, w654);
  FullAdder U128 (w654, w545, IN19[3], w655, w656);
  FullAdder U129 (w656, w547, IN20[3], w657, w658);
  FullAdder U130 (w658, w549, IN21[3], w659, w660);
  FullAdder U131 (w660, w551, IN22[3], w661, w662);
  FullAdder U132 (w662, w553, IN23[3], w663, w664);
  FullAdder U133 (w664, w555, IN24[3], w665, w666);
  FullAdder U134 (w666, w557, IN25[3], w667, w668);
  FullAdder U135 (w668, w559, IN26[3], w669, w670);
  FullAdder U136 (w670, w561, IN27[3], w671, w672);
  FullAdder U137 (w672, w563, IN28[3], w673, w674);
  FullAdder U138 (w674, w565, IN29[3], w675, w676);
  FullAdder U139 (w676, w567, IN30[3], w677, w678);
  FullAdder U140 (w678, w569, IN31[3], w679, w680);
  FullAdder U141 (w680, w571, IN32[3], w681, w682);
  FullAdder U142 (w682, w573, IN33[3], w683, w684);
  FullAdder U143 (w684, w575, IN34[3], w685, w686);
  FullAdder U144 (w686, w577, IN35[3], w687, w688);
  FullAdder U145 (w688, w579, IN36[3], w689, w690);
  FullAdder U146 (w690, w581, IN37[3], w691, w692);
  FullAdder U147 (w692, w583, IN38[3], w693, w694);
  FullAdder U148 (w694, w585, IN39[3], w695, w696);
  FullAdder U149 (w696, w587, IN40[3], w697, w698);
  FullAdder U150 (w698, w589, IN41[3], w699, w700);
  FullAdder U151 (w700, w591, IN42[3], w701, w702);
  FullAdder U152 (w702, w593, IN43[3], w703, w704);
  FullAdder U153 (w704, w595, IN44[3], w705, w706);
  FullAdder U154 (w706, w597, IN45[3], w707, w708);
  FullAdder U155 (w708, w599, IN46[3], w709, w710);
  FullAdder U156 (w710, w601, IN47[3], w711, w712);
  FullAdder U157 (w712, w603, IN48[3], w713, w714);
  FullAdder U158 (w714, w605, IN49[3], w715, w716);
  FullAdder U159 (w716, w607, IN50[3], w717, w718);
  FullAdder U160 (w718, w609, IN51[3], w719, w720);
  FullAdder U161 (w720, w611, IN52[3], w721, w722);
  FullAdder U162 (w722, w613, IN53[3], w723, w724);
  FullAdder U163 (w724, w615, IN54[3], w725, w726);
  FullAdder U164 (w726, w617, IN55[3], w727, w728);
  FullAdder U165 (w728, w619, IN56[3], w729, w730);
  FullAdder U166 (w730, w621, IN57[1], w731, w732);
  FullAdder U167 (w732, w622, IN58[0], w733, w734);
  HalfAdder U168 (w625, IN4[4], Out1[4], w736);
  FullAdder U169 (w736, w627, IN5[4], w737, w738);
  FullAdder U170 (w738, w629, IN6[4], w739, w740);
  FullAdder U171 (w740, w631, IN7[4], w741, w742);
  FullAdder U172 (w742, w633, IN8[4], w743, w744);
  FullAdder U173 (w744, w635, IN9[4], w745, w746);
  FullAdder U174 (w746, w637, IN10[4], w747, w748);
  FullAdder U175 (w748, w639, IN11[4], w749, w750);
  FullAdder U176 (w750, w641, IN12[4], w751, w752);
  FullAdder U177 (w752, w643, IN13[4], w753, w754);
  FullAdder U178 (w754, w645, IN14[4], w755, w756);
  FullAdder U179 (w756, w647, IN15[4], w757, w758);
  FullAdder U180 (w758, w649, IN16[4], w759, w760);
  FullAdder U181 (w760, w651, IN17[4], w761, w762);
  FullAdder U182 (w762, w653, IN18[4], w763, w764);
  FullAdder U183 (w764, w655, IN19[4], w765, w766);
  FullAdder U184 (w766, w657, IN20[4], w767, w768);
  FullAdder U185 (w768, w659, IN21[4], w769, w770);
  FullAdder U186 (w770, w661, IN22[4], w771, w772);
  FullAdder U187 (w772, w663, IN23[4], w773, w774);
  FullAdder U188 (w774, w665, IN24[4], w775, w776);
  FullAdder U189 (w776, w667, IN25[4], w777, w778);
  FullAdder U190 (w778, w669, IN26[4], w779, w780);
  FullAdder U191 (w780, w671, IN27[4], w781, w782);
  FullAdder U192 (w782, w673, IN28[4], w783, w784);
  FullAdder U193 (w784, w675, IN29[4], w785, w786);
  FullAdder U194 (w786, w677, IN30[4], w787, w788);
  FullAdder U195 (w788, w679, IN31[4], w789, w790);
  FullAdder U196 (w790, w681, IN32[4], w791, w792);
  FullAdder U197 (w792, w683, IN33[4], w793, w794);
  FullAdder U198 (w794, w685, IN34[4], w795, w796);
  FullAdder U199 (w796, w687, IN35[4], w797, w798);
  FullAdder U200 (w798, w689, IN36[4], w799, w800);
  FullAdder U201 (w800, w691, IN37[4], w801, w802);
  FullAdder U202 (w802, w693, IN38[4], w803, w804);
  FullAdder U203 (w804, w695, IN39[4], w805, w806);
  FullAdder U204 (w806, w697, IN40[4], w807, w808);
  FullAdder U205 (w808, w699, IN41[4], w809, w810);
  FullAdder U206 (w810, w701, IN42[4], w811, w812);
  FullAdder U207 (w812, w703, IN43[4], w813, w814);
  FullAdder U208 (w814, w705, IN44[4], w815, w816);
  FullAdder U209 (w816, w707, IN45[4], w817, w818);
  FullAdder U210 (w818, w709, IN46[4], w819, w820);
  FullAdder U211 (w820, w711, IN47[4], w821, w822);
  FullAdder U212 (w822, w713, IN48[4], w823, w824);
  FullAdder U213 (w824, w715, IN49[4], w825, w826);
  FullAdder U214 (w826, w717, IN50[4], w827, w828);
  FullAdder U215 (w828, w719, IN51[4], w829, w830);
  FullAdder U216 (w830, w721, IN52[4], w831, w832);
  FullAdder U217 (w832, w723, IN53[4], w833, w834);
  FullAdder U218 (w834, w725, IN54[4], w835, w836);
  FullAdder U219 (w836, w727, IN55[4], w837, w838);
  FullAdder U220 (w838, w729, IN56[4], w839, w840);
  FullAdder U221 (w840, w731, IN57[2], w841, w842);
  FullAdder U222 (w842, w733, IN58[1], w843, w844);
  FullAdder U223 (w844, w734, IN59[0], w845, w846);
  HalfAdder U224 (w737, IN5[5], Out1[5], w848);
  FullAdder U225 (w848, w739, IN6[5], w849, w850);
  FullAdder U226 (w850, w741, IN7[5], w851, w852);
  FullAdder U227 (w852, w743, IN8[5], w853, w854);
  FullAdder U228 (w854, w745, IN9[5], w855, w856);
  FullAdder U229 (w856, w747, IN10[5], w857, w858);
  FullAdder U230 (w858, w749, IN11[5], w859, w860);
  FullAdder U231 (w860, w751, IN12[5], w861, w862);
  FullAdder U232 (w862, w753, IN13[5], w863, w864);
  FullAdder U233 (w864, w755, IN14[5], w865, w866);
  FullAdder U234 (w866, w757, IN15[5], w867, w868);
  FullAdder U235 (w868, w759, IN16[5], w869, w870);
  FullAdder U236 (w870, w761, IN17[5], w871, w872);
  FullAdder U237 (w872, w763, IN18[5], w873, w874);
  FullAdder U238 (w874, w765, IN19[5], w875, w876);
  FullAdder U239 (w876, w767, IN20[5], w877, w878);
  FullAdder U240 (w878, w769, IN21[5], w879, w880);
  FullAdder U241 (w880, w771, IN22[5], w881, w882);
  FullAdder U242 (w882, w773, IN23[5], w883, w884);
  FullAdder U243 (w884, w775, IN24[5], w885, w886);
  FullAdder U244 (w886, w777, IN25[5], w887, w888);
  FullAdder U245 (w888, w779, IN26[5], w889, w890);
  FullAdder U246 (w890, w781, IN27[5], w891, w892);
  FullAdder U247 (w892, w783, IN28[5], w893, w894);
  FullAdder U248 (w894, w785, IN29[5], w895, w896);
  FullAdder U249 (w896, w787, IN30[5], w897, w898);
  FullAdder U250 (w898, w789, IN31[5], w899, w900);
  FullAdder U251 (w900, w791, IN32[5], w901, w902);
  FullAdder U252 (w902, w793, IN33[5], w903, w904);
  FullAdder U253 (w904, w795, IN34[5], w905, w906);
  FullAdder U254 (w906, w797, IN35[5], w907, w908);
  FullAdder U255 (w908, w799, IN36[5], w909, w910);
  FullAdder U256 (w910, w801, IN37[5], w911, w912);
  FullAdder U257 (w912, w803, IN38[5], w913, w914);
  FullAdder U258 (w914, w805, IN39[5], w915, w916);
  FullAdder U259 (w916, w807, IN40[5], w917, w918);
  FullAdder U260 (w918, w809, IN41[5], w919, w920);
  FullAdder U261 (w920, w811, IN42[5], w921, w922);
  FullAdder U262 (w922, w813, IN43[5], w923, w924);
  FullAdder U263 (w924, w815, IN44[5], w925, w926);
  FullAdder U264 (w926, w817, IN45[5], w927, w928);
  FullAdder U265 (w928, w819, IN46[5], w929, w930);
  FullAdder U266 (w930, w821, IN47[5], w931, w932);
  FullAdder U267 (w932, w823, IN48[5], w933, w934);
  FullAdder U268 (w934, w825, IN49[5], w935, w936);
  FullAdder U269 (w936, w827, IN50[5], w937, w938);
  FullAdder U270 (w938, w829, IN51[5], w939, w940);
  FullAdder U271 (w940, w831, IN52[5], w941, w942);
  FullAdder U272 (w942, w833, IN53[5], w943, w944);
  FullAdder U273 (w944, w835, IN54[5], w945, w946);
  FullAdder U274 (w946, w837, IN55[5], w947, w948);
  FullAdder U275 (w948, w839, IN56[5], w949, w950);
  FullAdder U276 (w950, w841, IN57[3], w951, w952);
  FullAdder U277 (w952, w843, IN58[2], w953, w954);
  FullAdder U278 (w954, w845, IN59[1], w955, w956);
  FullAdder U279 (w956, w846, IN60[0], w957, w958);
  HalfAdder U280 (w849, IN6[6], Out1[6], w960);
  FullAdder U281 (w960, w851, IN7[6], Out1[7], w962);
  FullAdder U282 (w962, w853, IN8[6], Out1[8], w964);
  FullAdder U283 (w964, w855, IN9[6], Out1[9], w966);
  FullAdder U284 (w966, w857, IN10[6], Out1[10], w968);
  FullAdder U285 (w968, w859, IN11[6], Out1[11], w970);
  FullAdder U286 (w970, w861, IN12[6], Out1[12], w972);
  FullAdder U287 (w972, w863, IN13[6], Out1[13], w974);
  FullAdder U288 (w974, w865, IN14[6], Out1[14], w976);
  FullAdder U289 (w976, w867, IN15[6], Out1[15], w978);
  FullAdder U290 (w978, w869, IN16[6], Out1[16], w980);
  FullAdder U291 (w980, w871, IN17[6], Out1[17], w982);
  FullAdder U292 (w982, w873, IN18[6], Out1[18], w984);
  FullAdder U293 (w984, w875, IN19[6], Out1[19], w986);
  FullAdder U294 (w986, w877, IN20[6], Out1[20], w988);
  FullAdder U295 (w988, w879, IN21[6], Out1[21], w990);
  FullAdder U296 (w990, w881, IN22[6], Out1[22], w992);
  FullAdder U297 (w992, w883, IN23[6], Out1[23], w994);
  FullAdder U298 (w994, w885, IN24[6], Out1[24], w996);
  FullAdder U299 (w996, w887, IN25[6], Out1[25], w998);
  FullAdder U300 (w998, w889, IN26[6], Out1[26], w1000);
  FullAdder U301 (w1000, w891, IN27[6], Out1[27], w1002);
  FullAdder U302 (w1002, w893, IN28[6], Out1[28], w1004);
  FullAdder U303 (w1004, w895, IN29[6], Out1[29], w1006);
  FullAdder U304 (w1006, w897, IN30[6], Out1[30], w1008);
  FullAdder U305 (w1008, w899, IN31[6], Out1[31], w1010);
  FullAdder U306 (w1010, w901, IN32[6], Out1[32], w1012);
  FullAdder U307 (w1012, w903, IN33[6], Out1[33], w1014);
  FullAdder U308 (w1014, w905, IN34[6], Out1[34], w1016);
  FullAdder U309 (w1016, w907, IN35[6], Out1[35], w1018);
  FullAdder U310 (w1018, w909, IN36[6], Out1[36], w1020);
  FullAdder U311 (w1020, w911, IN37[6], Out1[37], w1022);
  FullAdder U312 (w1022, w913, IN38[6], Out1[38], w1024);
  FullAdder U313 (w1024, w915, IN39[6], Out1[39], w1026);
  FullAdder U314 (w1026, w917, IN40[6], Out1[40], w1028);
  FullAdder U315 (w1028, w919, IN41[6], Out1[41], w1030);
  FullAdder U316 (w1030, w921, IN42[6], Out1[42], w1032);
  FullAdder U317 (w1032, w923, IN43[6], Out1[43], w1034);
  FullAdder U318 (w1034, w925, IN44[6], Out1[44], w1036);
  FullAdder U319 (w1036, w927, IN45[6], Out1[45], w1038);
  FullAdder U320 (w1038, w929, IN46[6], Out1[46], w1040);
  FullAdder U321 (w1040, w931, IN47[6], Out1[47], w1042);
  FullAdder U322 (w1042, w933, IN48[6], Out1[48], w1044);
  FullAdder U323 (w1044, w935, IN49[6], Out1[49], w1046);
  FullAdder U324 (w1046, w937, IN50[6], Out1[50], w1048);
  FullAdder U325 (w1048, w939, IN51[6], Out1[51], w1050);
  FullAdder U326 (w1050, w941, IN52[6], Out1[52], w1052);
  FullAdder U327 (w1052, w943, IN53[6], Out1[53], w1054);
  FullAdder U328 (w1054, w945, IN54[6], Out1[54], w1056);
  FullAdder U329 (w1056, w947, IN55[6], Out1[55], w1058);
  FullAdder U330 (w1058, w949, IN56[6], Out1[56], w1060);
  FullAdder U331 (w1060, w951, IN57[4], Out1[57], w1062);
  FullAdder U332 (w1062, w953, IN58[3], Out1[58], w1064);
  FullAdder U333 (w1064, w955, IN59[2], Out1[59], w1066);
  FullAdder U334 (w1066, w957, IN60[1], Out1[60], w1068);
  FullAdder U335 (w1068, w958, IN61[0], Out1[61], Out1[62]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN57[5];
  assign Out2[1] = IN58[4];
  assign Out2[2] = IN59[3];
  assign Out2[3] = IN60[2];
  assign Out2[4] = IN61[1];
  assign Out2[5] = IN62[0];

endmodule
module RC_6_6(IN1, IN2, Out);
  input [5:0] IN1;
  input [5:0] IN2;
  output [6:0] Out;
  wire w13;
  wire w15;
  wire w17;
  wire w19;
  wire w21;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w13);
  FullAdder U1 (IN1[1], IN2[1], w13, Out[1], w15);
  FullAdder U2 (IN1[2], IN2[2], w15, Out[2], w17);
  FullAdder U3 (IN1[3], IN2[3], w17, Out[3], w19);
  FullAdder U4 (IN1[4], IN2[4], w19, Out[4], w21);
  FullAdder U5 (IN1[5], IN2[5], w21, Out[5], Out[6]);

endmodule
module NR_57_7(IN1, IN2, Out);
  input [56:0] IN1;
  input [6:0] IN2;
  output [63:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [6:0] P37;
  wire [6:0] P38;
  wire [6:0] P39;
  wire [6:0] P40;
  wire [6:0] P41;
  wire [6:0] P42;
  wire [6:0] P43;
  wire [6:0] P44;
  wire [6:0] P45;
  wire [6:0] P46;
  wire [6:0] P47;
  wire [6:0] P48;
  wire [6:0] P49;
  wire [6:0] P50;
  wire [6:0] P51;
  wire [6:0] P52;
  wire [6:0] P53;
  wire [6:0] P54;
  wire [6:0] P55;
  wire [6:0] P56;
  wire [5:0] P57;
  wire [4:0] P58;
  wire [3:0] P59;
  wire [2:0] P60;
  wire [1:0] P61;
  wire [0:0] P62;
  wire [62:0] R1;
  wire [5:0] R2;
  wire [63:0] aOut;
  U_SP_57_7 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, R1, R2);
  RC_6_6 S2 (R1[62:57], R2, aOut[63:57]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign Out = aOut[63:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
