
module customAdder58_0(
    input [57 : 0] A,
    input [57 : 0] B,
    output [58 : 0] Sum
);

    assign Sum = A+B;

endmodule
