
module NR_62_1(
    input [61:0]IN1,
    input [0:0]IN2,
    output [61:0]Out
);
    assign Out = IN2;
endmodule
