
module NR_34_1(
    input [33:0]IN1,
    input [0:0]IN2,
    output [33:0]Out
);
    assign Out = IN2;
endmodule
