//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 4
  second input length: 48
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_4_48(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50);
  input [3:0] IN1;
  input [47:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [3:0] P4;
  output [3:0] P5;
  output [3:0] P6;
  output [3:0] P7;
  output [3:0] P8;
  output [3:0] P9;
  output [3:0] P10;
  output [3:0] P11;
  output [3:0] P12;
  output [3:0] P13;
  output [3:0] P14;
  output [3:0] P15;
  output [3:0] P16;
  output [3:0] P17;
  output [3:0] P18;
  output [3:0] P19;
  output [3:0] P20;
  output [3:0] P21;
  output [3:0] P22;
  output [3:0] P23;
  output [3:0] P24;
  output [3:0] P25;
  output [3:0] P26;
  output [3:0] P27;
  output [3:0] P28;
  output [3:0] P29;
  output [3:0] P30;
  output [3:0] P31;
  output [3:0] P32;
  output [3:0] P33;
  output [3:0] P34;
  output [3:0] P35;
  output [3:0] P36;
  output [3:0] P37;
  output [3:0] P38;
  output [3:0] P39;
  output [3:0] P40;
  output [3:0] P41;
  output [3:0] P42;
  output [3:0] P43;
  output [3:0] P44;
  output [3:0] P45;
  output [3:0] P46;
  output [3:0] P47;
  output [2:0] P48;
  output [1:0] P49;
  output [0:0] P50;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[0] = IN1[1]&IN2[47];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[1] = IN1[2]&IN2[46];
  assign P49[0] = IN1[2]&IN2[47];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[2] = IN1[3]&IN2[45];
  assign P49[1] = IN1[3]&IN2[46];
  assign P50[0] = IN1[3]&IN2[47];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [3:0] IN4;
  input [3:0] IN5;
  input [3:0] IN6;
  input [3:0] IN7;
  input [3:0] IN8;
  input [3:0] IN9;
  input [3:0] IN10;
  input [3:0] IN11;
  input [3:0] IN12;
  input [3:0] IN13;
  input [3:0] IN14;
  input [3:0] IN15;
  input [3:0] IN16;
  input [3:0] IN17;
  input [3:0] IN18;
  input [3:0] IN19;
  input [3:0] IN20;
  input [3:0] IN21;
  input [3:0] IN22;
  input [3:0] IN23;
  input [3:0] IN24;
  input [3:0] IN25;
  input [3:0] IN26;
  input [3:0] IN27;
  input [3:0] IN28;
  input [3:0] IN29;
  input [3:0] IN30;
  input [3:0] IN31;
  input [3:0] IN32;
  input [3:0] IN33;
  input [3:0] IN34;
  input [3:0] IN35;
  input [3:0] IN36;
  input [3:0] IN37;
  input [3:0] IN38;
  input [3:0] IN39;
  input [3:0] IN40;
  input [3:0] IN41;
  input [3:0] IN42;
  input [3:0] IN43;
  input [3:0] IN44;
  input [3:0] IN45;
  input [3:0] IN46;
  input [3:0] IN47;
  input [2:0] IN48;
  input [1:0] IN49;
  input [0:0] IN50;
  output [50:0] Out1;
  output [46:0] Out2;
  wire w193;
  wire w194;
  wire w195;
  wire w196;
  wire w197;
  wire w199;
  wire w200;
  wire w201;
  wire w202;
  wire w203;
  wire w205;
  wire w206;
  wire w207;
  wire w208;
  wire w209;
  wire w211;
  wire w212;
  wire w213;
  wire w214;
  wire w215;
  wire w217;
  wire w218;
  wire w219;
  wire w220;
  wire w221;
  wire w223;
  wire w224;
  wire w225;
  wire w226;
  wire w227;
  wire w229;
  wire w230;
  wire w231;
  wire w232;
  wire w233;
  wire w235;
  wire w236;
  wire w237;
  wire w238;
  wire w239;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w247;
  wire w248;
  wire w249;
  wire w250;
  wire w251;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w469;
  wire w471;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w193);
  FullAdder U1 (w193, IN2[0], IN2[1], w194, w195);
  FullAdder U2 (w195, IN3[0], IN3[1], w196, w197);
  HalfAdder U3 (w194, IN2[2], Out1[2], w199);
  FullAdder U4 (w199, w196, IN3[2], w200, w201);
  FullAdder U5 (w201, w197, IN4[0], w202, w203);
  HalfAdder U6 (w200, IN3[3], Out1[3], w205);
  FullAdder U7 (w205, w202, IN4[1], w206, w207);
  FullAdder U8 (w207, w203, IN5[0], w208, w209);
  HalfAdder U9 (w206, IN4[2], Out1[4], w211);
  FullAdder U10 (w211, w208, IN5[1], w212, w213);
  FullAdder U11 (w213, w209, IN6[0], w214, w215);
  HalfAdder U12 (w212, IN5[2], Out1[5], w217);
  FullAdder U13 (w217, w214, IN6[1], w218, w219);
  FullAdder U14 (w219, w215, IN7[0], w220, w221);
  HalfAdder U15 (w218, IN6[2], Out1[6], w223);
  FullAdder U16 (w223, w220, IN7[1], w224, w225);
  FullAdder U17 (w225, w221, IN8[0], w226, w227);
  HalfAdder U18 (w224, IN7[2], Out1[7], w229);
  FullAdder U19 (w229, w226, IN8[1], w230, w231);
  FullAdder U20 (w231, w227, IN9[0], w232, w233);
  HalfAdder U21 (w230, IN8[2], Out1[8], w235);
  FullAdder U22 (w235, w232, IN9[1], w236, w237);
  FullAdder U23 (w237, w233, IN10[0], w238, w239);
  HalfAdder U24 (w236, IN9[2], Out1[9], w241);
  FullAdder U25 (w241, w238, IN10[1], w242, w243);
  FullAdder U26 (w243, w239, IN11[0], w244, w245);
  HalfAdder U27 (w242, IN10[2], Out1[10], w247);
  FullAdder U28 (w247, w244, IN11[1], w248, w249);
  FullAdder U29 (w249, w245, IN12[0], w250, w251);
  HalfAdder U30 (w248, IN11[2], Out1[11], w253);
  FullAdder U31 (w253, w250, IN12[1], w254, w255);
  FullAdder U32 (w255, w251, IN13[0], w256, w257);
  HalfAdder U33 (w254, IN12[2], Out1[12], w259);
  FullAdder U34 (w259, w256, IN13[1], w260, w261);
  FullAdder U35 (w261, w257, IN14[0], w262, w263);
  HalfAdder U36 (w260, IN13[2], Out1[13], w265);
  FullAdder U37 (w265, w262, IN14[1], w266, w267);
  FullAdder U38 (w267, w263, IN15[0], w268, w269);
  HalfAdder U39 (w266, IN14[2], Out1[14], w271);
  FullAdder U40 (w271, w268, IN15[1], w272, w273);
  FullAdder U41 (w273, w269, IN16[0], w274, w275);
  HalfAdder U42 (w272, IN15[2], Out1[15], w277);
  FullAdder U43 (w277, w274, IN16[1], w278, w279);
  FullAdder U44 (w279, w275, IN17[0], w280, w281);
  HalfAdder U45 (w278, IN16[2], Out1[16], w283);
  FullAdder U46 (w283, w280, IN17[1], w284, w285);
  FullAdder U47 (w285, w281, IN18[0], w286, w287);
  HalfAdder U48 (w284, IN17[2], Out1[17], w289);
  FullAdder U49 (w289, w286, IN18[1], w290, w291);
  FullAdder U50 (w291, w287, IN19[0], w292, w293);
  HalfAdder U51 (w290, IN18[2], Out1[18], w295);
  FullAdder U52 (w295, w292, IN19[1], w296, w297);
  FullAdder U53 (w297, w293, IN20[0], w298, w299);
  HalfAdder U54 (w296, IN19[2], Out1[19], w301);
  FullAdder U55 (w301, w298, IN20[1], w302, w303);
  FullAdder U56 (w303, w299, IN21[0], w304, w305);
  HalfAdder U57 (w302, IN20[2], Out1[20], w307);
  FullAdder U58 (w307, w304, IN21[1], w308, w309);
  FullAdder U59 (w309, w305, IN22[0], w310, w311);
  HalfAdder U60 (w308, IN21[2], Out1[21], w313);
  FullAdder U61 (w313, w310, IN22[1], w314, w315);
  FullAdder U62 (w315, w311, IN23[0], w316, w317);
  HalfAdder U63 (w314, IN22[2], Out1[22], w319);
  FullAdder U64 (w319, w316, IN23[1], w320, w321);
  FullAdder U65 (w321, w317, IN24[0], w322, w323);
  HalfAdder U66 (w320, IN23[2], Out1[23], w325);
  FullAdder U67 (w325, w322, IN24[1], w326, w327);
  FullAdder U68 (w327, w323, IN25[0], w328, w329);
  HalfAdder U69 (w326, IN24[2], Out1[24], w331);
  FullAdder U70 (w331, w328, IN25[1], w332, w333);
  FullAdder U71 (w333, w329, IN26[0], w334, w335);
  HalfAdder U72 (w332, IN25[2], Out1[25], w337);
  FullAdder U73 (w337, w334, IN26[1], w338, w339);
  FullAdder U74 (w339, w335, IN27[0], w340, w341);
  HalfAdder U75 (w338, IN26[2], Out1[26], w343);
  FullAdder U76 (w343, w340, IN27[1], w344, w345);
  FullAdder U77 (w345, w341, IN28[0], w346, w347);
  HalfAdder U78 (w344, IN27[2], Out1[27], w349);
  FullAdder U79 (w349, w346, IN28[1], w350, w351);
  FullAdder U80 (w351, w347, IN29[0], w352, w353);
  HalfAdder U81 (w350, IN28[2], Out1[28], w355);
  FullAdder U82 (w355, w352, IN29[1], w356, w357);
  FullAdder U83 (w357, w353, IN30[0], w358, w359);
  HalfAdder U84 (w356, IN29[2], Out1[29], w361);
  FullAdder U85 (w361, w358, IN30[1], w362, w363);
  FullAdder U86 (w363, w359, IN31[0], w364, w365);
  HalfAdder U87 (w362, IN30[2], Out1[30], w367);
  FullAdder U88 (w367, w364, IN31[1], w368, w369);
  FullAdder U89 (w369, w365, IN32[0], w370, w371);
  HalfAdder U90 (w368, IN31[2], Out1[31], w373);
  FullAdder U91 (w373, w370, IN32[1], w374, w375);
  FullAdder U92 (w375, w371, IN33[0], w376, w377);
  HalfAdder U93 (w374, IN32[2], Out1[32], w379);
  FullAdder U94 (w379, w376, IN33[1], w380, w381);
  FullAdder U95 (w381, w377, IN34[0], w382, w383);
  HalfAdder U96 (w380, IN33[2], Out1[33], w385);
  FullAdder U97 (w385, w382, IN34[1], w386, w387);
  FullAdder U98 (w387, w383, IN35[0], w388, w389);
  HalfAdder U99 (w386, IN34[2], Out1[34], w391);
  FullAdder U100 (w391, w388, IN35[1], w392, w393);
  FullAdder U101 (w393, w389, IN36[0], w394, w395);
  HalfAdder U102 (w392, IN35[2], Out1[35], w397);
  FullAdder U103 (w397, w394, IN36[1], w398, w399);
  FullAdder U104 (w399, w395, IN37[0], w400, w401);
  HalfAdder U105 (w398, IN36[2], Out1[36], w403);
  FullAdder U106 (w403, w400, IN37[1], w404, w405);
  FullAdder U107 (w405, w401, IN38[0], w406, w407);
  HalfAdder U108 (w404, IN37[2], Out1[37], w409);
  FullAdder U109 (w409, w406, IN38[1], w410, w411);
  FullAdder U110 (w411, w407, IN39[0], w412, w413);
  HalfAdder U111 (w410, IN38[2], Out1[38], w415);
  FullAdder U112 (w415, w412, IN39[1], w416, w417);
  FullAdder U113 (w417, w413, IN40[0], w418, w419);
  HalfAdder U114 (w416, IN39[2], Out1[39], w421);
  FullAdder U115 (w421, w418, IN40[1], w422, w423);
  FullAdder U116 (w423, w419, IN41[0], w424, w425);
  HalfAdder U117 (w422, IN40[2], Out1[40], w427);
  FullAdder U118 (w427, w424, IN41[1], w428, w429);
  FullAdder U119 (w429, w425, IN42[0], w430, w431);
  HalfAdder U120 (w428, IN41[2], Out1[41], w433);
  FullAdder U121 (w433, w430, IN42[1], w434, w435);
  FullAdder U122 (w435, w431, IN43[0], w436, w437);
  HalfAdder U123 (w434, IN42[2], Out1[42], w439);
  FullAdder U124 (w439, w436, IN43[1], w440, w441);
  FullAdder U125 (w441, w437, IN44[0], w442, w443);
  HalfAdder U126 (w440, IN43[2], Out1[43], w445);
  FullAdder U127 (w445, w442, IN44[1], w446, w447);
  FullAdder U128 (w447, w443, IN45[0], w448, w449);
  HalfAdder U129 (w446, IN44[2], Out1[44], w451);
  FullAdder U130 (w451, w448, IN45[1], w452, w453);
  FullAdder U131 (w453, w449, IN46[0], w454, w455);
  HalfAdder U132 (w452, IN45[2], Out1[45], w457);
  FullAdder U133 (w457, w454, IN46[1], w458, w459);
  FullAdder U134 (w459, w455, IN47[0], w460, w461);
  HalfAdder U135 (w458, IN46[2], Out1[46], w463);
  FullAdder U136 (w463, w460, IN47[1], w464, w465);
  FullAdder U137 (w465, w461, IN48[0], w466, w467);
  HalfAdder U138 (w464, IN47[2], Out1[47], w469);
  FullAdder U139 (w469, w466, IN48[1], Out1[48], w471);
  FullAdder U140 (w471, w467, IN49[0], Out1[49], Out1[50]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN4[3];
  assign Out2[1] = IN5[3];
  assign Out2[2] = IN6[3];
  assign Out2[3] = IN7[3];
  assign Out2[4] = IN8[3];
  assign Out2[5] = IN9[3];
  assign Out2[6] = IN10[3];
  assign Out2[7] = IN11[3];
  assign Out2[8] = IN12[3];
  assign Out2[9] = IN13[3];
  assign Out2[10] = IN14[3];
  assign Out2[11] = IN15[3];
  assign Out2[12] = IN16[3];
  assign Out2[13] = IN17[3];
  assign Out2[14] = IN18[3];
  assign Out2[15] = IN19[3];
  assign Out2[16] = IN20[3];
  assign Out2[17] = IN21[3];
  assign Out2[18] = IN22[3];
  assign Out2[19] = IN23[3];
  assign Out2[20] = IN24[3];
  assign Out2[21] = IN25[3];
  assign Out2[22] = IN26[3];
  assign Out2[23] = IN27[3];
  assign Out2[24] = IN28[3];
  assign Out2[25] = IN29[3];
  assign Out2[26] = IN30[3];
  assign Out2[27] = IN31[3];
  assign Out2[28] = IN32[3];
  assign Out2[29] = IN33[3];
  assign Out2[30] = IN34[3];
  assign Out2[31] = IN35[3];
  assign Out2[32] = IN36[3];
  assign Out2[33] = IN37[3];
  assign Out2[34] = IN38[3];
  assign Out2[35] = IN39[3];
  assign Out2[36] = IN40[3];
  assign Out2[37] = IN41[3];
  assign Out2[38] = IN42[3];
  assign Out2[39] = IN43[3];
  assign Out2[40] = IN44[3];
  assign Out2[41] = IN45[3];
  assign Out2[42] = IN46[3];
  assign Out2[43] = IN47[3];
  assign Out2[44] = IN48[2];
  assign Out2[45] = IN49[1];
  assign Out2[46] = IN50[0];

endmodule
module RC_47_47(IN1, IN2, Out);
  input [46:0] IN1;
  input [46:0] IN2;
  output [47:0] Out;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w95);
  FullAdder U1 (IN1[1], IN2[1], w95, Out[1], w97);
  FullAdder U2 (IN1[2], IN2[2], w97, Out[2], w99);
  FullAdder U3 (IN1[3], IN2[3], w99, Out[3], w101);
  FullAdder U4 (IN1[4], IN2[4], w101, Out[4], w103);
  FullAdder U5 (IN1[5], IN2[5], w103, Out[5], w105);
  FullAdder U6 (IN1[6], IN2[6], w105, Out[6], w107);
  FullAdder U7 (IN1[7], IN2[7], w107, Out[7], w109);
  FullAdder U8 (IN1[8], IN2[8], w109, Out[8], w111);
  FullAdder U9 (IN1[9], IN2[9], w111, Out[9], w113);
  FullAdder U10 (IN1[10], IN2[10], w113, Out[10], w115);
  FullAdder U11 (IN1[11], IN2[11], w115, Out[11], w117);
  FullAdder U12 (IN1[12], IN2[12], w117, Out[12], w119);
  FullAdder U13 (IN1[13], IN2[13], w119, Out[13], w121);
  FullAdder U14 (IN1[14], IN2[14], w121, Out[14], w123);
  FullAdder U15 (IN1[15], IN2[15], w123, Out[15], w125);
  FullAdder U16 (IN1[16], IN2[16], w125, Out[16], w127);
  FullAdder U17 (IN1[17], IN2[17], w127, Out[17], w129);
  FullAdder U18 (IN1[18], IN2[18], w129, Out[18], w131);
  FullAdder U19 (IN1[19], IN2[19], w131, Out[19], w133);
  FullAdder U20 (IN1[20], IN2[20], w133, Out[20], w135);
  FullAdder U21 (IN1[21], IN2[21], w135, Out[21], w137);
  FullAdder U22 (IN1[22], IN2[22], w137, Out[22], w139);
  FullAdder U23 (IN1[23], IN2[23], w139, Out[23], w141);
  FullAdder U24 (IN1[24], IN2[24], w141, Out[24], w143);
  FullAdder U25 (IN1[25], IN2[25], w143, Out[25], w145);
  FullAdder U26 (IN1[26], IN2[26], w145, Out[26], w147);
  FullAdder U27 (IN1[27], IN2[27], w147, Out[27], w149);
  FullAdder U28 (IN1[28], IN2[28], w149, Out[28], w151);
  FullAdder U29 (IN1[29], IN2[29], w151, Out[29], w153);
  FullAdder U30 (IN1[30], IN2[30], w153, Out[30], w155);
  FullAdder U31 (IN1[31], IN2[31], w155, Out[31], w157);
  FullAdder U32 (IN1[32], IN2[32], w157, Out[32], w159);
  FullAdder U33 (IN1[33], IN2[33], w159, Out[33], w161);
  FullAdder U34 (IN1[34], IN2[34], w161, Out[34], w163);
  FullAdder U35 (IN1[35], IN2[35], w163, Out[35], w165);
  FullAdder U36 (IN1[36], IN2[36], w165, Out[36], w167);
  FullAdder U37 (IN1[37], IN2[37], w167, Out[37], w169);
  FullAdder U38 (IN1[38], IN2[38], w169, Out[38], w171);
  FullAdder U39 (IN1[39], IN2[39], w171, Out[39], w173);
  FullAdder U40 (IN1[40], IN2[40], w173, Out[40], w175);
  FullAdder U41 (IN1[41], IN2[41], w175, Out[41], w177);
  FullAdder U42 (IN1[42], IN2[42], w177, Out[42], w179);
  FullAdder U43 (IN1[43], IN2[43], w179, Out[43], w181);
  FullAdder U44 (IN1[44], IN2[44], w181, Out[44], w183);
  FullAdder U45 (IN1[45], IN2[45], w183, Out[45], w185);
  FullAdder U46 (IN1[46], IN2[46], w185, Out[46], Out[47]);

endmodule
module NR_4_48(IN1, IN2, Out);
  input [3:0] IN1;
  input [47:0] IN2;
  output [51:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [3:0] P4;
  wire [3:0] P5;
  wire [3:0] P6;
  wire [3:0] P7;
  wire [3:0] P8;
  wire [3:0] P9;
  wire [3:0] P10;
  wire [3:0] P11;
  wire [3:0] P12;
  wire [3:0] P13;
  wire [3:0] P14;
  wire [3:0] P15;
  wire [3:0] P16;
  wire [3:0] P17;
  wire [3:0] P18;
  wire [3:0] P19;
  wire [3:0] P20;
  wire [3:0] P21;
  wire [3:0] P22;
  wire [3:0] P23;
  wire [3:0] P24;
  wire [3:0] P25;
  wire [3:0] P26;
  wire [3:0] P27;
  wire [3:0] P28;
  wire [3:0] P29;
  wire [3:0] P30;
  wire [3:0] P31;
  wire [3:0] P32;
  wire [3:0] P33;
  wire [3:0] P34;
  wire [3:0] P35;
  wire [3:0] P36;
  wire [3:0] P37;
  wire [3:0] P38;
  wire [3:0] P39;
  wire [3:0] P40;
  wire [3:0] P41;
  wire [3:0] P42;
  wire [3:0] P43;
  wire [3:0] P44;
  wire [3:0] P45;
  wire [3:0] P46;
  wire [3:0] P47;
  wire [2:0] P48;
  wire [1:0] P49;
  wire [0:0] P50;
  wire [50:0] R1;
  wire [46:0] R2;
  wire [51:0] aOut;
  U_SP_4_48 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, R1, R2);
  RC_47_47 S2 (R1[50:4], R2, aOut[51:4]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign Out = aOut[51:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
