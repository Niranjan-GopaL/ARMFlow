
module NR_1_53(
    input [0:0]IN1,
    input [52:0]IN2,
    output [52:0]Out
);
    assign Out = IN2;
endmodule
