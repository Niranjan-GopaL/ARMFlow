
module customAdder48_0(
    input [47 : 0] A,
    input [47 : 0] B,
    output [48 : 0] Sum
);

    assign Sum = A+B;

endmodule
