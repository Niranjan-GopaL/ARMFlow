//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 10
  second input length: 55
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_10_55(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63);
  input [9:0] IN1;
  input [54:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [9:0] P10;
  output [9:0] P11;
  output [9:0] P12;
  output [9:0] P13;
  output [9:0] P14;
  output [9:0] P15;
  output [9:0] P16;
  output [9:0] P17;
  output [9:0] P18;
  output [9:0] P19;
  output [9:0] P20;
  output [9:0] P21;
  output [9:0] P22;
  output [9:0] P23;
  output [9:0] P24;
  output [9:0] P25;
  output [9:0] P26;
  output [9:0] P27;
  output [9:0] P28;
  output [9:0] P29;
  output [9:0] P30;
  output [9:0] P31;
  output [9:0] P32;
  output [9:0] P33;
  output [9:0] P34;
  output [9:0] P35;
  output [9:0] P36;
  output [9:0] P37;
  output [9:0] P38;
  output [9:0] P39;
  output [9:0] P40;
  output [9:0] P41;
  output [9:0] P42;
  output [9:0] P43;
  output [9:0] P44;
  output [9:0] P45;
  output [9:0] P46;
  output [9:0] P47;
  output [9:0] P48;
  output [9:0] P49;
  output [9:0] P50;
  output [9:0] P51;
  output [9:0] P52;
  output [9:0] P53;
  output [9:0] P54;
  output [8:0] P55;
  output [7:0] P56;
  output [6:0] P57;
  output [5:0] P58;
  output [4:0] P59;
  output [3:0] P60;
  output [2:0] P61;
  output [1:0] P62;
  output [0:0] P63;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[0] = IN1[1]&IN2[54];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[1] = IN1[2]&IN2[53];
  assign P56[0] = IN1[2]&IN2[54];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[2] = IN1[3]&IN2[52];
  assign P56[1] = IN1[3]&IN2[53];
  assign P57[0] = IN1[3]&IN2[54];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[3] = IN1[4]&IN2[51];
  assign P56[2] = IN1[4]&IN2[52];
  assign P57[1] = IN1[4]&IN2[53];
  assign P58[0] = IN1[4]&IN2[54];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[4] = IN1[5]&IN2[50];
  assign P56[3] = IN1[5]&IN2[51];
  assign P57[2] = IN1[5]&IN2[52];
  assign P58[1] = IN1[5]&IN2[53];
  assign P59[0] = IN1[5]&IN2[54];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[5] = IN1[6]&IN2[49];
  assign P56[4] = IN1[6]&IN2[50];
  assign P57[3] = IN1[6]&IN2[51];
  assign P58[2] = IN1[6]&IN2[52];
  assign P59[1] = IN1[6]&IN2[53];
  assign P60[0] = IN1[6]&IN2[54];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[7] = IN1[7]&IN2[47];
  assign P55[6] = IN1[7]&IN2[48];
  assign P56[5] = IN1[7]&IN2[49];
  assign P57[4] = IN1[7]&IN2[50];
  assign P58[3] = IN1[7]&IN2[51];
  assign P59[2] = IN1[7]&IN2[52];
  assign P60[1] = IN1[7]&IN2[53];
  assign P61[0] = IN1[7]&IN2[54];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[8] = IN1[8]&IN2[45];
  assign P54[8] = IN1[8]&IN2[46];
  assign P55[7] = IN1[8]&IN2[47];
  assign P56[6] = IN1[8]&IN2[48];
  assign P57[5] = IN1[8]&IN2[49];
  assign P58[4] = IN1[8]&IN2[50];
  assign P59[3] = IN1[8]&IN2[51];
  assign P60[2] = IN1[8]&IN2[52];
  assign P61[1] = IN1[8]&IN2[53];
  assign P62[0] = IN1[8]&IN2[54];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[9] = IN1[9]&IN2[44];
  assign P54[9] = IN1[9]&IN2[45];
  assign P55[8] = IN1[9]&IN2[46];
  assign P56[7] = IN1[9]&IN2[47];
  assign P57[6] = IN1[9]&IN2[48];
  assign P58[5] = IN1[9]&IN2[49];
  assign P59[4] = IN1[9]&IN2[50];
  assign P60[3] = IN1[9]&IN2[51];
  assign P61[2] = IN1[9]&IN2[52];
  assign P62[1] = IN1[9]&IN2[53];
  assign P63[0] = IN1[9]&IN2[54];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [9:0] IN10;
  input [9:0] IN11;
  input [9:0] IN12;
  input [9:0] IN13;
  input [9:0] IN14;
  input [9:0] IN15;
  input [9:0] IN16;
  input [9:0] IN17;
  input [9:0] IN18;
  input [9:0] IN19;
  input [9:0] IN20;
  input [9:0] IN21;
  input [9:0] IN22;
  input [9:0] IN23;
  input [9:0] IN24;
  input [9:0] IN25;
  input [9:0] IN26;
  input [9:0] IN27;
  input [9:0] IN28;
  input [9:0] IN29;
  input [9:0] IN30;
  input [9:0] IN31;
  input [9:0] IN32;
  input [9:0] IN33;
  input [9:0] IN34;
  input [9:0] IN35;
  input [9:0] IN36;
  input [9:0] IN37;
  input [9:0] IN38;
  input [9:0] IN39;
  input [9:0] IN40;
  input [9:0] IN41;
  input [9:0] IN42;
  input [9:0] IN43;
  input [9:0] IN44;
  input [9:0] IN45;
  input [9:0] IN46;
  input [9:0] IN47;
  input [9:0] IN48;
  input [9:0] IN49;
  input [9:0] IN50;
  input [9:0] IN51;
  input [9:0] IN52;
  input [9:0] IN53;
  input [9:0] IN54;
  input [8:0] IN55;
  input [7:0] IN56;
  input [6:0] IN57;
  input [5:0] IN58;
  input [4:0] IN59;
  input [3:0] IN60;
  input [2:0] IN61;
  input [1:0] IN62;
  input [0:0] IN63;
  output [63:0] Out1;
  output [53:0] Out2;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1505;
  wire w1507;
  wire w1509;
  wire w1511;
  wire w1513;
  wire w1515;
  wire w1517;
  wire w1519;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w551);
  FullAdder U1 (w551, IN2[0], IN2[1], w552, w553);
  FullAdder U2 (w553, IN3[0], IN3[1], w554, w555);
  FullAdder U3 (w555, IN4[0], IN4[1], w556, w557);
  FullAdder U4 (w557, IN5[0], IN5[1], w558, w559);
  FullAdder U5 (w559, IN6[0], IN6[1], w560, w561);
  FullAdder U6 (w561, IN7[0], IN7[1], w562, w563);
  FullAdder U7 (w563, IN8[0], IN8[1], w564, w565);
  FullAdder U8 (w565, IN9[0], IN9[1], w566, w567);
  HalfAdder U9 (w552, IN2[2], Out1[2], w569);
  FullAdder U10 (w569, w554, IN3[2], w570, w571);
  FullAdder U11 (w571, w556, IN4[2], w572, w573);
  FullAdder U12 (w573, w558, IN5[2], w574, w575);
  FullAdder U13 (w575, w560, IN6[2], w576, w577);
  FullAdder U14 (w577, w562, IN7[2], w578, w579);
  FullAdder U15 (w579, w564, IN8[2], w580, w581);
  FullAdder U16 (w581, w566, IN9[2], w582, w583);
  FullAdder U17 (w583, w567, IN10[0], w584, w585);
  HalfAdder U18 (w570, IN3[3], Out1[3], w587);
  FullAdder U19 (w587, w572, IN4[3], w588, w589);
  FullAdder U20 (w589, w574, IN5[3], w590, w591);
  FullAdder U21 (w591, w576, IN6[3], w592, w593);
  FullAdder U22 (w593, w578, IN7[3], w594, w595);
  FullAdder U23 (w595, w580, IN8[3], w596, w597);
  FullAdder U24 (w597, w582, IN9[3], w598, w599);
  FullAdder U25 (w599, w584, IN10[1], w600, w601);
  FullAdder U26 (w601, w585, IN11[0], w602, w603);
  HalfAdder U27 (w588, IN4[4], Out1[4], w605);
  FullAdder U28 (w605, w590, IN5[4], w606, w607);
  FullAdder U29 (w607, w592, IN6[4], w608, w609);
  FullAdder U30 (w609, w594, IN7[4], w610, w611);
  FullAdder U31 (w611, w596, IN8[4], w612, w613);
  FullAdder U32 (w613, w598, IN9[4], w614, w615);
  FullAdder U33 (w615, w600, IN10[2], w616, w617);
  FullAdder U34 (w617, w602, IN11[1], w618, w619);
  FullAdder U35 (w619, w603, IN12[0], w620, w621);
  HalfAdder U36 (w606, IN5[5], Out1[5], w623);
  FullAdder U37 (w623, w608, IN6[5], w624, w625);
  FullAdder U38 (w625, w610, IN7[5], w626, w627);
  FullAdder U39 (w627, w612, IN8[5], w628, w629);
  FullAdder U40 (w629, w614, IN9[5], w630, w631);
  FullAdder U41 (w631, w616, IN10[3], w632, w633);
  FullAdder U42 (w633, w618, IN11[2], w634, w635);
  FullAdder U43 (w635, w620, IN12[1], w636, w637);
  FullAdder U44 (w637, w621, IN13[0], w638, w639);
  HalfAdder U45 (w624, IN6[6], Out1[6], w641);
  FullAdder U46 (w641, w626, IN7[6], w642, w643);
  FullAdder U47 (w643, w628, IN8[6], w644, w645);
  FullAdder U48 (w645, w630, IN9[6], w646, w647);
  FullAdder U49 (w647, w632, IN10[4], w648, w649);
  FullAdder U50 (w649, w634, IN11[3], w650, w651);
  FullAdder U51 (w651, w636, IN12[2], w652, w653);
  FullAdder U52 (w653, w638, IN13[1], w654, w655);
  FullAdder U53 (w655, w639, IN14[0], w656, w657);
  HalfAdder U54 (w642, IN7[7], Out1[7], w659);
  FullAdder U55 (w659, w644, IN8[7], w660, w661);
  FullAdder U56 (w661, w646, IN9[7], w662, w663);
  FullAdder U57 (w663, w648, IN10[5], w664, w665);
  FullAdder U58 (w665, w650, IN11[4], w666, w667);
  FullAdder U59 (w667, w652, IN12[3], w668, w669);
  FullAdder U60 (w669, w654, IN13[2], w670, w671);
  FullAdder U61 (w671, w656, IN14[1], w672, w673);
  FullAdder U62 (w673, w657, IN15[0], w674, w675);
  HalfAdder U63 (w660, IN8[8], Out1[8], w677);
  FullAdder U64 (w677, w662, IN9[8], w678, w679);
  FullAdder U65 (w679, w664, IN10[6], w680, w681);
  FullAdder U66 (w681, w666, IN11[5], w682, w683);
  FullAdder U67 (w683, w668, IN12[4], w684, w685);
  FullAdder U68 (w685, w670, IN13[3], w686, w687);
  FullAdder U69 (w687, w672, IN14[2], w688, w689);
  FullAdder U70 (w689, w674, IN15[1], w690, w691);
  FullAdder U71 (w691, w675, IN16[0], w692, w693);
  HalfAdder U72 (w678, IN9[9], Out1[9], w695);
  FullAdder U73 (w695, w680, IN10[7], w696, w697);
  FullAdder U74 (w697, w682, IN11[6], w698, w699);
  FullAdder U75 (w699, w684, IN12[5], w700, w701);
  FullAdder U76 (w701, w686, IN13[4], w702, w703);
  FullAdder U77 (w703, w688, IN14[3], w704, w705);
  FullAdder U78 (w705, w690, IN15[2], w706, w707);
  FullAdder U79 (w707, w692, IN16[1], w708, w709);
  FullAdder U80 (w709, w693, IN17[0], w710, w711);
  HalfAdder U81 (w696, IN10[8], Out1[10], w713);
  FullAdder U82 (w713, w698, IN11[7], w714, w715);
  FullAdder U83 (w715, w700, IN12[6], w716, w717);
  FullAdder U84 (w717, w702, IN13[5], w718, w719);
  FullAdder U85 (w719, w704, IN14[4], w720, w721);
  FullAdder U86 (w721, w706, IN15[3], w722, w723);
  FullAdder U87 (w723, w708, IN16[2], w724, w725);
  FullAdder U88 (w725, w710, IN17[1], w726, w727);
  FullAdder U89 (w727, w711, IN18[0], w728, w729);
  HalfAdder U90 (w714, IN11[8], Out1[11], w731);
  FullAdder U91 (w731, w716, IN12[7], w732, w733);
  FullAdder U92 (w733, w718, IN13[6], w734, w735);
  FullAdder U93 (w735, w720, IN14[5], w736, w737);
  FullAdder U94 (w737, w722, IN15[4], w738, w739);
  FullAdder U95 (w739, w724, IN16[3], w740, w741);
  FullAdder U96 (w741, w726, IN17[2], w742, w743);
  FullAdder U97 (w743, w728, IN18[1], w744, w745);
  FullAdder U98 (w745, w729, IN19[0], w746, w747);
  HalfAdder U99 (w732, IN12[8], Out1[12], w749);
  FullAdder U100 (w749, w734, IN13[7], w750, w751);
  FullAdder U101 (w751, w736, IN14[6], w752, w753);
  FullAdder U102 (w753, w738, IN15[5], w754, w755);
  FullAdder U103 (w755, w740, IN16[4], w756, w757);
  FullAdder U104 (w757, w742, IN17[3], w758, w759);
  FullAdder U105 (w759, w744, IN18[2], w760, w761);
  FullAdder U106 (w761, w746, IN19[1], w762, w763);
  FullAdder U107 (w763, w747, IN20[0], w764, w765);
  HalfAdder U108 (w750, IN13[8], Out1[13], w767);
  FullAdder U109 (w767, w752, IN14[7], w768, w769);
  FullAdder U110 (w769, w754, IN15[6], w770, w771);
  FullAdder U111 (w771, w756, IN16[5], w772, w773);
  FullAdder U112 (w773, w758, IN17[4], w774, w775);
  FullAdder U113 (w775, w760, IN18[3], w776, w777);
  FullAdder U114 (w777, w762, IN19[2], w778, w779);
  FullAdder U115 (w779, w764, IN20[1], w780, w781);
  FullAdder U116 (w781, w765, IN21[0], w782, w783);
  HalfAdder U117 (w768, IN14[8], Out1[14], w785);
  FullAdder U118 (w785, w770, IN15[7], w786, w787);
  FullAdder U119 (w787, w772, IN16[6], w788, w789);
  FullAdder U120 (w789, w774, IN17[5], w790, w791);
  FullAdder U121 (w791, w776, IN18[4], w792, w793);
  FullAdder U122 (w793, w778, IN19[3], w794, w795);
  FullAdder U123 (w795, w780, IN20[2], w796, w797);
  FullAdder U124 (w797, w782, IN21[1], w798, w799);
  FullAdder U125 (w799, w783, IN22[0], w800, w801);
  HalfAdder U126 (w786, IN15[8], Out1[15], w803);
  FullAdder U127 (w803, w788, IN16[7], w804, w805);
  FullAdder U128 (w805, w790, IN17[6], w806, w807);
  FullAdder U129 (w807, w792, IN18[5], w808, w809);
  FullAdder U130 (w809, w794, IN19[4], w810, w811);
  FullAdder U131 (w811, w796, IN20[3], w812, w813);
  FullAdder U132 (w813, w798, IN21[2], w814, w815);
  FullAdder U133 (w815, w800, IN22[1], w816, w817);
  FullAdder U134 (w817, w801, IN23[0], w818, w819);
  HalfAdder U135 (w804, IN16[8], Out1[16], w821);
  FullAdder U136 (w821, w806, IN17[7], w822, w823);
  FullAdder U137 (w823, w808, IN18[6], w824, w825);
  FullAdder U138 (w825, w810, IN19[5], w826, w827);
  FullAdder U139 (w827, w812, IN20[4], w828, w829);
  FullAdder U140 (w829, w814, IN21[3], w830, w831);
  FullAdder U141 (w831, w816, IN22[2], w832, w833);
  FullAdder U142 (w833, w818, IN23[1], w834, w835);
  FullAdder U143 (w835, w819, IN24[0], w836, w837);
  HalfAdder U144 (w822, IN17[8], Out1[17], w839);
  FullAdder U145 (w839, w824, IN18[7], w840, w841);
  FullAdder U146 (w841, w826, IN19[6], w842, w843);
  FullAdder U147 (w843, w828, IN20[5], w844, w845);
  FullAdder U148 (w845, w830, IN21[4], w846, w847);
  FullAdder U149 (w847, w832, IN22[3], w848, w849);
  FullAdder U150 (w849, w834, IN23[2], w850, w851);
  FullAdder U151 (w851, w836, IN24[1], w852, w853);
  FullAdder U152 (w853, w837, IN25[0], w854, w855);
  HalfAdder U153 (w840, IN18[8], Out1[18], w857);
  FullAdder U154 (w857, w842, IN19[7], w858, w859);
  FullAdder U155 (w859, w844, IN20[6], w860, w861);
  FullAdder U156 (w861, w846, IN21[5], w862, w863);
  FullAdder U157 (w863, w848, IN22[4], w864, w865);
  FullAdder U158 (w865, w850, IN23[3], w866, w867);
  FullAdder U159 (w867, w852, IN24[2], w868, w869);
  FullAdder U160 (w869, w854, IN25[1], w870, w871);
  FullAdder U161 (w871, w855, IN26[0], w872, w873);
  HalfAdder U162 (w858, IN19[8], Out1[19], w875);
  FullAdder U163 (w875, w860, IN20[7], w876, w877);
  FullAdder U164 (w877, w862, IN21[6], w878, w879);
  FullAdder U165 (w879, w864, IN22[5], w880, w881);
  FullAdder U166 (w881, w866, IN23[4], w882, w883);
  FullAdder U167 (w883, w868, IN24[3], w884, w885);
  FullAdder U168 (w885, w870, IN25[2], w886, w887);
  FullAdder U169 (w887, w872, IN26[1], w888, w889);
  FullAdder U170 (w889, w873, IN27[0], w890, w891);
  HalfAdder U171 (w876, IN20[8], Out1[20], w893);
  FullAdder U172 (w893, w878, IN21[7], w894, w895);
  FullAdder U173 (w895, w880, IN22[6], w896, w897);
  FullAdder U174 (w897, w882, IN23[5], w898, w899);
  FullAdder U175 (w899, w884, IN24[4], w900, w901);
  FullAdder U176 (w901, w886, IN25[3], w902, w903);
  FullAdder U177 (w903, w888, IN26[2], w904, w905);
  FullAdder U178 (w905, w890, IN27[1], w906, w907);
  FullAdder U179 (w907, w891, IN28[0], w908, w909);
  HalfAdder U180 (w894, IN21[8], Out1[21], w911);
  FullAdder U181 (w911, w896, IN22[7], w912, w913);
  FullAdder U182 (w913, w898, IN23[6], w914, w915);
  FullAdder U183 (w915, w900, IN24[5], w916, w917);
  FullAdder U184 (w917, w902, IN25[4], w918, w919);
  FullAdder U185 (w919, w904, IN26[3], w920, w921);
  FullAdder U186 (w921, w906, IN27[2], w922, w923);
  FullAdder U187 (w923, w908, IN28[1], w924, w925);
  FullAdder U188 (w925, w909, IN29[0], w926, w927);
  HalfAdder U189 (w912, IN22[8], Out1[22], w929);
  FullAdder U190 (w929, w914, IN23[7], w930, w931);
  FullAdder U191 (w931, w916, IN24[6], w932, w933);
  FullAdder U192 (w933, w918, IN25[5], w934, w935);
  FullAdder U193 (w935, w920, IN26[4], w936, w937);
  FullAdder U194 (w937, w922, IN27[3], w938, w939);
  FullAdder U195 (w939, w924, IN28[2], w940, w941);
  FullAdder U196 (w941, w926, IN29[1], w942, w943);
  FullAdder U197 (w943, w927, IN30[0], w944, w945);
  HalfAdder U198 (w930, IN23[8], Out1[23], w947);
  FullAdder U199 (w947, w932, IN24[7], w948, w949);
  FullAdder U200 (w949, w934, IN25[6], w950, w951);
  FullAdder U201 (w951, w936, IN26[5], w952, w953);
  FullAdder U202 (w953, w938, IN27[4], w954, w955);
  FullAdder U203 (w955, w940, IN28[3], w956, w957);
  FullAdder U204 (w957, w942, IN29[2], w958, w959);
  FullAdder U205 (w959, w944, IN30[1], w960, w961);
  FullAdder U206 (w961, w945, IN31[0], w962, w963);
  HalfAdder U207 (w948, IN24[8], Out1[24], w965);
  FullAdder U208 (w965, w950, IN25[7], w966, w967);
  FullAdder U209 (w967, w952, IN26[6], w968, w969);
  FullAdder U210 (w969, w954, IN27[5], w970, w971);
  FullAdder U211 (w971, w956, IN28[4], w972, w973);
  FullAdder U212 (w973, w958, IN29[3], w974, w975);
  FullAdder U213 (w975, w960, IN30[2], w976, w977);
  FullAdder U214 (w977, w962, IN31[1], w978, w979);
  FullAdder U215 (w979, w963, IN32[0], w980, w981);
  HalfAdder U216 (w966, IN25[8], Out1[25], w983);
  FullAdder U217 (w983, w968, IN26[7], w984, w985);
  FullAdder U218 (w985, w970, IN27[6], w986, w987);
  FullAdder U219 (w987, w972, IN28[5], w988, w989);
  FullAdder U220 (w989, w974, IN29[4], w990, w991);
  FullAdder U221 (w991, w976, IN30[3], w992, w993);
  FullAdder U222 (w993, w978, IN31[2], w994, w995);
  FullAdder U223 (w995, w980, IN32[1], w996, w997);
  FullAdder U224 (w997, w981, IN33[0], w998, w999);
  HalfAdder U225 (w984, IN26[8], Out1[26], w1001);
  FullAdder U226 (w1001, w986, IN27[7], w1002, w1003);
  FullAdder U227 (w1003, w988, IN28[6], w1004, w1005);
  FullAdder U228 (w1005, w990, IN29[5], w1006, w1007);
  FullAdder U229 (w1007, w992, IN30[4], w1008, w1009);
  FullAdder U230 (w1009, w994, IN31[3], w1010, w1011);
  FullAdder U231 (w1011, w996, IN32[2], w1012, w1013);
  FullAdder U232 (w1013, w998, IN33[1], w1014, w1015);
  FullAdder U233 (w1015, w999, IN34[0], w1016, w1017);
  HalfAdder U234 (w1002, IN27[8], Out1[27], w1019);
  FullAdder U235 (w1019, w1004, IN28[7], w1020, w1021);
  FullAdder U236 (w1021, w1006, IN29[6], w1022, w1023);
  FullAdder U237 (w1023, w1008, IN30[5], w1024, w1025);
  FullAdder U238 (w1025, w1010, IN31[4], w1026, w1027);
  FullAdder U239 (w1027, w1012, IN32[3], w1028, w1029);
  FullAdder U240 (w1029, w1014, IN33[2], w1030, w1031);
  FullAdder U241 (w1031, w1016, IN34[1], w1032, w1033);
  FullAdder U242 (w1033, w1017, IN35[0], w1034, w1035);
  HalfAdder U243 (w1020, IN28[8], Out1[28], w1037);
  FullAdder U244 (w1037, w1022, IN29[7], w1038, w1039);
  FullAdder U245 (w1039, w1024, IN30[6], w1040, w1041);
  FullAdder U246 (w1041, w1026, IN31[5], w1042, w1043);
  FullAdder U247 (w1043, w1028, IN32[4], w1044, w1045);
  FullAdder U248 (w1045, w1030, IN33[3], w1046, w1047);
  FullAdder U249 (w1047, w1032, IN34[2], w1048, w1049);
  FullAdder U250 (w1049, w1034, IN35[1], w1050, w1051);
  FullAdder U251 (w1051, w1035, IN36[0], w1052, w1053);
  HalfAdder U252 (w1038, IN29[8], Out1[29], w1055);
  FullAdder U253 (w1055, w1040, IN30[7], w1056, w1057);
  FullAdder U254 (w1057, w1042, IN31[6], w1058, w1059);
  FullAdder U255 (w1059, w1044, IN32[5], w1060, w1061);
  FullAdder U256 (w1061, w1046, IN33[4], w1062, w1063);
  FullAdder U257 (w1063, w1048, IN34[3], w1064, w1065);
  FullAdder U258 (w1065, w1050, IN35[2], w1066, w1067);
  FullAdder U259 (w1067, w1052, IN36[1], w1068, w1069);
  FullAdder U260 (w1069, w1053, IN37[0], w1070, w1071);
  HalfAdder U261 (w1056, IN30[8], Out1[30], w1073);
  FullAdder U262 (w1073, w1058, IN31[7], w1074, w1075);
  FullAdder U263 (w1075, w1060, IN32[6], w1076, w1077);
  FullAdder U264 (w1077, w1062, IN33[5], w1078, w1079);
  FullAdder U265 (w1079, w1064, IN34[4], w1080, w1081);
  FullAdder U266 (w1081, w1066, IN35[3], w1082, w1083);
  FullAdder U267 (w1083, w1068, IN36[2], w1084, w1085);
  FullAdder U268 (w1085, w1070, IN37[1], w1086, w1087);
  FullAdder U269 (w1087, w1071, IN38[0], w1088, w1089);
  HalfAdder U270 (w1074, IN31[8], Out1[31], w1091);
  FullAdder U271 (w1091, w1076, IN32[7], w1092, w1093);
  FullAdder U272 (w1093, w1078, IN33[6], w1094, w1095);
  FullAdder U273 (w1095, w1080, IN34[5], w1096, w1097);
  FullAdder U274 (w1097, w1082, IN35[4], w1098, w1099);
  FullAdder U275 (w1099, w1084, IN36[3], w1100, w1101);
  FullAdder U276 (w1101, w1086, IN37[2], w1102, w1103);
  FullAdder U277 (w1103, w1088, IN38[1], w1104, w1105);
  FullAdder U278 (w1105, w1089, IN39[0], w1106, w1107);
  HalfAdder U279 (w1092, IN32[8], Out1[32], w1109);
  FullAdder U280 (w1109, w1094, IN33[7], w1110, w1111);
  FullAdder U281 (w1111, w1096, IN34[6], w1112, w1113);
  FullAdder U282 (w1113, w1098, IN35[5], w1114, w1115);
  FullAdder U283 (w1115, w1100, IN36[4], w1116, w1117);
  FullAdder U284 (w1117, w1102, IN37[3], w1118, w1119);
  FullAdder U285 (w1119, w1104, IN38[2], w1120, w1121);
  FullAdder U286 (w1121, w1106, IN39[1], w1122, w1123);
  FullAdder U287 (w1123, w1107, IN40[0], w1124, w1125);
  HalfAdder U288 (w1110, IN33[8], Out1[33], w1127);
  FullAdder U289 (w1127, w1112, IN34[7], w1128, w1129);
  FullAdder U290 (w1129, w1114, IN35[6], w1130, w1131);
  FullAdder U291 (w1131, w1116, IN36[5], w1132, w1133);
  FullAdder U292 (w1133, w1118, IN37[4], w1134, w1135);
  FullAdder U293 (w1135, w1120, IN38[3], w1136, w1137);
  FullAdder U294 (w1137, w1122, IN39[2], w1138, w1139);
  FullAdder U295 (w1139, w1124, IN40[1], w1140, w1141);
  FullAdder U296 (w1141, w1125, IN41[0], w1142, w1143);
  HalfAdder U297 (w1128, IN34[8], Out1[34], w1145);
  FullAdder U298 (w1145, w1130, IN35[7], w1146, w1147);
  FullAdder U299 (w1147, w1132, IN36[6], w1148, w1149);
  FullAdder U300 (w1149, w1134, IN37[5], w1150, w1151);
  FullAdder U301 (w1151, w1136, IN38[4], w1152, w1153);
  FullAdder U302 (w1153, w1138, IN39[3], w1154, w1155);
  FullAdder U303 (w1155, w1140, IN40[2], w1156, w1157);
  FullAdder U304 (w1157, w1142, IN41[1], w1158, w1159);
  FullAdder U305 (w1159, w1143, IN42[0], w1160, w1161);
  HalfAdder U306 (w1146, IN35[8], Out1[35], w1163);
  FullAdder U307 (w1163, w1148, IN36[7], w1164, w1165);
  FullAdder U308 (w1165, w1150, IN37[6], w1166, w1167);
  FullAdder U309 (w1167, w1152, IN38[5], w1168, w1169);
  FullAdder U310 (w1169, w1154, IN39[4], w1170, w1171);
  FullAdder U311 (w1171, w1156, IN40[3], w1172, w1173);
  FullAdder U312 (w1173, w1158, IN41[2], w1174, w1175);
  FullAdder U313 (w1175, w1160, IN42[1], w1176, w1177);
  FullAdder U314 (w1177, w1161, IN43[0], w1178, w1179);
  HalfAdder U315 (w1164, IN36[8], Out1[36], w1181);
  FullAdder U316 (w1181, w1166, IN37[7], w1182, w1183);
  FullAdder U317 (w1183, w1168, IN38[6], w1184, w1185);
  FullAdder U318 (w1185, w1170, IN39[5], w1186, w1187);
  FullAdder U319 (w1187, w1172, IN40[4], w1188, w1189);
  FullAdder U320 (w1189, w1174, IN41[3], w1190, w1191);
  FullAdder U321 (w1191, w1176, IN42[2], w1192, w1193);
  FullAdder U322 (w1193, w1178, IN43[1], w1194, w1195);
  FullAdder U323 (w1195, w1179, IN44[0], w1196, w1197);
  HalfAdder U324 (w1182, IN37[8], Out1[37], w1199);
  FullAdder U325 (w1199, w1184, IN38[7], w1200, w1201);
  FullAdder U326 (w1201, w1186, IN39[6], w1202, w1203);
  FullAdder U327 (w1203, w1188, IN40[5], w1204, w1205);
  FullAdder U328 (w1205, w1190, IN41[4], w1206, w1207);
  FullAdder U329 (w1207, w1192, IN42[3], w1208, w1209);
  FullAdder U330 (w1209, w1194, IN43[2], w1210, w1211);
  FullAdder U331 (w1211, w1196, IN44[1], w1212, w1213);
  FullAdder U332 (w1213, w1197, IN45[0], w1214, w1215);
  HalfAdder U333 (w1200, IN38[8], Out1[38], w1217);
  FullAdder U334 (w1217, w1202, IN39[7], w1218, w1219);
  FullAdder U335 (w1219, w1204, IN40[6], w1220, w1221);
  FullAdder U336 (w1221, w1206, IN41[5], w1222, w1223);
  FullAdder U337 (w1223, w1208, IN42[4], w1224, w1225);
  FullAdder U338 (w1225, w1210, IN43[3], w1226, w1227);
  FullAdder U339 (w1227, w1212, IN44[2], w1228, w1229);
  FullAdder U340 (w1229, w1214, IN45[1], w1230, w1231);
  FullAdder U341 (w1231, w1215, IN46[0], w1232, w1233);
  HalfAdder U342 (w1218, IN39[8], Out1[39], w1235);
  FullAdder U343 (w1235, w1220, IN40[7], w1236, w1237);
  FullAdder U344 (w1237, w1222, IN41[6], w1238, w1239);
  FullAdder U345 (w1239, w1224, IN42[5], w1240, w1241);
  FullAdder U346 (w1241, w1226, IN43[4], w1242, w1243);
  FullAdder U347 (w1243, w1228, IN44[3], w1244, w1245);
  FullAdder U348 (w1245, w1230, IN45[2], w1246, w1247);
  FullAdder U349 (w1247, w1232, IN46[1], w1248, w1249);
  FullAdder U350 (w1249, w1233, IN47[0], w1250, w1251);
  HalfAdder U351 (w1236, IN40[8], Out1[40], w1253);
  FullAdder U352 (w1253, w1238, IN41[7], w1254, w1255);
  FullAdder U353 (w1255, w1240, IN42[6], w1256, w1257);
  FullAdder U354 (w1257, w1242, IN43[5], w1258, w1259);
  FullAdder U355 (w1259, w1244, IN44[4], w1260, w1261);
  FullAdder U356 (w1261, w1246, IN45[3], w1262, w1263);
  FullAdder U357 (w1263, w1248, IN46[2], w1264, w1265);
  FullAdder U358 (w1265, w1250, IN47[1], w1266, w1267);
  FullAdder U359 (w1267, w1251, IN48[0], w1268, w1269);
  HalfAdder U360 (w1254, IN41[8], Out1[41], w1271);
  FullAdder U361 (w1271, w1256, IN42[7], w1272, w1273);
  FullAdder U362 (w1273, w1258, IN43[6], w1274, w1275);
  FullAdder U363 (w1275, w1260, IN44[5], w1276, w1277);
  FullAdder U364 (w1277, w1262, IN45[4], w1278, w1279);
  FullAdder U365 (w1279, w1264, IN46[3], w1280, w1281);
  FullAdder U366 (w1281, w1266, IN47[2], w1282, w1283);
  FullAdder U367 (w1283, w1268, IN48[1], w1284, w1285);
  FullAdder U368 (w1285, w1269, IN49[0], w1286, w1287);
  HalfAdder U369 (w1272, IN42[8], Out1[42], w1289);
  FullAdder U370 (w1289, w1274, IN43[7], w1290, w1291);
  FullAdder U371 (w1291, w1276, IN44[6], w1292, w1293);
  FullAdder U372 (w1293, w1278, IN45[5], w1294, w1295);
  FullAdder U373 (w1295, w1280, IN46[4], w1296, w1297);
  FullAdder U374 (w1297, w1282, IN47[3], w1298, w1299);
  FullAdder U375 (w1299, w1284, IN48[2], w1300, w1301);
  FullAdder U376 (w1301, w1286, IN49[1], w1302, w1303);
  FullAdder U377 (w1303, w1287, IN50[0], w1304, w1305);
  HalfAdder U378 (w1290, IN43[8], Out1[43], w1307);
  FullAdder U379 (w1307, w1292, IN44[7], w1308, w1309);
  FullAdder U380 (w1309, w1294, IN45[6], w1310, w1311);
  FullAdder U381 (w1311, w1296, IN46[5], w1312, w1313);
  FullAdder U382 (w1313, w1298, IN47[4], w1314, w1315);
  FullAdder U383 (w1315, w1300, IN48[3], w1316, w1317);
  FullAdder U384 (w1317, w1302, IN49[2], w1318, w1319);
  FullAdder U385 (w1319, w1304, IN50[1], w1320, w1321);
  FullAdder U386 (w1321, w1305, IN51[0], w1322, w1323);
  HalfAdder U387 (w1308, IN44[8], Out1[44], w1325);
  FullAdder U388 (w1325, w1310, IN45[7], w1326, w1327);
  FullAdder U389 (w1327, w1312, IN46[6], w1328, w1329);
  FullAdder U390 (w1329, w1314, IN47[5], w1330, w1331);
  FullAdder U391 (w1331, w1316, IN48[4], w1332, w1333);
  FullAdder U392 (w1333, w1318, IN49[3], w1334, w1335);
  FullAdder U393 (w1335, w1320, IN50[2], w1336, w1337);
  FullAdder U394 (w1337, w1322, IN51[1], w1338, w1339);
  FullAdder U395 (w1339, w1323, IN52[0], w1340, w1341);
  HalfAdder U396 (w1326, IN45[8], Out1[45], w1343);
  FullAdder U397 (w1343, w1328, IN46[7], w1344, w1345);
  FullAdder U398 (w1345, w1330, IN47[6], w1346, w1347);
  FullAdder U399 (w1347, w1332, IN48[5], w1348, w1349);
  FullAdder U400 (w1349, w1334, IN49[4], w1350, w1351);
  FullAdder U401 (w1351, w1336, IN50[3], w1352, w1353);
  FullAdder U402 (w1353, w1338, IN51[2], w1354, w1355);
  FullAdder U403 (w1355, w1340, IN52[1], w1356, w1357);
  FullAdder U404 (w1357, w1341, IN53[0], w1358, w1359);
  HalfAdder U405 (w1344, IN46[8], Out1[46], w1361);
  FullAdder U406 (w1361, w1346, IN47[7], w1362, w1363);
  FullAdder U407 (w1363, w1348, IN48[6], w1364, w1365);
  FullAdder U408 (w1365, w1350, IN49[5], w1366, w1367);
  FullAdder U409 (w1367, w1352, IN50[4], w1368, w1369);
  FullAdder U410 (w1369, w1354, IN51[3], w1370, w1371);
  FullAdder U411 (w1371, w1356, IN52[2], w1372, w1373);
  FullAdder U412 (w1373, w1358, IN53[1], w1374, w1375);
  FullAdder U413 (w1375, w1359, IN54[0], w1376, w1377);
  HalfAdder U414 (w1362, IN47[8], Out1[47], w1379);
  FullAdder U415 (w1379, w1364, IN48[7], w1380, w1381);
  FullAdder U416 (w1381, w1366, IN49[6], w1382, w1383);
  FullAdder U417 (w1383, w1368, IN50[5], w1384, w1385);
  FullAdder U418 (w1385, w1370, IN51[4], w1386, w1387);
  FullAdder U419 (w1387, w1372, IN52[3], w1388, w1389);
  FullAdder U420 (w1389, w1374, IN53[2], w1390, w1391);
  FullAdder U421 (w1391, w1376, IN54[1], w1392, w1393);
  FullAdder U422 (w1393, w1377, IN55[0], w1394, w1395);
  HalfAdder U423 (w1380, IN48[8], Out1[48], w1397);
  FullAdder U424 (w1397, w1382, IN49[7], w1398, w1399);
  FullAdder U425 (w1399, w1384, IN50[6], w1400, w1401);
  FullAdder U426 (w1401, w1386, IN51[5], w1402, w1403);
  FullAdder U427 (w1403, w1388, IN52[4], w1404, w1405);
  FullAdder U428 (w1405, w1390, IN53[3], w1406, w1407);
  FullAdder U429 (w1407, w1392, IN54[2], w1408, w1409);
  FullAdder U430 (w1409, w1394, IN55[1], w1410, w1411);
  FullAdder U431 (w1411, w1395, IN56[0], w1412, w1413);
  HalfAdder U432 (w1398, IN49[8], Out1[49], w1415);
  FullAdder U433 (w1415, w1400, IN50[7], w1416, w1417);
  FullAdder U434 (w1417, w1402, IN51[6], w1418, w1419);
  FullAdder U435 (w1419, w1404, IN52[5], w1420, w1421);
  FullAdder U436 (w1421, w1406, IN53[4], w1422, w1423);
  FullAdder U437 (w1423, w1408, IN54[3], w1424, w1425);
  FullAdder U438 (w1425, w1410, IN55[2], w1426, w1427);
  FullAdder U439 (w1427, w1412, IN56[1], w1428, w1429);
  FullAdder U440 (w1429, w1413, IN57[0], w1430, w1431);
  HalfAdder U441 (w1416, IN50[8], Out1[50], w1433);
  FullAdder U442 (w1433, w1418, IN51[7], w1434, w1435);
  FullAdder U443 (w1435, w1420, IN52[6], w1436, w1437);
  FullAdder U444 (w1437, w1422, IN53[5], w1438, w1439);
  FullAdder U445 (w1439, w1424, IN54[4], w1440, w1441);
  FullAdder U446 (w1441, w1426, IN55[3], w1442, w1443);
  FullAdder U447 (w1443, w1428, IN56[2], w1444, w1445);
  FullAdder U448 (w1445, w1430, IN57[1], w1446, w1447);
  FullAdder U449 (w1447, w1431, IN58[0], w1448, w1449);
  HalfAdder U450 (w1434, IN51[8], Out1[51], w1451);
  FullAdder U451 (w1451, w1436, IN52[7], w1452, w1453);
  FullAdder U452 (w1453, w1438, IN53[6], w1454, w1455);
  FullAdder U453 (w1455, w1440, IN54[5], w1456, w1457);
  FullAdder U454 (w1457, w1442, IN55[4], w1458, w1459);
  FullAdder U455 (w1459, w1444, IN56[3], w1460, w1461);
  FullAdder U456 (w1461, w1446, IN57[2], w1462, w1463);
  FullAdder U457 (w1463, w1448, IN58[1], w1464, w1465);
  FullAdder U458 (w1465, w1449, IN59[0], w1466, w1467);
  HalfAdder U459 (w1452, IN52[8], Out1[52], w1469);
  FullAdder U460 (w1469, w1454, IN53[7], w1470, w1471);
  FullAdder U461 (w1471, w1456, IN54[6], w1472, w1473);
  FullAdder U462 (w1473, w1458, IN55[5], w1474, w1475);
  FullAdder U463 (w1475, w1460, IN56[4], w1476, w1477);
  FullAdder U464 (w1477, w1462, IN57[3], w1478, w1479);
  FullAdder U465 (w1479, w1464, IN58[2], w1480, w1481);
  FullAdder U466 (w1481, w1466, IN59[1], w1482, w1483);
  FullAdder U467 (w1483, w1467, IN60[0], w1484, w1485);
  HalfAdder U468 (w1470, IN53[8], Out1[53], w1487);
  FullAdder U469 (w1487, w1472, IN54[7], w1488, w1489);
  FullAdder U470 (w1489, w1474, IN55[6], w1490, w1491);
  FullAdder U471 (w1491, w1476, IN56[5], w1492, w1493);
  FullAdder U472 (w1493, w1478, IN57[4], w1494, w1495);
  FullAdder U473 (w1495, w1480, IN58[3], w1496, w1497);
  FullAdder U474 (w1497, w1482, IN59[2], w1498, w1499);
  FullAdder U475 (w1499, w1484, IN60[1], w1500, w1501);
  FullAdder U476 (w1501, w1485, IN61[0], w1502, w1503);
  HalfAdder U477 (w1488, IN54[8], Out1[54], w1505);
  FullAdder U478 (w1505, w1490, IN55[7], Out1[55], w1507);
  FullAdder U479 (w1507, w1492, IN56[6], Out1[56], w1509);
  FullAdder U480 (w1509, w1494, IN57[5], Out1[57], w1511);
  FullAdder U481 (w1511, w1496, IN58[4], Out1[58], w1513);
  FullAdder U482 (w1513, w1498, IN59[3], Out1[59], w1515);
  FullAdder U483 (w1515, w1500, IN60[2], Out1[60], w1517);
  FullAdder U484 (w1517, w1502, IN61[1], Out1[61], w1519);
  FullAdder U485 (w1519, w1503, IN62[0], Out1[62], Out1[63]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN10[9];
  assign Out2[1] = IN11[9];
  assign Out2[2] = IN12[9];
  assign Out2[3] = IN13[9];
  assign Out2[4] = IN14[9];
  assign Out2[5] = IN15[9];
  assign Out2[6] = IN16[9];
  assign Out2[7] = IN17[9];
  assign Out2[8] = IN18[9];
  assign Out2[9] = IN19[9];
  assign Out2[10] = IN20[9];
  assign Out2[11] = IN21[9];
  assign Out2[12] = IN22[9];
  assign Out2[13] = IN23[9];
  assign Out2[14] = IN24[9];
  assign Out2[15] = IN25[9];
  assign Out2[16] = IN26[9];
  assign Out2[17] = IN27[9];
  assign Out2[18] = IN28[9];
  assign Out2[19] = IN29[9];
  assign Out2[20] = IN30[9];
  assign Out2[21] = IN31[9];
  assign Out2[22] = IN32[9];
  assign Out2[23] = IN33[9];
  assign Out2[24] = IN34[9];
  assign Out2[25] = IN35[9];
  assign Out2[26] = IN36[9];
  assign Out2[27] = IN37[9];
  assign Out2[28] = IN38[9];
  assign Out2[29] = IN39[9];
  assign Out2[30] = IN40[9];
  assign Out2[31] = IN41[9];
  assign Out2[32] = IN42[9];
  assign Out2[33] = IN43[9];
  assign Out2[34] = IN44[9];
  assign Out2[35] = IN45[9];
  assign Out2[36] = IN46[9];
  assign Out2[37] = IN47[9];
  assign Out2[38] = IN48[9];
  assign Out2[39] = IN49[9];
  assign Out2[40] = IN50[9];
  assign Out2[41] = IN51[9];
  assign Out2[42] = IN52[9];
  assign Out2[43] = IN53[9];
  assign Out2[44] = IN54[9];
  assign Out2[45] = IN55[8];
  assign Out2[46] = IN56[7];
  assign Out2[47] = IN57[6];
  assign Out2[48] = IN58[5];
  assign Out2[49] = IN59[4];
  assign Out2[50] = IN60[3];
  assign Out2[51] = IN61[2];
  assign Out2[52] = IN62[1];
  assign Out2[53] = IN63[0];

endmodule
module RC_54_54(IN1, IN2, Out);
  input [53:0] IN1;
  input [53:0] IN2;
  output [54:0] Out;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w109);
  FullAdder U1 (IN1[1], IN2[1], w109, Out[1], w111);
  FullAdder U2 (IN1[2], IN2[2], w111, Out[2], w113);
  FullAdder U3 (IN1[3], IN2[3], w113, Out[3], w115);
  FullAdder U4 (IN1[4], IN2[4], w115, Out[4], w117);
  FullAdder U5 (IN1[5], IN2[5], w117, Out[5], w119);
  FullAdder U6 (IN1[6], IN2[6], w119, Out[6], w121);
  FullAdder U7 (IN1[7], IN2[7], w121, Out[7], w123);
  FullAdder U8 (IN1[8], IN2[8], w123, Out[8], w125);
  FullAdder U9 (IN1[9], IN2[9], w125, Out[9], w127);
  FullAdder U10 (IN1[10], IN2[10], w127, Out[10], w129);
  FullAdder U11 (IN1[11], IN2[11], w129, Out[11], w131);
  FullAdder U12 (IN1[12], IN2[12], w131, Out[12], w133);
  FullAdder U13 (IN1[13], IN2[13], w133, Out[13], w135);
  FullAdder U14 (IN1[14], IN2[14], w135, Out[14], w137);
  FullAdder U15 (IN1[15], IN2[15], w137, Out[15], w139);
  FullAdder U16 (IN1[16], IN2[16], w139, Out[16], w141);
  FullAdder U17 (IN1[17], IN2[17], w141, Out[17], w143);
  FullAdder U18 (IN1[18], IN2[18], w143, Out[18], w145);
  FullAdder U19 (IN1[19], IN2[19], w145, Out[19], w147);
  FullAdder U20 (IN1[20], IN2[20], w147, Out[20], w149);
  FullAdder U21 (IN1[21], IN2[21], w149, Out[21], w151);
  FullAdder U22 (IN1[22], IN2[22], w151, Out[22], w153);
  FullAdder U23 (IN1[23], IN2[23], w153, Out[23], w155);
  FullAdder U24 (IN1[24], IN2[24], w155, Out[24], w157);
  FullAdder U25 (IN1[25], IN2[25], w157, Out[25], w159);
  FullAdder U26 (IN1[26], IN2[26], w159, Out[26], w161);
  FullAdder U27 (IN1[27], IN2[27], w161, Out[27], w163);
  FullAdder U28 (IN1[28], IN2[28], w163, Out[28], w165);
  FullAdder U29 (IN1[29], IN2[29], w165, Out[29], w167);
  FullAdder U30 (IN1[30], IN2[30], w167, Out[30], w169);
  FullAdder U31 (IN1[31], IN2[31], w169, Out[31], w171);
  FullAdder U32 (IN1[32], IN2[32], w171, Out[32], w173);
  FullAdder U33 (IN1[33], IN2[33], w173, Out[33], w175);
  FullAdder U34 (IN1[34], IN2[34], w175, Out[34], w177);
  FullAdder U35 (IN1[35], IN2[35], w177, Out[35], w179);
  FullAdder U36 (IN1[36], IN2[36], w179, Out[36], w181);
  FullAdder U37 (IN1[37], IN2[37], w181, Out[37], w183);
  FullAdder U38 (IN1[38], IN2[38], w183, Out[38], w185);
  FullAdder U39 (IN1[39], IN2[39], w185, Out[39], w187);
  FullAdder U40 (IN1[40], IN2[40], w187, Out[40], w189);
  FullAdder U41 (IN1[41], IN2[41], w189, Out[41], w191);
  FullAdder U42 (IN1[42], IN2[42], w191, Out[42], w193);
  FullAdder U43 (IN1[43], IN2[43], w193, Out[43], w195);
  FullAdder U44 (IN1[44], IN2[44], w195, Out[44], w197);
  FullAdder U45 (IN1[45], IN2[45], w197, Out[45], w199);
  FullAdder U46 (IN1[46], IN2[46], w199, Out[46], w201);
  FullAdder U47 (IN1[47], IN2[47], w201, Out[47], w203);
  FullAdder U48 (IN1[48], IN2[48], w203, Out[48], w205);
  FullAdder U49 (IN1[49], IN2[49], w205, Out[49], w207);
  FullAdder U50 (IN1[50], IN2[50], w207, Out[50], w209);
  FullAdder U51 (IN1[51], IN2[51], w209, Out[51], w211);
  FullAdder U52 (IN1[52], IN2[52], w211, Out[52], w213);
  FullAdder U53 (IN1[53], IN2[53], w213, Out[53], Out[54]);

endmodule
module NR_10_55(IN1, IN2, Out);
  input [9:0] IN1;
  input [54:0] IN2;
  output [64:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [9:0] P10;
  wire [9:0] P11;
  wire [9:0] P12;
  wire [9:0] P13;
  wire [9:0] P14;
  wire [9:0] P15;
  wire [9:0] P16;
  wire [9:0] P17;
  wire [9:0] P18;
  wire [9:0] P19;
  wire [9:0] P20;
  wire [9:0] P21;
  wire [9:0] P22;
  wire [9:0] P23;
  wire [9:0] P24;
  wire [9:0] P25;
  wire [9:0] P26;
  wire [9:0] P27;
  wire [9:0] P28;
  wire [9:0] P29;
  wire [9:0] P30;
  wire [9:0] P31;
  wire [9:0] P32;
  wire [9:0] P33;
  wire [9:0] P34;
  wire [9:0] P35;
  wire [9:0] P36;
  wire [9:0] P37;
  wire [9:0] P38;
  wire [9:0] P39;
  wire [9:0] P40;
  wire [9:0] P41;
  wire [9:0] P42;
  wire [9:0] P43;
  wire [9:0] P44;
  wire [9:0] P45;
  wire [9:0] P46;
  wire [9:0] P47;
  wire [9:0] P48;
  wire [9:0] P49;
  wire [9:0] P50;
  wire [9:0] P51;
  wire [9:0] P52;
  wire [9:0] P53;
  wire [9:0] P54;
  wire [8:0] P55;
  wire [7:0] P56;
  wire [6:0] P57;
  wire [5:0] P58;
  wire [4:0] P59;
  wire [3:0] P60;
  wire [2:0] P61;
  wire [1:0] P62;
  wire [0:0] P63;
  wire [63:0] R1;
  wire [53:0] R2;
  wire [64:0] aOut;
  U_SP_10_55 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, R1, R2);
  RC_54_54 S2 (R1[63:10], R2, aOut[64:10]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign Out = aOut[64:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
