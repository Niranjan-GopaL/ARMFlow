
module NR_1_42(
    input [0:0]IN1,
    input [41:0]IN2,
    output [41:0]Out
);
    assign Out = IN2;
endmodule
