//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 47
  second input length: 11
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_47_11(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56);
  input [46:0] IN1;
  input [10:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [10:0] P11;
  output [10:0] P12;
  output [10:0] P13;
  output [10:0] P14;
  output [10:0] P15;
  output [10:0] P16;
  output [10:0] P17;
  output [10:0] P18;
  output [10:0] P19;
  output [10:0] P20;
  output [10:0] P21;
  output [10:0] P22;
  output [10:0] P23;
  output [10:0] P24;
  output [10:0] P25;
  output [10:0] P26;
  output [10:0] P27;
  output [10:0] P28;
  output [10:0] P29;
  output [10:0] P30;
  output [10:0] P31;
  output [10:0] P32;
  output [10:0] P33;
  output [10:0] P34;
  output [10:0] P35;
  output [10:0] P36;
  output [10:0] P37;
  output [10:0] P38;
  output [10:0] P39;
  output [10:0] P40;
  output [10:0] P41;
  output [10:0] P42;
  output [10:0] P43;
  output [10:0] P44;
  output [10:0] P45;
  output [10:0] P46;
  output [9:0] P47;
  output [8:0] P48;
  output [7:0] P49;
  output [6:0] P50;
  output [5:0] P51;
  output [4:0] P52;
  output [3:0] P53;
  output [2:0] P54;
  output [1:0] P55;
  output [0:0] P56;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[0] = IN1[1]&IN2[10];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[1] = IN1[2]&IN2[9];
  assign P12[0] = IN1[2]&IN2[10];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[2] = IN1[3]&IN2[8];
  assign P12[1] = IN1[3]&IN2[9];
  assign P13[0] = IN1[3]&IN2[10];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[3] = IN1[4]&IN2[7];
  assign P12[2] = IN1[4]&IN2[8];
  assign P13[1] = IN1[4]&IN2[9];
  assign P14[0] = IN1[4]&IN2[10];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[4] = IN1[5]&IN2[6];
  assign P12[3] = IN1[5]&IN2[7];
  assign P13[2] = IN1[5]&IN2[8];
  assign P14[1] = IN1[5]&IN2[9];
  assign P15[0] = IN1[5]&IN2[10];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[5] = IN1[6]&IN2[5];
  assign P12[4] = IN1[6]&IN2[6];
  assign P13[3] = IN1[6]&IN2[7];
  assign P14[2] = IN1[6]&IN2[8];
  assign P15[1] = IN1[6]&IN2[9];
  assign P16[0] = IN1[6]&IN2[10];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[6] = IN1[7]&IN2[4];
  assign P12[5] = IN1[7]&IN2[5];
  assign P13[4] = IN1[7]&IN2[6];
  assign P14[3] = IN1[7]&IN2[7];
  assign P15[2] = IN1[7]&IN2[8];
  assign P16[1] = IN1[7]&IN2[9];
  assign P17[0] = IN1[7]&IN2[10];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[7] = IN1[8]&IN2[3];
  assign P12[6] = IN1[8]&IN2[4];
  assign P13[5] = IN1[8]&IN2[5];
  assign P14[4] = IN1[8]&IN2[6];
  assign P15[3] = IN1[8]&IN2[7];
  assign P16[2] = IN1[8]&IN2[8];
  assign P17[1] = IN1[8]&IN2[9];
  assign P18[0] = IN1[8]&IN2[10];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[8] = IN1[9]&IN2[2];
  assign P12[7] = IN1[9]&IN2[3];
  assign P13[6] = IN1[9]&IN2[4];
  assign P14[5] = IN1[9]&IN2[5];
  assign P15[4] = IN1[9]&IN2[6];
  assign P16[3] = IN1[9]&IN2[7];
  assign P17[2] = IN1[9]&IN2[8];
  assign P18[1] = IN1[9]&IN2[9];
  assign P19[0] = IN1[9]&IN2[10];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[9] = IN1[10]&IN2[1];
  assign P12[8] = IN1[10]&IN2[2];
  assign P13[7] = IN1[10]&IN2[3];
  assign P14[6] = IN1[10]&IN2[4];
  assign P15[5] = IN1[10]&IN2[5];
  assign P16[4] = IN1[10]&IN2[6];
  assign P17[3] = IN1[10]&IN2[7];
  assign P18[2] = IN1[10]&IN2[8];
  assign P19[1] = IN1[10]&IN2[9];
  assign P20[0] = IN1[10]&IN2[10];
  assign P11[10] = IN1[11]&IN2[0];
  assign P12[9] = IN1[11]&IN2[1];
  assign P13[8] = IN1[11]&IN2[2];
  assign P14[7] = IN1[11]&IN2[3];
  assign P15[6] = IN1[11]&IN2[4];
  assign P16[5] = IN1[11]&IN2[5];
  assign P17[4] = IN1[11]&IN2[6];
  assign P18[3] = IN1[11]&IN2[7];
  assign P19[2] = IN1[11]&IN2[8];
  assign P20[1] = IN1[11]&IN2[9];
  assign P21[0] = IN1[11]&IN2[10];
  assign P12[10] = IN1[12]&IN2[0];
  assign P13[9] = IN1[12]&IN2[1];
  assign P14[8] = IN1[12]&IN2[2];
  assign P15[7] = IN1[12]&IN2[3];
  assign P16[6] = IN1[12]&IN2[4];
  assign P17[5] = IN1[12]&IN2[5];
  assign P18[4] = IN1[12]&IN2[6];
  assign P19[3] = IN1[12]&IN2[7];
  assign P20[2] = IN1[12]&IN2[8];
  assign P21[1] = IN1[12]&IN2[9];
  assign P22[0] = IN1[12]&IN2[10];
  assign P13[10] = IN1[13]&IN2[0];
  assign P14[9] = IN1[13]&IN2[1];
  assign P15[8] = IN1[13]&IN2[2];
  assign P16[7] = IN1[13]&IN2[3];
  assign P17[6] = IN1[13]&IN2[4];
  assign P18[5] = IN1[13]&IN2[5];
  assign P19[4] = IN1[13]&IN2[6];
  assign P20[3] = IN1[13]&IN2[7];
  assign P21[2] = IN1[13]&IN2[8];
  assign P22[1] = IN1[13]&IN2[9];
  assign P23[0] = IN1[13]&IN2[10];
  assign P14[10] = IN1[14]&IN2[0];
  assign P15[9] = IN1[14]&IN2[1];
  assign P16[8] = IN1[14]&IN2[2];
  assign P17[7] = IN1[14]&IN2[3];
  assign P18[6] = IN1[14]&IN2[4];
  assign P19[5] = IN1[14]&IN2[5];
  assign P20[4] = IN1[14]&IN2[6];
  assign P21[3] = IN1[14]&IN2[7];
  assign P22[2] = IN1[14]&IN2[8];
  assign P23[1] = IN1[14]&IN2[9];
  assign P24[0] = IN1[14]&IN2[10];
  assign P15[10] = IN1[15]&IN2[0];
  assign P16[9] = IN1[15]&IN2[1];
  assign P17[8] = IN1[15]&IN2[2];
  assign P18[7] = IN1[15]&IN2[3];
  assign P19[6] = IN1[15]&IN2[4];
  assign P20[5] = IN1[15]&IN2[5];
  assign P21[4] = IN1[15]&IN2[6];
  assign P22[3] = IN1[15]&IN2[7];
  assign P23[2] = IN1[15]&IN2[8];
  assign P24[1] = IN1[15]&IN2[9];
  assign P25[0] = IN1[15]&IN2[10];
  assign P16[10] = IN1[16]&IN2[0];
  assign P17[9] = IN1[16]&IN2[1];
  assign P18[8] = IN1[16]&IN2[2];
  assign P19[7] = IN1[16]&IN2[3];
  assign P20[6] = IN1[16]&IN2[4];
  assign P21[5] = IN1[16]&IN2[5];
  assign P22[4] = IN1[16]&IN2[6];
  assign P23[3] = IN1[16]&IN2[7];
  assign P24[2] = IN1[16]&IN2[8];
  assign P25[1] = IN1[16]&IN2[9];
  assign P26[0] = IN1[16]&IN2[10];
  assign P17[10] = IN1[17]&IN2[0];
  assign P18[9] = IN1[17]&IN2[1];
  assign P19[8] = IN1[17]&IN2[2];
  assign P20[7] = IN1[17]&IN2[3];
  assign P21[6] = IN1[17]&IN2[4];
  assign P22[5] = IN1[17]&IN2[5];
  assign P23[4] = IN1[17]&IN2[6];
  assign P24[3] = IN1[17]&IN2[7];
  assign P25[2] = IN1[17]&IN2[8];
  assign P26[1] = IN1[17]&IN2[9];
  assign P27[0] = IN1[17]&IN2[10];
  assign P18[10] = IN1[18]&IN2[0];
  assign P19[9] = IN1[18]&IN2[1];
  assign P20[8] = IN1[18]&IN2[2];
  assign P21[7] = IN1[18]&IN2[3];
  assign P22[6] = IN1[18]&IN2[4];
  assign P23[5] = IN1[18]&IN2[5];
  assign P24[4] = IN1[18]&IN2[6];
  assign P25[3] = IN1[18]&IN2[7];
  assign P26[2] = IN1[18]&IN2[8];
  assign P27[1] = IN1[18]&IN2[9];
  assign P28[0] = IN1[18]&IN2[10];
  assign P19[10] = IN1[19]&IN2[0];
  assign P20[9] = IN1[19]&IN2[1];
  assign P21[8] = IN1[19]&IN2[2];
  assign P22[7] = IN1[19]&IN2[3];
  assign P23[6] = IN1[19]&IN2[4];
  assign P24[5] = IN1[19]&IN2[5];
  assign P25[4] = IN1[19]&IN2[6];
  assign P26[3] = IN1[19]&IN2[7];
  assign P27[2] = IN1[19]&IN2[8];
  assign P28[1] = IN1[19]&IN2[9];
  assign P29[0] = IN1[19]&IN2[10];
  assign P20[10] = IN1[20]&IN2[0];
  assign P21[9] = IN1[20]&IN2[1];
  assign P22[8] = IN1[20]&IN2[2];
  assign P23[7] = IN1[20]&IN2[3];
  assign P24[6] = IN1[20]&IN2[4];
  assign P25[5] = IN1[20]&IN2[5];
  assign P26[4] = IN1[20]&IN2[6];
  assign P27[3] = IN1[20]&IN2[7];
  assign P28[2] = IN1[20]&IN2[8];
  assign P29[1] = IN1[20]&IN2[9];
  assign P30[0] = IN1[20]&IN2[10];
  assign P21[10] = IN1[21]&IN2[0];
  assign P22[9] = IN1[21]&IN2[1];
  assign P23[8] = IN1[21]&IN2[2];
  assign P24[7] = IN1[21]&IN2[3];
  assign P25[6] = IN1[21]&IN2[4];
  assign P26[5] = IN1[21]&IN2[5];
  assign P27[4] = IN1[21]&IN2[6];
  assign P28[3] = IN1[21]&IN2[7];
  assign P29[2] = IN1[21]&IN2[8];
  assign P30[1] = IN1[21]&IN2[9];
  assign P31[0] = IN1[21]&IN2[10];
  assign P22[10] = IN1[22]&IN2[0];
  assign P23[9] = IN1[22]&IN2[1];
  assign P24[8] = IN1[22]&IN2[2];
  assign P25[7] = IN1[22]&IN2[3];
  assign P26[6] = IN1[22]&IN2[4];
  assign P27[5] = IN1[22]&IN2[5];
  assign P28[4] = IN1[22]&IN2[6];
  assign P29[3] = IN1[22]&IN2[7];
  assign P30[2] = IN1[22]&IN2[8];
  assign P31[1] = IN1[22]&IN2[9];
  assign P32[0] = IN1[22]&IN2[10];
  assign P23[10] = IN1[23]&IN2[0];
  assign P24[9] = IN1[23]&IN2[1];
  assign P25[8] = IN1[23]&IN2[2];
  assign P26[7] = IN1[23]&IN2[3];
  assign P27[6] = IN1[23]&IN2[4];
  assign P28[5] = IN1[23]&IN2[5];
  assign P29[4] = IN1[23]&IN2[6];
  assign P30[3] = IN1[23]&IN2[7];
  assign P31[2] = IN1[23]&IN2[8];
  assign P32[1] = IN1[23]&IN2[9];
  assign P33[0] = IN1[23]&IN2[10];
  assign P24[10] = IN1[24]&IN2[0];
  assign P25[9] = IN1[24]&IN2[1];
  assign P26[8] = IN1[24]&IN2[2];
  assign P27[7] = IN1[24]&IN2[3];
  assign P28[6] = IN1[24]&IN2[4];
  assign P29[5] = IN1[24]&IN2[5];
  assign P30[4] = IN1[24]&IN2[6];
  assign P31[3] = IN1[24]&IN2[7];
  assign P32[2] = IN1[24]&IN2[8];
  assign P33[1] = IN1[24]&IN2[9];
  assign P34[0] = IN1[24]&IN2[10];
  assign P25[10] = IN1[25]&IN2[0];
  assign P26[9] = IN1[25]&IN2[1];
  assign P27[8] = IN1[25]&IN2[2];
  assign P28[7] = IN1[25]&IN2[3];
  assign P29[6] = IN1[25]&IN2[4];
  assign P30[5] = IN1[25]&IN2[5];
  assign P31[4] = IN1[25]&IN2[6];
  assign P32[3] = IN1[25]&IN2[7];
  assign P33[2] = IN1[25]&IN2[8];
  assign P34[1] = IN1[25]&IN2[9];
  assign P35[0] = IN1[25]&IN2[10];
  assign P26[10] = IN1[26]&IN2[0];
  assign P27[9] = IN1[26]&IN2[1];
  assign P28[8] = IN1[26]&IN2[2];
  assign P29[7] = IN1[26]&IN2[3];
  assign P30[6] = IN1[26]&IN2[4];
  assign P31[5] = IN1[26]&IN2[5];
  assign P32[4] = IN1[26]&IN2[6];
  assign P33[3] = IN1[26]&IN2[7];
  assign P34[2] = IN1[26]&IN2[8];
  assign P35[1] = IN1[26]&IN2[9];
  assign P36[0] = IN1[26]&IN2[10];
  assign P27[10] = IN1[27]&IN2[0];
  assign P28[9] = IN1[27]&IN2[1];
  assign P29[8] = IN1[27]&IN2[2];
  assign P30[7] = IN1[27]&IN2[3];
  assign P31[6] = IN1[27]&IN2[4];
  assign P32[5] = IN1[27]&IN2[5];
  assign P33[4] = IN1[27]&IN2[6];
  assign P34[3] = IN1[27]&IN2[7];
  assign P35[2] = IN1[27]&IN2[8];
  assign P36[1] = IN1[27]&IN2[9];
  assign P37[0] = IN1[27]&IN2[10];
  assign P28[10] = IN1[28]&IN2[0];
  assign P29[9] = IN1[28]&IN2[1];
  assign P30[8] = IN1[28]&IN2[2];
  assign P31[7] = IN1[28]&IN2[3];
  assign P32[6] = IN1[28]&IN2[4];
  assign P33[5] = IN1[28]&IN2[5];
  assign P34[4] = IN1[28]&IN2[6];
  assign P35[3] = IN1[28]&IN2[7];
  assign P36[2] = IN1[28]&IN2[8];
  assign P37[1] = IN1[28]&IN2[9];
  assign P38[0] = IN1[28]&IN2[10];
  assign P29[10] = IN1[29]&IN2[0];
  assign P30[9] = IN1[29]&IN2[1];
  assign P31[8] = IN1[29]&IN2[2];
  assign P32[7] = IN1[29]&IN2[3];
  assign P33[6] = IN1[29]&IN2[4];
  assign P34[5] = IN1[29]&IN2[5];
  assign P35[4] = IN1[29]&IN2[6];
  assign P36[3] = IN1[29]&IN2[7];
  assign P37[2] = IN1[29]&IN2[8];
  assign P38[1] = IN1[29]&IN2[9];
  assign P39[0] = IN1[29]&IN2[10];
  assign P30[10] = IN1[30]&IN2[0];
  assign P31[9] = IN1[30]&IN2[1];
  assign P32[8] = IN1[30]&IN2[2];
  assign P33[7] = IN1[30]&IN2[3];
  assign P34[6] = IN1[30]&IN2[4];
  assign P35[5] = IN1[30]&IN2[5];
  assign P36[4] = IN1[30]&IN2[6];
  assign P37[3] = IN1[30]&IN2[7];
  assign P38[2] = IN1[30]&IN2[8];
  assign P39[1] = IN1[30]&IN2[9];
  assign P40[0] = IN1[30]&IN2[10];
  assign P31[10] = IN1[31]&IN2[0];
  assign P32[9] = IN1[31]&IN2[1];
  assign P33[8] = IN1[31]&IN2[2];
  assign P34[7] = IN1[31]&IN2[3];
  assign P35[6] = IN1[31]&IN2[4];
  assign P36[5] = IN1[31]&IN2[5];
  assign P37[4] = IN1[31]&IN2[6];
  assign P38[3] = IN1[31]&IN2[7];
  assign P39[2] = IN1[31]&IN2[8];
  assign P40[1] = IN1[31]&IN2[9];
  assign P41[0] = IN1[31]&IN2[10];
  assign P32[10] = IN1[32]&IN2[0];
  assign P33[9] = IN1[32]&IN2[1];
  assign P34[8] = IN1[32]&IN2[2];
  assign P35[7] = IN1[32]&IN2[3];
  assign P36[6] = IN1[32]&IN2[4];
  assign P37[5] = IN1[32]&IN2[5];
  assign P38[4] = IN1[32]&IN2[6];
  assign P39[3] = IN1[32]&IN2[7];
  assign P40[2] = IN1[32]&IN2[8];
  assign P41[1] = IN1[32]&IN2[9];
  assign P42[0] = IN1[32]&IN2[10];
  assign P33[10] = IN1[33]&IN2[0];
  assign P34[9] = IN1[33]&IN2[1];
  assign P35[8] = IN1[33]&IN2[2];
  assign P36[7] = IN1[33]&IN2[3];
  assign P37[6] = IN1[33]&IN2[4];
  assign P38[5] = IN1[33]&IN2[5];
  assign P39[4] = IN1[33]&IN2[6];
  assign P40[3] = IN1[33]&IN2[7];
  assign P41[2] = IN1[33]&IN2[8];
  assign P42[1] = IN1[33]&IN2[9];
  assign P43[0] = IN1[33]&IN2[10];
  assign P34[10] = IN1[34]&IN2[0];
  assign P35[9] = IN1[34]&IN2[1];
  assign P36[8] = IN1[34]&IN2[2];
  assign P37[7] = IN1[34]&IN2[3];
  assign P38[6] = IN1[34]&IN2[4];
  assign P39[5] = IN1[34]&IN2[5];
  assign P40[4] = IN1[34]&IN2[6];
  assign P41[3] = IN1[34]&IN2[7];
  assign P42[2] = IN1[34]&IN2[8];
  assign P43[1] = IN1[34]&IN2[9];
  assign P44[0] = IN1[34]&IN2[10];
  assign P35[10] = IN1[35]&IN2[0];
  assign P36[9] = IN1[35]&IN2[1];
  assign P37[8] = IN1[35]&IN2[2];
  assign P38[7] = IN1[35]&IN2[3];
  assign P39[6] = IN1[35]&IN2[4];
  assign P40[5] = IN1[35]&IN2[5];
  assign P41[4] = IN1[35]&IN2[6];
  assign P42[3] = IN1[35]&IN2[7];
  assign P43[2] = IN1[35]&IN2[8];
  assign P44[1] = IN1[35]&IN2[9];
  assign P45[0] = IN1[35]&IN2[10];
  assign P36[10] = IN1[36]&IN2[0];
  assign P37[9] = IN1[36]&IN2[1];
  assign P38[8] = IN1[36]&IN2[2];
  assign P39[7] = IN1[36]&IN2[3];
  assign P40[6] = IN1[36]&IN2[4];
  assign P41[5] = IN1[36]&IN2[5];
  assign P42[4] = IN1[36]&IN2[6];
  assign P43[3] = IN1[36]&IN2[7];
  assign P44[2] = IN1[36]&IN2[8];
  assign P45[1] = IN1[36]&IN2[9];
  assign P46[0] = IN1[36]&IN2[10];
  assign P37[10] = IN1[37]&IN2[0];
  assign P38[9] = IN1[37]&IN2[1];
  assign P39[8] = IN1[37]&IN2[2];
  assign P40[7] = IN1[37]&IN2[3];
  assign P41[6] = IN1[37]&IN2[4];
  assign P42[5] = IN1[37]&IN2[5];
  assign P43[4] = IN1[37]&IN2[6];
  assign P44[3] = IN1[37]&IN2[7];
  assign P45[2] = IN1[37]&IN2[8];
  assign P46[1] = IN1[37]&IN2[9];
  assign P47[0] = IN1[37]&IN2[10];
  assign P38[10] = IN1[38]&IN2[0];
  assign P39[9] = IN1[38]&IN2[1];
  assign P40[8] = IN1[38]&IN2[2];
  assign P41[7] = IN1[38]&IN2[3];
  assign P42[6] = IN1[38]&IN2[4];
  assign P43[5] = IN1[38]&IN2[5];
  assign P44[4] = IN1[38]&IN2[6];
  assign P45[3] = IN1[38]&IN2[7];
  assign P46[2] = IN1[38]&IN2[8];
  assign P47[1] = IN1[38]&IN2[9];
  assign P48[0] = IN1[38]&IN2[10];
  assign P39[10] = IN1[39]&IN2[0];
  assign P40[9] = IN1[39]&IN2[1];
  assign P41[8] = IN1[39]&IN2[2];
  assign P42[7] = IN1[39]&IN2[3];
  assign P43[6] = IN1[39]&IN2[4];
  assign P44[5] = IN1[39]&IN2[5];
  assign P45[4] = IN1[39]&IN2[6];
  assign P46[3] = IN1[39]&IN2[7];
  assign P47[2] = IN1[39]&IN2[8];
  assign P48[1] = IN1[39]&IN2[9];
  assign P49[0] = IN1[39]&IN2[10];
  assign P40[10] = IN1[40]&IN2[0];
  assign P41[9] = IN1[40]&IN2[1];
  assign P42[8] = IN1[40]&IN2[2];
  assign P43[7] = IN1[40]&IN2[3];
  assign P44[6] = IN1[40]&IN2[4];
  assign P45[5] = IN1[40]&IN2[5];
  assign P46[4] = IN1[40]&IN2[6];
  assign P47[3] = IN1[40]&IN2[7];
  assign P48[2] = IN1[40]&IN2[8];
  assign P49[1] = IN1[40]&IN2[9];
  assign P50[0] = IN1[40]&IN2[10];
  assign P41[10] = IN1[41]&IN2[0];
  assign P42[9] = IN1[41]&IN2[1];
  assign P43[8] = IN1[41]&IN2[2];
  assign P44[7] = IN1[41]&IN2[3];
  assign P45[6] = IN1[41]&IN2[4];
  assign P46[5] = IN1[41]&IN2[5];
  assign P47[4] = IN1[41]&IN2[6];
  assign P48[3] = IN1[41]&IN2[7];
  assign P49[2] = IN1[41]&IN2[8];
  assign P50[1] = IN1[41]&IN2[9];
  assign P51[0] = IN1[41]&IN2[10];
  assign P42[10] = IN1[42]&IN2[0];
  assign P43[9] = IN1[42]&IN2[1];
  assign P44[8] = IN1[42]&IN2[2];
  assign P45[7] = IN1[42]&IN2[3];
  assign P46[6] = IN1[42]&IN2[4];
  assign P47[5] = IN1[42]&IN2[5];
  assign P48[4] = IN1[42]&IN2[6];
  assign P49[3] = IN1[42]&IN2[7];
  assign P50[2] = IN1[42]&IN2[8];
  assign P51[1] = IN1[42]&IN2[9];
  assign P52[0] = IN1[42]&IN2[10];
  assign P43[10] = IN1[43]&IN2[0];
  assign P44[9] = IN1[43]&IN2[1];
  assign P45[8] = IN1[43]&IN2[2];
  assign P46[7] = IN1[43]&IN2[3];
  assign P47[6] = IN1[43]&IN2[4];
  assign P48[5] = IN1[43]&IN2[5];
  assign P49[4] = IN1[43]&IN2[6];
  assign P50[3] = IN1[43]&IN2[7];
  assign P51[2] = IN1[43]&IN2[8];
  assign P52[1] = IN1[43]&IN2[9];
  assign P53[0] = IN1[43]&IN2[10];
  assign P44[10] = IN1[44]&IN2[0];
  assign P45[9] = IN1[44]&IN2[1];
  assign P46[8] = IN1[44]&IN2[2];
  assign P47[7] = IN1[44]&IN2[3];
  assign P48[6] = IN1[44]&IN2[4];
  assign P49[5] = IN1[44]&IN2[5];
  assign P50[4] = IN1[44]&IN2[6];
  assign P51[3] = IN1[44]&IN2[7];
  assign P52[2] = IN1[44]&IN2[8];
  assign P53[1] = IN1[44]&IN2[9];
  assign P54[0] = IN1[44]&IN2[10];
  assign P45[10] = IN1[45]&IN2[0];
  assign P46[9] = IN1[45]&IN2[1];
  assign P47[8] = IN1[45]&IN2[2];
  assign P48[7] = IN1[45]&IN2[3];
  assign P49[6] = IN1[45]&IN2[4];
  assign P50[5] = IN1[45]&IN2[5];
  assign P51[4] = IN1[45]&IN2[6];
  assign P52[3] = IN1[45]&IN2[7];
  assign P53[2] = IN1[45]&IN2[8];
  assign P54[1] = IN1[45]&IN2[9];
  assign P55[0] = IN1[45]&IN2[10];
  assign P46[10] = IN1[46]&IN2[0];
  assign P47[9] = IN1[46]&IN2[1];
  assign P48[8] = IN1[46]&IN2[2];
  assign P49[7] = IN1[46]&IN2[3];
  assign P50[6] = IN1[46]&IN2[4];
  assign P51[5] = IN1[46]&IN2[5];
  assign P52[4] = IN1[46]&IN2[6];
  assign P53[3] = IN1[46]&IN2[7];
  assign P54[2] = IN1[46]&IN2[8];
  assign P55[1] = IN1[46]&IN2[9];
  assign P56[0] = IN1[46]&IN2[10];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [10:0] IN11;
  input [10:0] IN12;
  input [10:0] IN13;
  input [10:0] IN14;
  input [10:0] IN15;
  input [10:0] IN16;
  input [10:0] IN17;
  input [10:0] IN18;
  input [10:0] IN19;
  input [10:0] IN20;
  input [10:0] IN21;
  input [10:0] IN22;
  input [10:0] IN23;
  input [10:0] IN24;
  input [10:0] IN25;
  input [10:0] IN26;
  input [10:0] IN27;
  input [10:0] IN28;
  input [10:0] IN29;
  input [10:0] IN30;
  input [10:0] IN31;
  input [10:0] IN32;
  input [10:0] IN33;
  input [10:0] IN34;
  input [10:0] IN35;
  input [10:0] IN36;
  input [10:0] IN37;
  input [10:0] IN38;
  input [10:0] IN39;
  input [10:0] IN40;
  input [10:0] IN41;
  input [10:0] IN42;
  input [10:0] IN43;
  input [10:0] IN44;
  input [10:0] IN45;
  input [10:0] IN46;
  input [9:0] IN47;
  input [8:0] IN48;
  input [7:0] IN49;
  input [6:0] IN50;
  input [5:0] IN51;
  input [4:0] IN52;
  input [3:0] IN53;
  input [2:0] IN54;
  input [1:0] IN55;
  input [0:0] IN56;
  output [56:0] Out1;
  output [9:0] Out2;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1346;
  wire w1348;
  wire w1350;
  wire w1352;
  wire w1354;
  wire w1356;
  wire w1358;
  wire w1360;
  wire w1362;
  wire w1364;
  wire w1366;
  wire w1368;
  wire w1370;
  wire w1372;
  wire w1374;
  wire w1376;
  wire w1378;
  wire w1380;
  wire w1382;
  wire w1384;
  wire w1386;
  wire w1388;
  wire w1390;
  wire w1392;
  wire w1394;
  wire w1396;
  wire w1398;
  wire w1400;
  wire w1402;
  wire w1404;
  wire w1406;
  wire w1408;
  wire w1410;
  wire w1412;
  wire w1414;
  wire w1416;
  wire w1418;
  wire w1420;
  wire w1422;
  wire w1424;
  wire w1426;
  wire w1428;
  wire w1430;
  wire w1432;
  wire w1434;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w518);
  FullAdder U1 (w518, IN2[0], IN2[1], w519, w520);
  FullAdder U2 (w520, IN3[0], IN3[1], w521, w522);
  FullAdder U3 (w522, IN4[0], IN4[1], w523, w524);
  FullAdder U4 (w524, IN5[0], IN5[1], w525, w526);
  FullAdder U5 (w526, IN6[0], IN6[1], w527, w528);
  FullAdder U6 (w528, IN7[0], IN7[1], w529, w530);
  FullAdder U7 (w530, IN8[0], IN8[1], w531, w532);
  FullAdder U8 (w532, IN9[0], IN9[1], w533, w534);
  FullAdder U9 (w534, IN10[0], IN10[1], w535, w536);
  FullAdder U10 (w536, IN11[0], IN11[1], w537, w538);
  FullAdder U11 (w538, IN12[0], IN12[1], w539, w540);
  FullAdder U12 (w540, IN13[0], IN13[1], w541, w542);
  FullAdder U13 (w542, IN14[0], IN14[1], w543, w544);
  FullAdder U14 (w544, IN15[0], IN15[1], w545, w546);
  FullAdder U15 (w546, IN16[0], IN16[1], w547, w548);
  FullAdder U16 (w548, IN17[0], IN17[1], w549, w550);
  FullAdder U17 (w550, IN18[0], IN18[1], w551, w552);
  FullAdder U18 (w552, IN19[0], IN19[1], w553, w554);
  FullAdder U19 (w554, IN20[0], IN20[1], w555, w556);
  FullAdder U20 (w556, IN21[0], IN21[1], w557, w558);
  FullAdder U21 (w558, IN22[0], IN22[1], w559, w560);
  FullAdder U22 (w560, IN23[0], IN23[1], w561, w562);
  FullAdder U23 (w562, IN24[0], IN24[1], w563, w564);
  FullAdder U24 (w564, IN25[0], IN25[1], w565, w566);
  FullAdder U25 (w566, IN26[0], IN26[1], w567, w568);
  FullAdder U26 (w568, IN27[0], IN27[1], w569, w570);
  FullAdder U27 (w570, IN28[0], IN28[1], w571, w572);
  FullAdder U28 (w572, IN29[0], IN29[1], w573, w574);
  FullAdder U29 (w574, IN30[0], IN30[1], w575, w576);
  FullAdder U30 (w576, IN31[0], IN31[1], w577, w578);
  FullAdder U31 (w578, IN32[0], IN32[1], w579, w580);
  FullAdder U32 (w580, IN33[0], IN33[1], w581, w582);
  FullAdder U33 (w582, IN34[0], IN34[1], w583, w584);
  FullAdder U34 (w584, IN35[0], IN35[1], w585, w586);
  FullAdder U35 (w586, IN36[0], IN36[1], w587, w588);
  FullAdder U36 (w588, IN37[0], IN37[1], w589, w590);
  FullAdder U37 (w590, IN38[0], IN38[1], w591, w592);
  FullAdder U38 (w592, IN39[0], IN39[1], w593, w594);
  FullAdder U39 (w594, IN40[0], IN40[1], w595, w596);
  FullAdder U40 (w596, IN41[0], IN41[1], w597, w598);
  FullAdder U41 (w598, IN42[0], IN42[1], w599, w600);
  FullAdder U42 (w600, IN43[0], IN43[1], w601, w602);
  FullAdder U43 (w602, IN44[0], IN44[1], w603, w604);
  FullAdder U44 (w604, IN45[0], IN45[1], w605, w606);
  FullAdder U45 (w606, IN46[0], IN46[1], w607, w608);
  HalfAdder U46 (w519, IN2[2], Out1[2], w610);
  FullAdder U47 (w610, w521, IN3[2], w611, w612);
  FullAdder U48 (w612, w523, IN4[2], w613, w614);
  FullAdder U49 (w614, w525, IN5[2], w615, w616);
  FullAdder U50 (w616, w527, IN6[2], w617, w618);
  FullAdder U51 (w618, w529, IN7[2], w619, w620);
  FullAdder U52 (w620, w531, IN8[2], w621, w622);
  FullAdder U53 (w622, w533, IN9[2], w623, w624);
  FullAdder U54 (w624, w535, IN10[2], w625, w626);
  FullAdder U55 (w626, w537, IN11[2], w627, w628);
  FullAdder U56 (w628, w539, IN12[2], w629, w630);
  FullAdder U57 (w630, w541, IN13[2], w631, w632);
  FullAdder U58 (w632, w543, IN14[2], w633, w634);
  FullAdder U59 (w634, w545, IN15[2], w635, w636);
  FullAdder U60 (w636, w547, IN16[2], w637, w638);
  FullAdder U61 (w638, w549, IN17[2], w639, w640);
  FullAdder U62 (w640, w551, IN18[2], w641, w642);
  FullAdder U63 (w642, w553, IN19[2], w643, w644);
  FullAdder U64 (w644, w555, IN20[2], w645, w646);
  FullAdder U65 (w646, w557, IN21[2], w647, w648);
  FullAdder U66 (w648, w559, IN22[2], w649, w650);
  FullAdder U67 (w650, w561, IN23[2], w651, w652);
  FullAdder U68 (w652, w563, IN24[2], w653, w654);
  FullAdder U69 (w654, w565, IN25[2], w655, w656);
  FullAdder U70 (w656, w567, IN26[2], w657, w658);
  FullAdder U71 (w658, w569, IN27[2], w659, w660);
  FullAdder U72 (w660, w571, IN28[2], w661, w662);
  FullAdder U73 (w662, w573, IN29[2], w663, w664);
  FullAdder U74 (w664, w575, IN30[2], w665, w666);
  FullAdder U75 (w666, w577, IN31[2], w667, w668);
  FullAdder U76 (w668, w579, IN32[2], w669, w670);
  FullAdder U77 (w670, w581, IN33[2], w671, w672);
  FullAdder U78 (w672, w583, IN34[2], w673, w674);
  FullAdder U79 (w674, w585, IN35[2], w675, w676);
  FullAdder U80 (w676, w587, IN36[2], w677, w678);
  FullAdder U81 (w678, w589, IN37[2], w679, w680);
  FullAdder U82 (w680, w591, IN38[2], w681, w682);
  FullAdder U83 (w682, w593, IN39[2], w683, w684);
  FullAdder U84 (w684, w595, IN40[2], w685, w686);
  FullAdder U85 (w686, w597, IN41[2], w687, w688);
  FullAdder U86 (w688, w599, IN42[2], w689, w690);
  FullAdder U87 (w690, w601, IN43[2], w691, w692);
  FullAdder U88 (w692, w603, IN44[2], w693, w694);
  FullAdder U89 (w694, w605, IN45[2], w695, w696);
  FullAdder U90 (w696, w607, IN46[2], w697, w698);
  FullAdder U91 (w698, w608, IN47[0], w699, w700);
  HalfAdder U92 (w611, IN3[3], Out1[3], w702);
  FullAdder U93 (w702, w613, IN4[3], w703, w704);
  FullAdder U94 (w704, w615, IN5[3], w705, w706);
  FullAdder U95 (w706, w617, IN6[3], w707, w708);
  FullAdder U96 (w708, w619, IN7[3], w709, w710);
  FullAdder U97 (w710, w621, IN8[3], w711, w712);
  FullAdder U98 (w712, w623, IN9[3], w713, w714);
  FullAdder U99 (w714, w625, IN10[3], w715, w716);
  FullAdder U100 (w716, w627, IN11[3], w717, w718);
  FullAdder U101 (w718, w629, IN12[3], w719, w720);
  FullAdder U102 (w720, w631, IN13[3], w721, w722);
  FullAdder U103 (w722, w633, IN14[3], w723, w724);
  FullAdder U104 (w724, w635, IN15[3], w725, w726);
  FullAdder U105 (w726, w637, IN16[3], w727, w728);
  FullAdder U106 (w728, w639, IN17[3], w729, w730);
  FullAdder U107 (w730, w641, IN18[3], w731, w732);
  FullAdder U108 (w732, w643, IN19[3], w733, w734);
  FullAdder U109 (w734, w645, IN20[3], w735, w736);
  FullAdder U110 (w736, w647, IN21[3], w737, w738);
  FullAdder U111 (w738, w649, IN22[3], w739, w740);
  FullAdder U112 (w740, w651, IN23[3], w741, w742);
  FullAdder U113 (w742, w653, IN24[3], w743, w744);
  FullAdder U114 (w744, w655, IN25[3], w745, w746);
  FullAdder U115 (w746, w657, IN26[3], w747, w748);
  FullAdder U116 (w748, w659, IN27[3], w749, w750);
  FullAdder U117 (w750, w661, IN28[3], w751, w752);
  FullAdder U118 (w752, w663, IN29[3], w753, w754);
  FullAdder U119 (w754, w665, IN30[3], w755, w756);
  FullAdder U120 (w756, w667, IN31[3], w757, w758);
  FullAdder U121 (w758, w669, IN32[3], w759, w760);
  FullAdder U122 (w760, w671, IN33[3], w761, w762);
  FullAdder U123 (w762, w673, IN34[3], w763, w764);
  FullAdder U124 (w764, w675, IN35[3], w765, w766);
  FullAdder U125 (w766, w677, IN36[3], w767, w768);
  FullAdder U126 (w768, w679, IN37[3], w769, w770);
  FullAdder U127 (w770, w681, IN38[3], w771, w772);
  FullAdder U128 (w772, w683, IN39[3], w773, w774);
  FullAdder U129 (w774, w685, IN40[3], w775, w776);
  FullAdder U130 (w776, w687, IN41[3], w777, w778);
  FullAdder U131 (w778, w689, IN42[3], w779, w780);
  FullAdder U132 (w780, w691, IN43[3], w781, w782);
  FullAdder U133 (w782, w693, IN44[3], w783, w784);
  FullAdder U134 (w784, w695, IN45[3], w785, w786);
  FullAdder U135 (w786, w697, IN46[3], w787, w788);
  FullAdder U136 (w788, w699, IN47[1], w789, w790);
  FullAdder U137 (w790, w700, IN48[0], w791, w792);
  HalfAdder U138 (w703, IN4[4], Out1[4], w794);
  FullAdder U139 (w794, w705, IN5[4], w795, w796);
  FullAdder U140 (w796, w707, IN6[4], w797, w798);
  FullAdder U141 (w798, w709, IN7[4], w799, w800);
  FullAdder U142 (w800, w711, IN8[4], w801, w802);
  FullAdder U143 (w802, w713, IN9[4], w803, w804);
  FullAdder U144 (w804, w715, IN10[4], w805, w806);
  FullAdder U145 (w806, w717, IN11[4], w807, w808);
  FullAdder U146 (w808, w719, IN12[4], w809, w810);
  FullAdder U147 (w810, w721, IN13[4], w811, w812);
  FullAdder U148 (w812, w723, IN14[4], w813, w814);
  FullAdder U149 (w814, w725, IN15[4], w815, w816);
  FullAdder U150 (w816, w727, IN16[4], w817, w818);
  FullAdder U151 (w818, w729, IN17[4], w819, w820);
  FullAdder U152 (w820, w731, IN18[4], w821, w822);
  FullAdder U153 (w822, w733, IN19[4], w823, w824);
  FullAdder U154 (w824, w735, IN20[4], w825, w826);
  FullAdder U155 (w826, w737, IN21[4], w827, w828);
  FullAdder U156 (w828, w739, IN22[4], w829, w830);
  FullAdder U157 (w830, w741, IN23[4], w831, w832);
  FullAdder U158 (w832, w743, IN24[4], w833, w834);
  FullAdder U159 (w834, w745, IN25[4], w835, w836);
  FullAdder U160 (w836, w747, IN26[4], w837, w838);
  FullAdder U161 (w838, w749, IN27[4], w839, w840);
  FullAdder U162 (w840, w751, IN28[4], w841, w842);
  FullAdder U163 (w842, w753, IN29[4], w843, w844);
  FullAdder U164 (w844, w755, IN30[4], w845, w846);
  FullAdder U165 (w846, w757, IN31[4], w847, w848);
  FullAdder U166 (w848, w759, IN32[4], w849, w850);
  FullAdder U167 (w850, w761, IN33[4], w851, w852);
  FullAdder U168 (w852, w763, IN34[4], w853, w854);
  FullAdder U169 (w854, w765, IN35[4], w855, w856);
  FullAdder U170 (w856, w767, IN36[4], w857, w858);
  FullAdder U171 (w858, w769, IN37[4], w859, w860);
  FullAdder U172 (w860, w771, IN38[4], w861, w862);
  FullAdder U173 (w862, w773, IN39[4], w863, w864);
  FullAdder U174 (w864, w775, IN40[4], w865, w866);
  FullAdder U175 (w866, w777, IN41[4], w867, w868);
  FullAdder U176 (w868, w779, IN42[4], w869, w870);
  FullAdder U177 (w870, w781, IN43[4], w871, w872);
  FullAdder U178 (w872, w783, IN44[4], w873, w874);
  FullAdder U179 (w874, w785, IN45[4], w875, w876);
  FullAdder U180 (w876, w787, IN46[4], w877, w878);
  FullAdder U181 (w878, w789, IN47[2], w879, w880);
  FullAdder U182 (w880, w791, IN48[1], w881, w882);
  FullAdder U183 (w882, w792, IN49[0], w883, w884);
  HalfAdder U184 (w795, IN5[5], Out1[5], w886);
  FullAdder U185 (w886, w797, IN6[5], w887, w888);
  FullAdder U186 (w888, w799, IN7[5], w889, w890);
  FullAdder U187 (w890, w801, IN8[5], w891, w892);
  FullAdder U188 (w892, w803, IN9[5], w893, w894);
  FullAdder U189 (w894, w805, IN10[5], w895, w896);
  FullAdder U190 (w896, w807, IN11[5], w897, w898);
  FullAdder U191 (w898, w809, IN12[5], w899, w900);
  FullAdder U192 (w900, w811, IN13[5], w901, w902);
  FullAdder U193 (w902, w813, IN14[5], w903, w904);
  FullAdder U194 (w904, w815, IN15[5], w905, w906);
  FullAdder U195 (w906, w817, IN16[5], w907, w908);
  FullAdder U196 (w908, w819, IN17[5], w909, w910);
  FullAdder U197 (w910, w821, IN18[5], w911, w912);
  FullAdder U198 (w912, w823, IN19[5], w913, w914);
  FullAdder U199 (w914, w825, IN20[5], w915, w916);
  FullAdder U200 (w916, w827, IN21[5], w917, w918);
  FullAdder U201 (w918, w829, IN22[5], w919, w920);
  FullAdder U202 (w920, w831, IN23[5], w921, w922);
  FullAdder U203 (w922, w833, IN24[5], w923, w924);
  FullAdder U204 (w924, w835, IN25[5], w925, w926);
  FullAdder U205 (w926, w837, IN26[5], w927, w928);
  FullAdder U206 (w928, w839, IN27[5], w929, w930);
  FullAdder U207 (w930, w841, IN28[5], w931, w932);
  FullAdder U208 (w932, w843, IN29[5], w933, w934);
  FullAdder U209 (w934, w845, IN30[5], w935, w936);
  FullAdder U210 (w936, w847, IN31[5], w937, w938);
  FullAdder U211 (w938, w849, IN32[5], w939, w940);
  FullAdder U212 (w940, w851, IN33[5], w941, w942);
  FullAdder U213 (w942, w853, IN34[5], w943, w944);
  FullAdder U214 (w944, w855, IN35[5], w945, w946);
  FullAdder U215 (w946, w857, IN36[5], w947, w948);
  FullAdder U216 (w948, w859, IN37[5], w949, w950);
  FullAdder U217 (w950, w861, IN38[5], w951, w952);
  FullAdder U218 (w952, w863, IN39[5], w953, w954);
  FullAdder U219 (w954, w865, IN40[5], w955, w956);
  FullAdder U220 (w956, w867, IN41[5], w957, w958);
  FullAdder U221 (w958, w869, IN42[5], w959, w960);
  FullAdder U222 (w960, w871, IN43[5], w961, w962);
  FullAdder U223 (w962, w873, IN44[5], w963, w964);
  FullAdder U224 (w964, w875, IN45[5], w965, w966);
  FullAdder U225 (w966, w877, IN46[5], w967, w968);
  FullAdder U226 (w968, w879, IN47[3], w969, w970);
  FullAdder U227 (w970, w881, IN48[2], w971, w972);
  FullAdder U228 (w972, w883, IN49[1], w973, w974);
  FullAdder U229 (w974, w884, IN50[0], w975, w976);
  HalfAdder U230 (w887, IN6[6], Out1[6], w978);
  FullAdder U231 (w978, w889, IN7[6], w979, w980);
  FullAdder U232 (w980, w891, IN8[6], w981, w982);
  FullAdder U233 (w982, w893, IN9[6], w983, w984);
  FullAdder U234 (w984, w895, IN10[6], w985, w986);
  FullAdder U235 (w986, w897, IN11[6], w987, w988);
  FullAdder U236 (w988, w899, IN12[6], w989, w990);
  FullAdder U237 (w990, w901, IN13[6], w991, w992);
  FullAdder U238 (w992, w903, IN14[6], w993, w994);
  FullAdder U239 (w994, w905, IN15[6], w995, w996);
  FullAdder U240 (w996, w907, IN16[6], w997, w998);
  FullAdder U241 (w998, w909, IN17[6], w999, w1000);
  FullAdder U242 (w1000, w911, IN18[6], w1001, w1002);
  FullAdder U243 (w1002, w913, IN19[6], w1003, w1004);
  FullAdder U244 (w1004, w915, IN20[6], w1005, w1006);
  FullAdder U245 (w1006, w917, IN21[6], w1007, w1008);
  FullAdder U246 (w1008, w919, IN22[6], w1009, w1010);
  FullAdder U247 (w1010, w921, IN23[6], w1011, w1012);
  FullAdder U248 (w1012, w923, IN24[6], w1013, w1014);
  FullAdder U249 (w1014, w925, IN25[6], w1015, w1016);
  FullAdder U250 (w1016, w927, IN26[6], w1017, w1018);
  FullAdder U251 (w1018, w929, IN27[6], w1019, w1020);
  FullAdder U252 (w1020, w931, IN28[6], w1021, w1022);
  FullAdder U253 (w1022, w933, IN29[6], w1023, w1024);
  FullAdder U254 (w1024, w935, IN30[6], w1025, w1026);
  FullAdder U255 (w1026, w937, IN31[6], w1027, w1028);
  FullAdder U256 (w1028, w939, IN32[6], w1029, w1030);
  FullAdder U257 (w1030, w941, IN33[6], w1031, w1032);
  FullAdder U258 (w1032, w943, IN34[6], w1033, w1034);
  FullAdder U259 (w1034, w945, IN35[6], w1035, w1036);
  FullAdder U260 (w1036, w947, IN36[6], w1037, w1038);
  FullAdder U261 (w1038, w949, IN37[6], w1039, w1040);
  FullAdder U262 (w1040, w951, IN38[6], w1041, w1042);
  FullAdder U263 (w1042, w953, IN39[6], w1043, w1044);
  FullAdder U264 (w1044, w955, IN40[6], w1045, w1046);
  FullAdder U265 (w1046, w957, IN41[6], w1047, w1048);
  FullAdder U266 (w1048, w959, IN42[6], w1049, w1050);
  FullAdder U267 (w1050, w961, IN43[6], w1051, w1052);
  FullAdder U268 (w1052, w963, IN44[6], w1053, w1054);
  FullAdder U269 (w1054, w965, IN45[6], w1055, w1056);
  FullAdder U270 (w1056, w967, IN46[6], w1057, w1058);
  FullAdder U271 (w1058, w969, IN47[4], w1059, w1060);
  FullAdder U272 (w1060, w971, IN48[3], w1061, w1062);
  FullAdder U273 (w1062, w973, IN49[2], w1063, w1064);
  FullAdder U274 (w1064, w975, IN50[1], w1065, w1066);
  FullAdder U275 (w1066, w976, IN51[0], w1067, w1068);
  HalfAdder U276 (w979, IN7[7], Out1[7], w1070);
  FullAdder U277 (w1070, w981, IN8[7], w1071, w1072);
  FullAdder U278 (w1072, w983, IN9[7], w1073, w1074);
  FullAdder U279 (w1074, w985, IN10[7], w1075, w1076);
  FullAdder U280 (w1076, w987, IN11[7], w1077, w1078);
  FullAdder U281 (w1078, w989, IN12[7], w1079, w1080);
  FullAdder U282 (w1080, w991, IN13[7], w1081, w1082);
  FullAdder U283 (w1082, w993, IN14[7], w1083, w1084);
  FullAdder U284 (w1084, w995, IN15[7], w1085, w1086);
  FullAdder U285 (w1086, w997, IN16[7], w1087, w1088);
  FullAdder U286 (w1088, w999, IN17[7], w1089, w1090);
  FullAdder U287 (w1090, w1001, IN18[7], w1091, w1092);
  FullAdder U288 (w1092, w1003, IN19[7], w1093, w1094);
  FullAdder U289 (w1094, w1005, IN20[7], w1095, w1096);
  FullAdder U290 (w1096, w1007, IN21[7], w1097, w1098);
  FullAdder U291 (w1098, w1009, IN22[7], w1099, w1100);
  FullAdder U292 (w1100, w1011, IN23[7], w1101, w1102);
  FullAdder U293 (w1102, w1013, IN24[7], w1103, w1104);
  FullAdder U294 (w1104, w1015, IN25[7], w1105, w1106);
  FullAdder U295 (w1106, w1017, IN26[7], w1107, w1108);
  FullAdder U296 (w1108, w1019, IN27[7], w1109, w1110);
  FullAdder U297 (w1110, w1021, IN28[7], w1111, w1112);
  FullAdder U298 (w1112, w1023, IN29[7], w1113, w1114);
  FullAdder U299 (w1114, w1025, IN30[7], w1115, w1116);
  FullAdder U300 (w1116, w1027, IN31[7], w1117, w1118);
  FullAdder U301 (w1118, w1029, IN32[7], w1119, w1120);
  FullAdder U302 (w1120, w1031, IN33[7], w1121, w1122);
  FullAdder U303 (w1122, w1033, IN34[7], w1123, w1124);
  FullAdder U304 (w1124, w1035, IN35[7], w1125, w1126);
  FullAdder U305 (w1126, w1037, IN36[7], w1127, w1128);
  FullAdder U306 (w1128, w1039, IN37[7], w1129, w1130);
  FullAdder U307 (w1130, w1041, IN38[7], w1131, w1132);
  FullAdder U308 (w1132, w1043, IN39[7], w1133, w1134);
  FullAdder U309 (w1134, w1045, IN40[7], w1135, w1136);
  FullAdder U310 (w1136, w1047, IN41[7], w1137, w1138);
  FullAdder U311 (w1138, w1049, IN42[7], w1139, w1140);
  FullAdder U312 (w1140, w1051, IN43[7], w1141, w1142);
  FullAdder U313 (w1142, w1053, IN44[7], w1143, w1144);
  FullAdder U314 (w1144, w1055, IN45[7], w1145, w1146);
  FullAdder U315 (w1146, w1057, IN46[7], w1147, w1148);
  FullAdder U316 (w1148, w1059, IN47[5], w1149, w1150);
  FullAdder U317 (w1150, w1061, IN48[4], w1151, w1152);
  FullAdder U318 (w1152, w1063, IN49[3], w1153, w1154);
  FullAdder U319 (w1154, w1065, IN50[2], w1155, w1156);
  FullAdder U320 (w1156, w1067, IN51[1], w1157, w1158);
  FullAdder U321 (w1158, w1068, IN52[0], w1159, w1160);
  HalfAdder U322 (w1071, IN8[8], Out1[8], w1162);
  FullAdder U323 (w1162, w1073, IN9[8], w1163, w1164);
  FullAdder U324 (w1164, w1075, IN10[8], w1165, w1166);
  FullAdder U325 (w1166, w1077, IN11[8], w1167, w1168);
  FullAdder U326 (w1168, w1079, IN12[8], w1169, w1170);
  FullAdder U327 (w1170, w1081, IN13[8], w1171, w1172);
  FullAdder U328 (w1172, w1083, IN14[8], w1173, w1174);
  FullAdder U329 (w1174, w1085, IN15[8], w1175, w1176);
  FullAdder U330 (w1176, w1087, IN16[8], w1177, w1178);
  FullAdder U331 (w1178, w1089, IN17[8], w1179, w1180);
  FullAdder U332 (w1180, w1091, IN18[8], w1181, w1182);
  FullAdder U333 (w1182, w1093, IN19[8], w1183, w1184);
  FullAdder U334 (w1184, w1095, IN20[8], w1185, w1186);
  FullAdder U335 (w1186, w1097, IN21[8], w1187, w1188);
  FullAdder U336 (w1188, w1099, IN22[8], w1189, w1190);
  FullAdder U337 (w1190, w1101, IN23[8], w1191, w1192);
  FullAdder U338 (w1192, w1103, IN24[8], w1193, w1194);
  FullAdder U339 (w1194, w1105, IN25[8], w1195, w1196);
  FullAdder U340 (w1196, w1107, IN26[8], w1197, w1198);
  FullAdder U341 (w1198, w1109, IN27[8], w1199, w1200);
  FullAdder U342 (w1200, w1111, IN28[8], w1201, w1202);
  FullAdder U343 (w1202, w1113, IN29[8], w1203, w1204);
  FullAdder U344 (w1204, w1115, IN30[8], w1205, w1206);
  FullAdder U345 (w1206, w1117, IN31[8], w1207, w1208);
  FullAdder U346 (w1208, w1119, IN32[8], w1209, w1210);
  FullAdder U347 (w1210, w1121, IN33[8], w1211, w1212);
  FullAdder U348 (w1212, w1123, IN34[8], w1213, w1214);
  FullAdder U349 (w1214, w1125, IN35[8], w1215, w1216);
  FullAdder U350 (w1216, w1127, IN36[8], w1217, w1218);
  FullAdder U351 (w1218, w1129, IN37[8], w1219, w1220);
  FullAdder U352 (w1220, w1131, IN38[8], w1221, w1222);
  FullAdder U353 (w1222, w1133, IN39[8], w1223, w1224);
  FullAdder U354 (w1224, w1135, IN40[8], w1225, w1226);
  FullAdder U355 (w1226, w1137, IN41[8], w1227, w1228);
  FullAdder U356 (w1228, w1139, IN42[8], w1229, w1230);
  FullAdder U357 (w1230, w1141, IN43[8], w1231, w1232);
  FullAdder U358 (w1232, w1143, IN44[8], w1233, w1234);
  FullAdder U359 (w1234, w1145, IN45[8], w1235, w1236);
  FullAdder U360 (w1236, w1147, IN46[8], w1237, w1238);
  FullAdder U361 (w1238, w1149, IN47[6], w1239, w1240);
  FullAdder U362 (w1240, w1151, IN48[5], w1241, w1242);
  FullAdder U363 (w1242, w1153, IN49[4], w1243, w1244);
  FullAdder U364 (w1244, w1155, IN50[3], w1245, w1246);
  FullAdder U365 (w1246, w1157, IN51[2], w1247, w1248);
  FullAdder U366 (w1248, w1159, IN52[1], w1249, w1250);
  FullAdder U367 (w1250, w1160, IN53[0], w1251, w1252);
  HalfAdder U368 (w1163, IN9[9], Out1[9], w1254);
  FullAdder U369 (w1254, w1165, IN10[9], w1255, w1256);
  FullAdder U370 (w1256, w1167, IN11[9], w1257, w1258);
  FullAdder U371 (w1258, w1169, IN12[9], w1259, w1260);
  FullAdder U372 (w1260, w1171, IN13[9], w1261, w1262);
  FullAdder U373 (w1262, w1173, IN14[9], w1263, w1264);
  FullAdder U374 (w1264, w1175, IN15[9], w1265, w1266);
  FullAdder U375 (w1266, w1177, IN16[9], w1267, w1268);
  FullAdder U376 (w1268, w1179, IN17[9], w1269, w1270);
  FullAdder U377 (w1270, w1181, IN18[9], w1271, w1272);
  FullAdder U378 (w1272, w1183, IN19[9], w1273, w1274);
  FullAdder U379 (w1274, w1185, IN20[9], w1275, w1276);
  FullAdder U380 (w1276, w1187, IN21[9], w1277, w1278);
  FullAdder U381 (w1278, w1189, IN22[9], w1279, w1280);
  FullAdder U382 (w1280, w1191, IN23[9], w1281, w1282);
  FullAdder U383 (w1282, w1193, IN24[9], w1283, w1284);
  FullAdder U384 (w1284, w1195, IN25[9], w1285, w1286);
  FullAdder U385 (w1286, w1197, IN26[9], w1287, w1288);
  FullAdder U386 (w1288, w1199, IN27[9], w1289, w1290);
  FullAdder U387 (w1290, w1201, IN28[9], w1291, w1292);
  FullAdder U388 (w1292, w1203, IN29[9], w1293, w1294);
  FullAdder U389 (w1294, w1205, IN30[9], w1295, w1296);
  FullAdder U390 (w1296, w1207, IN31[9], w1297, w1298);
  FullAdder U391 (w1298, w1209, IN32[9], w1299, w1300);
  FullAdder U392 (w1300, w1211, IN33[9], w1301, w1302);
  FullAdder U393 (w1302, w1213, IN34[9], w1303, w1304);
  FullAdder U394 (w1304, w1215, IN35[9], w1305, w1306);
  FullAdder U395 (w1306, w1217, IN36[9], w1307, w1308);
  FullAdder U396 (w1308, w1219, IN37[9], w1309, w1310);
  FullAdder U397 (w1310, w1221, IN38[9], w1311, w1312);
  FullAdder U398 (w1312, w1223, IN39[9], w1313, w1314);
  FullAdder U399 (w1314, w1225, IN40[9], w1315, w1316);
  FullAdder U400 (w1316, w1227, IN41[9], w1317, w1318);
  FullAdder U401 (w1318, w1229, IN42[9], w1319, w1320);
  FullAdder U402 (w1320, w1231, IN43[9], w1321, w1322);
  FullAdder U403 (w1322, w1233, IN44[9], w1323, w1324);
  FullAdder U404 (w1324, w1235, IN45[9], w1325, w1326);
  FullAdder U405 (w1326, w1237, IN46[9], w1327, w1328);
  FullAdder U406 (w1328, w1239, IN47[7], w1329, w1330);
  FullAdder U407 (w1330, w1241, IN48[6], w1331, w1332);
  FullAdder U408 (w1332, w1243, IN49[5], w1333, w1334);
  FullAdder U409 (w1334, w1245, IN50[4], w1335, w1336);
  FullAdder U410 (w1336, w1247, IN51[3], w1337, w1338);
  FullAdder U411 (w1338, w1249, IN52[2], w1339, w1340);
  FullAdder U412 (w1340, w1251, IN53[1], w1341, w1342);
  FullAdder U413 (w1342, w1252, IN54[0], w1343, w1344);
  HalfAdder U414 (w1255, IN10[10], Out1[10], w1346);
  FullAdder U415 (w1346, w1257, IN11[10], Out1[11], w1348);
  FullAdder U416 (w1348, w1259, IN12[10], Out1[12], w1350);
  FullAdder U417 (w1350, w1261, IN13[10], Out1[13], w1352);
  FullAdder U418 (w1352, w1263, IN14[10], Out1[14], w1354);
  FullAdder U419 (w1354, w1265, IN15[10], Out1[15], w1356);
  FullAdder U420 (w1356, w1267, IN16[10], Out1[16], w1358);
  FullAdder U421 (w1358, w1269, IN17[10], Out1[17], w1360);
  FullAdder U422 (w1360, w1271, IN18[10], Out1[18], w1362);
  FullAdder U423 (w1362, w1273, IN19[10], Out1[19], w1364);
  FullAdder U424 (w1364, w1275, IN20[10], Out1[20], w1366);
  FullAdder U425 (w1366, w1277, IN21[10], Out1[21], w1368);
  FullAdder U426 (w1368, w1279, IN22[10], Out1[22], w1370);
  FullAdder U427 (w1370, w1281, IN23[10], Out1[23], w1372);
  FullAdder U428 (w1372, w1283, IN24[10], Out1[24], w1374);
  FullAdder U429 (w1374, w1285, IN25[10], Out1[25], w1376);
  FullAdder U430 (w1376, w1287, IN26[10], Out1[26], w1378);
  FullAdder U431 (w1378, w1289, IN27[10], Out1[27], w1380);
  FullAdder U432 (w1380, w1291, IN28[10], Out1[28], w1382);
  FullAdder U433 (w1382, w1293, IN29[10], Out1[29], w1384);
  FullAdder U434 (w1384, w1295, IN30[10], Out1[30], w1386);
  FullAdder U435 (w1386, w1297, IN31[10], Out1[31], w1388);
  FullAdder U436 (w1388, w1299, IN32[10], Out1[32], w1390);
  FullAdder U437 (w1390, w1301, IN33[10], Out1[33], w1392);
  FullAdder U438 (w1392, w1303, IN34[10], Out1[34], w1394);
  FullAdder U439 (w1394, w1305, IN35[10], Out1[35], w1396);
  FullAdder U440 (w1396, w1307, IN36[10], Out1[36], w1398);
  FullAdder U441 (w1398, w1309, IN37[10], Out1[37], w1400);
  FullAdder U442 (w1400, w1311, IN38[10], Out1[38], w1402);
  FullAdder U443 (w1402, w1313, IN39[10], Out1[39], w1404);
  FullAdder U444 (w1404, w1315, IN40[10], Out1[40], w1406);
  FullAdder U445 (w1406, w1317, IN41[10], Out1[41], w1408);
  FullAdder U446 (w1408, w1319, IN42[10], Out1[42], w1410);
  FullAdder U447 (w1410, w1321, IN43[10], Out1[43], w1412);
  FullAdder U448 (w1412, w1323, IN44[10], Out1[44], w1414);
  FullAdder U449 (w1414, w1325, IN45[10], Out1[45], w1416);
  FullAdder U450 (w1416, w1327, IN46[10], Out1[46], w1418);
  FullAdder U451 (w1418, w1329, IN47[8], Out1[47], w1420);
  FullAdder U452 (w1420, w1331, IN48[7], Out1[48], w1422);
  FullAdder U453 (w1422, w1333, IN49[6], Out1[49], w1424);
  FullAdder U454 (w1424, w1335, IN50[5], Out1[50], w1426);
  FullAdder U455 (w1426, w1337, IN51[4], Out1[51], w1428);
  FullAdder U456 (w1428, w1339, IN52[3], Out1[52], w1430);
  FullAdder U457 (w1430, w1341, IN53[2], Out1[53], w1432);
  FullAdder U458 (w1432, w1343, IN54[1], Out1[54], w1434);
  FullAdder U459 (w1434, w1344, IN55[0], Out1[55], Out1[56]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN47[9];
  assign Out2[1] = IN48[8];
  assign Out2[2] = IN49[7];
  assign Out2[3] = IN50[6];
  assign Out2[4] = IN51[5];
  assign Out2[5] = IN52[4];
  assign Out2[6] = IN53[3];
  assign Out2[7] = IN54[2];
  assign Out2[8] = IN55[1];
  assign Out2[9] = IN56[0];

endmodule
module RC_10_10(IN1, IN2, Out);
  input [9:0] IN1;
  input [9:0] IN2;
  output [10:0] Out;
  wire w21;
  wire w23;
  wire w25;
  wire w27;
  wire w29;
  wire w31;
  wire w33;
  wire w35;
  wire w37;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w21);
  FullAdder U1 (IN1[1], IN2[1], w21, Out[1], w23);
  FullAdder U2 (IN1[2], IN2[2], w23, Out[2], w25);
  FullAdder U3 (IN1[3], IN2[3], w25, Out[3], w27);
  FullAdder U4 (IN1[4], IN2[4], w27, Out[4], w29);
  FullAdder U5 (IN1[5], IN2[5], w29, Out[5], w31);
  FullAdder U6 (IN1[6], IN2[6], w31, Out[6], w33);
  FullAdder U7 (IN1[7], IN2[7], w33, Out[7], w35);
  FullAdder U8 (IN1[8], IN2[8], w35, Out[8], w37);
  FullAdder U9 (IN1[9], IN2[9], w37, Out[9], Out[10]);

endmodule
module NR_47_11(IN1, IN2, Out);
  input [46:0] IN1;
  input [10:0] IN2;
  output [57:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [10:0] P11;
  wire [10:0] P12;
  wire [10:0] P13;
  wire [10:0] P14;
  wire [10:0] P15;
  wire [10:0] P16;
  wire [10:0] P17;
  wire [10:0] P18;
  wire [10:0] P19;
  wire [10:0] P20;
  wire [10:0] P21;
  wire [10:0] P22;
  wire [10:0] P23;
  wire [10:0] P24;
  wire [10:0] P25;
  wire [10:0] P26;
  wire [10:0] P27;
  wire [10:0] P28;
  wire [10:0] P29;
  wire [10:0] P30;
  wire [10:0] P31;
  wire [10:0] P32;
  wire [10:0] P33;
  wire [10:0] P34;
  wire [10:0] P35;
  wire [10:0] P36;
  wire [10:0] P37;
  wire [10:0] P38;
  wire [10:0] P39;
  wire [10:0] P40;
  wire [10:0] P41;
  wire [10:0] P42;
  wire [10:0] P43;
  wire [10:0] P44;
  wire [10:0] P45;
  wire [10:0] P46;
  wire [9:0] P47;
  wire [8:0] P48;
  wire [7:0] P49;
  wire [6:0] P50;
  wire [5:0] P51;
  wire [4:0] P52;
  wire [3:0] P53;
  wire [2:0] P54;
  wire [1:0] P55;
  wire [0:0] P56;
  wire [56:0] R1;
  wire [9:0] R2;
  wire [57:0] aOut;
  U_SP_47_11 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, R1, R2);
  RC_10_10 S2 (R1[56:47], R2, aOut[57:47]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign Out = aOut[57:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
