
module NR_37_1(
    input [36:0]IN1,
    input [0:0]IN2,
    output [36:0]Out
);
    assign Out = IN2;
endmodule
