//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 51
  second input length: 62
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_51_62(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111);
  input [50:0] IN1;
  input [61:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [29:0] P29;
  output [30:0] P30;
  output [31:0] P31;
  output [32:0] P32;
  output [33:0] P33;
  output [34:0] P34;
  output [35:0] P35;
  output [36:0] P36;
  output [37:0] P37;
  output [38:0] P38;
  output [39:0] P39;
  output [40:0] P40;
  output [41:0] P41;
  output [42:0] P42;
  output [43:0] P43;
  output [44:0] P44;
  output [45:0] P45;
  output [46:0] P46;
  output [47:0] P47;
  output [48:0] P48;
  output [49:0] P49;
  output [50:0] P50;
  output [50:0] P51;
  output [50:0] P52;
  output [50:0] P53;
  output [50:0] P54;
  output [50:0] P55;
  output [50:0] P56;
  output [50:0] P57;
  output [50:0] P58;
  output [50:0] P59;
  output [50:0] P60;
  output [50:0] P61;
  output [49:0] P62;
  output [48:0] P63;
  output [47:0] P64;
  output [46:0] P65;
  output [45:0] P66;
  output [44:0] P67;
  output [43:0] P68;
  output [42:0] P69;
  output [41:0] P70;
  output [40:0] P71;
  output [39:0] P72;
  output [38:0] P73;
  output [37:0] P74;
  output [36:0] P75;
  output [35:0] P76;
  output [34:0] P77;
  output [33:0] P78;
  output [32:0] P79;
  output [31:0] P80;
  output [30:0] P81;
  output [29:0] P82;
  output [28:0] P83;
  output [27:0] P84;
  output [26:0] P85;
  output [25:0] P86;
  output [24:0] P87;
  output [23:0] P88;
  output [22:0] P89;
  output [21:0] P90;
  output [20:0] P91;
  output [19:0] P92;
  output [18:0] P93;
  output [17:0] P94;
  output [16:0] P95;
  output [15:0] P96;
  output [14:0] P97;
  output [13:0] P98;
  output [12:0] P99;
  output [11:0] P100;
  output [10:0] P101;
  output [9:0] P102;
  output [8:0] P103;
  output [7:0] P104;
  output [6:0] P105;
  output [5:0] P106;
  output [4:0] P107;
  output [3:0] P108;
  output [2:0] P109;
  output [1:0] P110;
  output [0:0] P111;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P59[0] = IN1[0]&IN2[59];
  assign P60[0] = IN1[0]&IN2[60];
  assign P61[0] = IN1[0]&IN2[61];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[1] = IN1[1]&IN2[58];
  assign P60[1] = IN1[1]&IN2[59];
  assign P61[1] = IN1[1]&IN2[60];
  assign P62[0] = IN1[1]&IN2[61];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[2] = IN1[2]&IN2[57];
  assign P60[2] = IN1[2]&IN2[58];
  assign P61[2] = IN1[2]&IN2[59];
  assign P62[1] = IN1[2]&IN2[60];
  assign P63[0] = IN1[2]&IN2[61];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[3] = IN1[3]&IN2[56];
  assign P60[3] = IN1[3]&IN2[57];
  assign P61[3] = IN1[3]&IN2[58];
  assign P62[2] = IN1[3]&IN2[59];
  assign P63[1] = IN1[3]&IN2[60];
  assign P64[0] = IN1[3]&IN2[61];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[4] = IN1[4]&IN2[55];
  assign P60[4] = IN1[4]&IN2[56];
  assign P61[4] = IN1[4]&IN2[57];
  assign P62[3] = IN1[4]&IN2[58];
  assign P63[2] = IN1[4]&IN2[59];
  assign P64[1] = IN1[4]&IN2[60];
  assign P65[0] = IN1[4]&IN2[61];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[5] = IN1[5]&IN2[54];
  assign P60[5] = IN1[5]&IN2[55];
  assign P61[5] = IN1[5]&IN2[56];
  assign P62[4] = IN1[5]&IN2[57];
  assign P63[3] = IN1[5]&IN2[58];
  assign P64[2] = IN1[5]&IN2[59];
  assign P65[1] = IN1[5]&IN2[60];
  assign P66[0] = IN1[5]&IN2[61];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[6] = IN1[6]&IN2[53];
  assign P60[6] = IN1[6]&IN2[54];
  assign P61[6] = IN1[6]&IN2[55];
  assign P62[5] = IN1[6]&IN2[56];
  assign P63[4] = IN1[6]&IN2[57];
  assign P64[3] = IN1[6]&IN2[58];
  assign P65[2] = IN1[6]&IN2[59];
  assign P66[1] = IN1[6]&IN2[60];
  assign P67[0] = IN1[6]&IN2[61];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[7] = IN1[7]&IN2[47];
  assign P55[7] = IN1[7]&IN2[48];
  assign P56[7] = IN1[7]&IN2[49];
  assign P57[7] = IN1[7]&IN2[50];
  assign P58[7] = IN1[7]&IN2[51];
  assign P59[7] = IN1[7]&IN2[52];
  assign P60[7] = IN1[7]&IN2[53];
  assign P61[7] = IN1[7]&IN2[54];
  assign P62[6] = IN1[7]&IN2[55];
  assign P63[5] = IN1[7]&IN2[56];
  assign P64[4] = IN1[7]&IN2[57];
  assign P65[3] = IN1[7]&IN2[58];
  assign P66[2] = IN1[7]&IN2[59];
  assign P67[1] = IN1[7]&IN2[60];
  assign P68[0] = IN1[7]&IN2[61];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[8] = IN1[8]&IN2[45];
  assign P54[8] = IN1[8]&IN2[46];
  assign P55[8] = IN1[8]&IN2[47];
  assign P56[8] = IN1[8]&IN2[48];
  assign P57[8] = IN1[8]&IN2[49];
  assign P58[8] = IN1[8]&IN2[50];
  assign P59[8] = IN1[8]&IN2[51];
  assign P60[8] = IN1[8]&IN2[52];
  assign P61[8] = IN1[8]&IN2[53];
  assign P62[7] = IN1[8]&IN2[54];
  assign P63[6] = IN1[8]&IN2[55];
  assign P64[5] = IN1[8]&IN2[56];
  assign P65[4] = IN1[8]&IN2[57];
  assign P66[3] = IN1[8]&IN2[58];
  assign P67[2] = IN1[8]&IN2[59];
  assign P68[1] = IN1[8]&IN2[60];
  assign P69[0] = IN1[8]&IN2[61];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[9] = IN1[9]&IN2[44];
  assign P54[9] = IN1[9]&IN2[45];
  assign P55[9] = IN1[9]&IN2[46];
  assign P56[9] = IN1[9]&IN2[47];
  assign P57[9] = IN1[9]&IN2[48];
  assign P58[9] = IN1[9]&IN2[49];
  assign P59[9] = IN1[9]&IN2[50];
  assign P60[9] = IN1[9]&IN2[51];
  assign P61[9] = IN1[9]&IN2[52];
  assign P62[8] = IN1[9]&IN2[53];
  assign P63[7] = IN1[9]&IN2[54];
  assign P64[6] = IN1[9]&IN2[55];
  assign P65[5] = IN1[9]&IN2[56];
  assign P66[4] = IN1[9]&IN2[57];
  assign P67[3] = IN1[9]&IN2[58];
  assign P68[2] = IN1[9]&IN2[59];
  assign P69[1] = IN1[9]&IN2[60];
  assign P70[0] = IN1[9]&IN2[61];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[10] = IN1[10]&IN2[39];
  assign P50[10] = IN1[10]&IN2[40];
  assign P51[10] = IN1[10]&IN2[41];
  assign P52[10] = IN1[10]&IN2[42];
  assign P53[10] = IN1[10]&IN2[43];
  assign P54[10] = IN1[10]&IN2[44];
  assign P55[10] = IN1[10]&IN2[45];
  assign P56[10] = IN1[10]&IN2[46];
  assign P57[10] = IN1[10]&IN2[47];
  assign P58[10] = IN1[10]&IN2[48];
  assign P59[10] = IN1[10]&IN2[49];
  assign P60[10] = IN1[10]&IN2[50];
  assign P61[10] = IN1[10]&IN2[51];
  assign P62[9] = IN1[10]&IN2[52];
  assign P63[8] = IN1[10]&IN2[53];
  assign P64[7] = IN1[10]&IN2[54];
  assign P65[6] = IN1[10]&IN2[55];
  assign P66[5] = IN1[10]&IN2[56];
  assign P67[4] = IN1[10]&IN2[57];
  assign P68[3] = IN1[10]&IN2[58];
  assign P69[2] = IN1[10]&IN2[59];
  assign P70[1] = IN1[10]&IN2[60];
  assign P71[0] = IN1[10]&IN2[61];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[11] = IN1[11]&IN2[38];
  assign P50[11] = IN1[11]&IN2[39];
  assign P51[11] = IN1[11]&IN2[40];
  assign P52[11] = IN1[11]&IN2[41];
  assign P53[11] = IN1[11]&IN2[42];
  assign P54[11] = IN1[11]&IN2[43];
  assign P55[11] = IN1[11]&IN2[44];
  assign P56[11] = IN1[11]&IN2[45];
  assign P57[11] = IN1[11]&IN2[46];
  assign P58[11] = IN1[11]&IN2[47];
  assign P59[11] = IN1[11]&IN2[48];
  assign P60[11] = IN1[11]&IN2[49];
  assign P61[11] = IN1[11]&IN2[50];
  assign P62[10] = IN1[11]&IN2[51];
  assign P63[9] = IN1[11]&IN2[52];
  assign P64[8] = IN1[11]&IN2[53];
  assign P65[7] = IN1[11]&IN2[54];
  assign P66[6] = IN1[11]&IN2[55];
  assign P67[5] = IN1[11]&IN2[56];
  assign P68[4] = IN1[11]&IN2[57];
  assign P69[3] = IN1[11]&IN2[58];
  assign P70[2] = IN1[11]&IN2[59];
  assign P71[1] = IN1[11]&IN2[60];
  assign P72[0] = IN1[11]&IN2[61];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[12] = IN1[12]&IN2[37];
  assign P50[12] = IN1[12]&IN2[38];
  assign P51[12] = IN1[12]&IN2[39];
  assign P52[12] = IN1[12]&IN2[40];
  assign P53[12] = IN1[12]&IN2[41];
  assign P54[12] = IN1[12]&IN2[42];
  assign P55[12] = IN1[12]&IN2[43];
  assign P56[12] = IN1[12]&IN2[44];
  assign P57[12] = IN1[12]&IN2[45];
  assign P58[12] = IN1[12]&IN2[46];
  assign P59[12] = IN1[12]&IN2[47];
  assign P60[12] = IN1[12]&IN2[48];
  assign P61[12] = IN1[12]&IN2[49];
  assign P62[11] = IN1[12]&IN2[50];
  assign P63[10] = IN1[12]&IN2[51];
  assign P64[9] = IN1[12]&IN2[52];
  assign P65[8] = IN1[12]&IN2[53];
  assign P66[7] = IN1[12]&IN2[54];
  assign P67[6] = IN1[12]&IN2[55];
  assign P68[5] = IN1[12]&IN2[56];
  assign P69[4] = IN1[12]&IN2[57];
  assign P70[3] = IN1[12]&IN2[58];
  assign P71[2] = IN1[12]&IN2[59];
  assign P72[1] = IN1[12]&IN2[60];
  assign P73[0] = IN1[12]&IN2[61];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[13] = IN1[13]&IN2[36];
  assign P50[13] = IN1[13]&IN2[37];
  assign P51[13] = IN1[13]&IN2[38];
  assign P52[13] = IN1[13]&IN2[39];
  assign P53[13] = IN1[13]&IN2[40];
  assign P54[13] = IN1[13]&IN2[41];
  assign P55[13] = IN1[13]&IN2[42];
  assign P56[13] = IN1[13]&IN2[43];
  assign P57[13] = IN1[13]&IN2[44];
  assign P58[13] = IN1[13]&IN2[45];
  assign P59[13] = IN1[13]&IN2[46];
  assign P60[13] = IN1[13]&IN2[47];
  assign P61[13] = IN1[13]&IN2[48];
  assign P62[12] = IN1[13]&IN2[49];
  assign P63[11] = IN1[13]&IN2[50];
  assign P64[10] = IN1[13]&IN2[51];
  assign P65[9] = IN1[13]&IN2[52];
  assign P66[8] = IN1[13]&IN2[53];
  assign P67[7] = IN1[13]&IN2[54];
  assign P68[6] = IN1[13]&IN2[55];
  assign P69[5] = IN1[13]&IN2[56];
  assign P70[4] = IN1[13]&IN2[57];
  assign P71[3] = IN1[13]&IN2[58];
  assign P72[2] = IN1[13]&IN2[59];
  assign P73[1] = IN1[13]&IN2[60];
  assign P74[0] = IN1[13]&IN2[61];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[14] = IN1[14]&IN2[24];
  assign P39[14] = IN1[14]&IN2[25];
  assign P40[14] = IN1[14]&IN2[26];
  assign P41[14] = IN1[14]&IN2[27];
  assign P42[14] = IN1[14]&IN2[28];
  assign P43[14] = IN1[14]&IN2[29];
  assign P44[14] = IN1[14]&IN2[30];
  assign P45[14] = IN1[14]&IN2[31];
  assign P46[14] = IN1[14]&IN2[32];
  assign P47[14] = IN1[14]&IN2[33];
  assign P48[14] = IN1[14]&IN2[34];
  assign P49[14] = IN1[14]&IN2[35];
  assign P50[14] = IN1[14]&IN2[36];
  assign P51[14] = IN1[14]&IN2[37];
  assign P52[14] = IN1[14]&IN2[38];
  assign P53[14] = IN1[14]&IN2[39];
  assign P54[14] = IN1[14]&IN2[40];
  assign P55[14] = IN1[14]&IN2[41];
  assign P56[14] = IN1[14]&IN2[42];
  assign P57[14] = IN1[14]&IN2[43];
  assign P58[14] = IN1[14]&IN2[44];
  assign P59[14] = IN1[14]&IN2[45];
  assign P60[14] = IN1[14]&IN2[46];
  assign P61[14] = IN1[14]&IN2[47];
  assign P62[13] = IN1[14]&IN2[48];
  assign P63[12] = IN1[14]&IN2[49];
  assign P64[11] = IN1[14]&IN2[50];
  assign P65[10] = IN1[14]&IN2[51];
  assign P66[9] = IN1[14]&IN2[52];
  assign P67[8] = IN1[14]&IN2[53];
  assign P68[7] = IN1[14]&IN2[54];
  assign P69[6] = IN1[14]&IN2[55];
  assign P70[5] = IN1[14]&IN2[56];
  assign P71[4] = IN1[14]&IN2[57];
  assign P72[3] = IN1[14]&IN2[58];
  assign P73[2] = IN1[14]&IN2[59];
  assign P74[1] = IN1[14]&IN2[60];
  assign P75[0] = IN1[14]&IN2[61];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[15] = IN1[15]&IN2[23];
  assign P39[15] = IN1[15]&IN2[24];
  assign P40[15] = IN1[15]&IN2[25];
  assign P41[15] = IN1[15]&IN2[26];
  assign P42[15] = IN1[15]&IN2[27];
  assign P43[15] = IN1[15]&IN2[28];
  assign P44[15] = IN1[15]&IN2[29];
  assign P45[15] = IN1[15]&IN2[30];
  assign P46[15] = IN1[15]&IN2[31];
  assign P47[15] = IN1[15]&IN2[32];
  assign P48[15] = IN1[15]&IN2[33];
  assign P49[15] = IN1[15]&IN2[34];
  assign P50[15] = IN1[15]&IN2[35];
  assign P51[15] = IN1[15]&IN2[36];
  assign P52[15] = IN1[15]&IN2[37];
  assign P53[15] = IN1[15]&IN2[38];
  assign P54[15] = IN1[15]&IN2[39];
  assign P55[15] = IN1[15]&IN2[40];
  assign P56[15] = IN1[15]&IN2[41];
  assign P57[15] = IN1[15]&IN2[42];
  assign P58[15] = IN1[15]&IN2[43];
  assign P59[15] = IN1[15]&IN2[44];
  assign P60[15] = IN1[15]&IN2[45];
  assign P61[15] = IN1[15]&IN2[46];
  assign P62[14] = IN1[15]&IN2[47];
  assign P63[13] = IN1[15]&IN2[48];
  assign P64[12] = IN1[15]&IN2[49];
  assign P65[11] = IN1[15]&IN2[50];
  assign P66[10] = IN1[15]&IN2[51];
  assign P67[9] = IN1[15]&IN2[52];
  assign P68[8] = IN1[15]&IN2[53];
  assign P69[7] = IN1[15]&IN2[54];
  assign P70[6] = IN1[15]&IN2[55];
  assign P71[5] = IN1[15]&IN2[56];
  assign P72[4] = IN1[15]&IN2[57];
  assign P73[3] = IN1[15]&IN2[58];
  assign P74[2] = IN1[15]&IN2[59];
  assign P75[1] = IN1[15]&IN2[60];
  assign P76[0] = IN1[15]&IN2[61];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[16] = IN1[16]&IN2[22];
  assign P39[16] = IN1[16]&IN2[23];
  assign P40[16] = IN1[16]&IN2[24];
  assign P41[16] = IN1[16]&IN2[25];
  assign P42[16] = IN1[16]&IN2[26];
  assign P43[16] = IN1[16]&IN2[27];
  assign P44[16] = IN1[16]&IN2[28];
  assign P45[16] = IN1[16]&IN2[29];
  assign P46[16] = IN1[16]&IN2[30];
  assign P47[16] = IN1[16]&IN2[31];
  assign P48[16] = IN1[16]&IN2[32];
  assign P49[16] = IN1[16]&IN2[33];
  assign P50[16] = IN1[16]&IN2[34];
  assign P51[16] = IN1[16]&IN2[35];
  assign P52[16] = IN1[16]&IN2[36];
  assign P53[16] = IN1[16]&IN2[37];
  assign P54[16] = IN1[16]&IN2[38];
  assign P55[16] = IN1[16]&IN2[39];
  assign P56[16] = IN1[16]&IN2[40];
  assign P57[16] = IN1[16]&IN2[41];
  assign P58[16] = IN1[16]&IN2[42];
  assign P59[16] = IN1[16]&IN2[43];
  assign P60[16] = IN1[16]&IN2[44];
  assign P61[16] = IN1[16]&IN2[45];
  assign P62[15] = IN1[16]&IN2[46];
  assign P63[14] = IN1[16]&IN2[47];
  assign P64[13] = IN1[16]&IN2[48];
  assign P65[12] = IN1[16]&IN2[49];
  assign P66[11] = IN1[16]&IN2[50];
  assign P67[10] = IN1[16]&IN2[51];
  assign P68[9] = IN1[16]&IN2[52];
  assign P69[8] = IN1[16]&IN2[53];
  assign P70[7] = IN1[16]&IN2[54];
  assign P71[6] = IN1[16]&IN2[55];
  assign P72[5] = IN1[16]&IN2[56];
  assign P73[4] = IN1[16]&IN2[57];
  assign P74[3] = IN1[16]&IN2[58];
  assign P75[2] = IN1[16]&IN2[59];
  assign P76[1] = IN1[16]&IN2[60];
  assign P77[0] = IN1[16]&IN2[61];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[17] = IN1[17]&IN2[21];
  assign P39[17] = IN1[17]&IN2[22];
  assign P40[17] = IN1[17]&IN2[23];
  assign P41[17] = IN1[17]&IN2[24];
  assign P42[17] = IN1[17]&IN2[25];
  assign P43[17] = IN1[17]&IN2[26];
  assign P44[17] = IN1[17]&IN2[27];
  assign P45[17] = IN1[17]&IN2[28];
  assign P46[17] = IN1[17]&IN2[29];
  assign P47[17] = IN1[17]&IN2[30];
  assign P48[17] = IN1[17]&IN2[31];
  assign P49[17] = IN1[17]&IN2[32];
  assign P50[17] = IN1[17]&IN2[33];
  assign P51[17] = IN1[17]&IN2[34];
  assign P52[17] = IN1[17]&IN2[35];
  assign P53[17] = IN1[17]&IN2[36];
  assign P54[17] = IN1[17]&IN2[37];
  assign P55[17] = IN1[17]&IN2[38];
  assign P56[17] = IN1[17]&IN2[39];
  assign P57[17] = IN1[17]&IN2[40];
  assign P58[17] = IN1[17]&IN2[41];
  assign P59[17] = IN1[17]&IN2[42];
  assign P60[17] = IN1[17]&IN2[43];
  assign P61[17] = IN1[17]&IN2[44];
  assign P62[16] = IN1[17]&IN2[45];
  assign P63[15] = IN1[17]&IN2[46];
  assign P64[14] = IN1[17]&IN2[47];
  assign P65[13] = IN1[17]&IN2[48];
  assign P66[12] = IN1[17]&IN2[49];
  assign P67[11] = IN1[17]&IN2[50];
  assign P68[10] = IN1[17]&IN2[51];
  assign P69[9] = IN1[17]&IN2[52];
  assign P70[8] = IN1[17]&IN2[53];
  assign P71[7] = IN1[17]&IN2[54];
  assign P72[6] = IN1[17]&IN2[55];
  assign P73[5] = IN1[17]&IN2[56];
  assign P74[4] = IN1[17]&IN2[57];
  assign P75[3] = IN1[17]&IN2[58];
  assign P76[2] = IN1[17]&IN2[59];
  assign P77[1] = IN1[17]&IN2[60];
  assign P78[0] = IN1[17]&IN2[61];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[18] = IN1[18]&IN2[20];
  assign P39[18] = IN1[18]&IN2[21];
  assign P40[18] = IN1[18]&IN2[22];
  assign P41[18] = IN1[18]&IN2[23];
  assign P42[18] = IN1[18]&IN2[24];
  assign P43[18] = IN1[18]&IN2[25];
  assign P44[18] = IN1[18]&IN2[26];
  assign P45[18] = IN1[18]&IN2[27];
  assign P46[18] = IN1[18]&IN2[28];
  assign P47[18] = IN1[18]&IN2[29];
  assign P48[18] = IN1[18]&IN2[30];
  assign P49[18] = IN1[18]&IN2[31];
  assign P50[18] = IN1[18]&IN2[32];
  assign P51[18] = IN1[18]&IN2[33];
  assign P52[18] = IN1[18]&IN2[34];
  assign P53[18] = IN1[18]&IN2[35];
  assign P54[18] = IN1[18]&IN2[36];
  assign P55[18] = IN1[18]&IN2[37];
  assign P56[18] = IN1[18]&IN2[38];
  assign P57[18] = IN1[18]&IN2[39];
  assign P58[18] = IN1[18]&IN2[40];
  assign P59[18] = IN1[18]&IN2[41];
  assign P60[18] = IN1[18]&IN2[42];
  assign P61[18] = IN1[18]&IN2[43];
  assign P62[17] = IN1[18]&IN2[44];
  assign P63[16] = IN1[18]&IN2[45];
  assign P64[15] = IN1[18]&IN2[46];
  assign P65[14] = IN1[18]&IN2[47];
  assign P66[13] = IN1[18]&IN2[48];
  assign P67[12] = IN1[18]&IN2[49];
  assign P68[11] = IN1[18]&IN2[50];
  assign P69[10] = IN1[18]&IN2[51];
  assign P70[9] = IN1[18]&IN2[52];
  assign P71[8] = IN1[18]&IN2[53];
  assign P72[7] = IN1[18]&IN2[54];
  assign P73[6] = IN1[18]&IN2[55];
  assign P74[5] = IN1[18]&IN2[56];
  assign P75[4] = IN1[18]&IN2[57];
  assign P76[3] = IN1[18]&IN2[58];
  assign P77[2] = IN1[18]&IN2[59];
  assign P78[1] = IN1[18]&IN2[60];
  assign P79[0] = IN1[18]&IN2[61];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[19] = IN1[19]&IN2[19];
  assign P39[19] = IN1[19]&IN2[20];
  assign P40[19] = IN1[19]&IN2[21];
  assign P41[19] = IN1[19]&IN2[22];
  assign P42[19] = IN1[19]&IN2[23];
  assign P43[19] = IN1[19]&IN2[24];
  assign P44[19] = IN1[19]&IN2[25];
  assign P45[19] = IN1[19]&IN2[26];
  assign P46[19] = IN1[19]&IN2[27];
  assign P47[19] = IN1[19]&IN2[28];
  assign P48[19] = IN1[19]&IN2[29];
  assign P49[19] = IN1[19]&IN2[30];
  assign P50[19] = IN1[19]&IN2[31];
  assign P51[19] = IN1[19]&IN2[32];
  assign P52[19] = IN1[19]&IN2[33];
  assign P53[19] = IN1[19]&IN2[34];
  assign P54[19] = IN1[19]&IN2[35];
  assign P55[19] = IN1[19]&IN2[36];
  assign P56[19] = IN1[19]&IN2[37];
  assign P57[19] = IN1[19]&IN2[38];
  assign P58[19] = IN1[19]&IN2[39];
  assign P59[19] = IN1[19]&IN2[40];
  assign P60[19] = IN1[19]&IN2[41];
  assign P61[19] = IN1[19]&IN2[42];
  assign P62[18] = IN1[19]&IN2[43];
  assign P63[17] = IN1[19]&IN2[44];
  assign P64[16] = IN1[19]&IN2[45];
  assign P65[15] = IN1[19]&IN2[46];
  assign P66[14] = IN1[19]&IN2[47];
  assign P67[13] = IN1[19]&IN2[48];
  assign P68[12] = IN1[19]&IN2[49];
  assign P69[11] = IN1[19]&IN2[50];
  assign P70[10] = IN1[19]&IN2[51];
  assign P71[9] = IN1[19]&IN2[52];
  assign P72[8] = IN1[19]&IN2[53];
  assign P73[7] = IN1[19]&IN2[54];
  assign P74[6] = IN1[19]&IN2[55];
  assign P75[5] = IN1[19]&IN2[56];
  assign P76[4] = IN1[19]&IN2[57];
  assign P77[3] = IN1[19]&IN2[58];
  assign P78[2] = IN1[19]&IN2[59];
  assign P79[1] = IN1[19]&IN2[60];
  assign P80[0] = IN1[19]&IN2[61];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[20] = IN1[20]&IN2[18];
  assign P39[20] = IN1[20]&IN2[19];
  assign P40[20] = IN1[20]&IN2[20];
  assign P41[20] = IN1[20]&IN2[21];
  assign P42[20] = IN1[20]&IN2[22];
  assign P43[20] = IN1[20]&IN2[23];
  assign P44[20] = IN1[20]&IN2[24];
  assign P45[20] = IN1[20]&IN2[25];
  assign P46[20] = IN1[20]&IN2[26];
  assign P47[20] = IN1[20]&IN2[27];
  assign P48[20] = IN1[20]&IN2[28];
  assign P49[20] = IN1[20]&IN2[29];
  assign P50[20] = IN1[20]&IN2[30];
  assign P51[20] = IN1[20]&IN2[31];
  assign P52[20] = IN1[20]&IN2[32];
  assign P53[20] = IN1[20]&IN2[33];
  assign P54[20] = IN1[20]&IN2[34];
  assign P55[20] = IN1[20]&IN2[35];
  assign P56[20] = IN1[20]&IN2[36];
  assign P57[20] = IN1[20]&IN2[37];
  assign P58[20] = IN1[20]&IN2[38];
  assign P59[20] = IN1[20]&IN2[39];
  assign P60[20] = IN1[20]&IN2[40];
  assign P61[20] = IN1[20]&IN2[41];
  assign P62[19] = IN1[20]&IN2[42];
  assign P63[18] = IN1[20]&IN2[43];
  assign P64[17] = IN1[20]&IN2[44];
  assign P65[16] = IN1[20]&IN2[45];
  assign P66[15] = IN1[20]&IN2[46];
  assign P67[14] = IN1[20]&IN2[47];
  assign P68[13] = IN1[20]&IN2[48];
  assign P69[12] = IN1[20]&IN2[49];
  assign P70[11] = IN1[20]&IN2[50];
  assign P71[10] = IN1[20]&IN2[51];
  assign P72[9] = IN1[20]&IN2[52];
  assign P73[8] = IN1[20]&IN2[53];
  assign P74[7] = IN1[20]&IN2[54];
  assign P75[6] = IN1[20]&IN2[55];
  assign P76[5] = IN1[20]&IN2[56];
  assign P77[4] = IN1[20]&IN2[57];
  assign P78[3] = IN1[20]&IN2[58];
  assign P79[2] = IN1[20]&IN2[59];
  assign P80[1] = IN1[20]&IN2[60];
  assign P81[0] = IN1[20]&IN2[61];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[21] = IN1[21]&IN2[14];
  assign P36[21] = IN1[21]&IN2[15];
  assign P37[21] = IN1[21]&IN2[16];
  assign P38[21] = IN1[21]&IN2[17];
  assign P39[21] = IN1[21]&IN2[18];
  assign P40[21] = IN1[21]&IN2[19];
  assign P41[21] = IN1[21]&IN2[20];
  assign P42[21] = IN1[21]&IN2[21];
  assign P43[21] = IN1[21]&IN2[22];
  assign P44[21] = IN1[21]&IN2[23];
  assign P45[21] = IN1[21]&IN2[24];
  assign P46[21] = IN1[21]&IN2[25];
  assign P47[21] = IN1[21]&IN2[26];
  assign P48[21] = IN1[21]&IN2[27];
  assign P49[21] = IN1[21]&IN2[28];
  assign P50[21] = IN1[21]&IN2[29];
  assign P51[21] = IN1[21]&IN2[30];
  assign P52[21] = IN1[21]&IN2[31];
  assign P53[21] = IN1[21]&IN2[32];
  assign P54[21] = IN1[21]&IN2[33];
  assign P55[21] = IN1[21]&IN2[34];
  assign P56[21] = IN1[21]&IN2[35];
  assign P57[21] = IN1[21]&IN2[36];
  assign P58[21] = IN1[21]&IN2[37];
  assign P59[21] = IN1[21]&IN2[38];
  assign P60[21] = IN1[21]&IN2[39];
  assign P61[21] = IN1[21]&IN2[40];
  assign P62[20] = IN1[21]&IN2[41];
  assign P63[19] = IN1[21]&IN2[42];
  assign P64[18] = IN1[21]&IN2[43];
  assign P65[17] = IN1[21]&IN2[44];
  assign P66[16] = IN1[21]&IN2[45];
  assign P67[15] = IN1[21]&IN2[46];
  assign P68[14] = IN1[21]&IN2[47];
  assign P69[13] = IN1[21]&IN2[48];
  assign P70[12] = IN1[21]&IN2[49];
  assign P71[11] = IN1[21]&IN2[50];
  assign P72[10] = IN1[21]&IN2[51];
  assign P73[9] = IN1[21]&IN2[52];
  assign P74[8] = IN1[21]&IN2[53];
  assign P75[7] = IN1[21]&IN2[54];
  assign P76[6] = IN1[21]&IN2[55];
  assign P77[5] = IN1[21]&IN2[56];
  assign P78[4] = IN1[21]&IN2[57];
  assign P79[3] = IN1[21]&IN2[58];
  assign P80[2] = IN1[21]&IN2[59];
  assign P81[1] = IN1[21]&IN2[60];
  assign P82[0] = IN1[21]&IN2[61];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[22] = IN1[22]&IN2[13];
  assign P36[22] = IN1[22]&IN2[14];
  assign P37[22] = IN1[22]&IN2[15];
  assign P38[22] = IN1[22]&IN2[16];
  assign P39[22] = IN1[22]&IN2[17];
  assign P40[22] = IN1[22]&IN2[18];
  assign P41[22] = IN1[22]&IN2[19];
  assign P42[22] = IN1[22]&IN2[20];
  assign P43[22] = IN1[22]&IN2[21];
  assign P44[22] = IN1[22]&IN2[22];
  assign P45[22] = IN1[22]&IN2[23];
  assign P46[22] = IN1[22]&IN2[24];
  assign P47[22] = IN1[22]&IN2[25];
  assign P48[22] = IN1[22]&IN2[26];
  assign P49[22] = IN1[22]&IN2[27];
  assign P50[22] = IN1[22]&IN2[28];
  assign P51[22] = IN1[22]&IN2[29];
  assign P52[22] = IN1[22]&IN2[30];
  assign P53[22] = IN1[22]&IN2[31];
  assign P54[22] = IN1[22]&IN2[32];
  assign P55[22] = IN1[22]&IN2[33];
  assign P56[22] = IN1[22]&IN2[34];
  assign P57[22] = IN1[22]&IN2[35];
  assign P58[22] = IN1[22]&IN2[36];
  assign P59[22] = IN1[22]&IN2[37];
  assign P60[22] = IN1[22]&IN2[38];
  assign P61[22] = IN1[22]&IN2[39];
  assign P62[21] = IN1[22]&IN2[40];
  assign P63[20] = IN1[22]&IN2[41];
  assign P64[19] = IN1[22]&IN2[42];
  assign P65[18] = IN1[22]&IN2[43];
  assign P66[17] = IN1[22]&IN2[44];
  assign P67[16] = IN1[22]&IN2[45];
  assign P68[15] = IN1[22]&IN2[46];
  assign P69[14] = IN1[22]&IN2[47];
  assign P70[13] = IN1[22]&IN2[48];
  assign P71[12] = IN1[22]&IN2[49];
  assign P72[11] = IN1[22]&IN2[50];
  assign P73[10] = IN1[22]&IN2[51];
  assign P74[9] = IN1[22]&IN2[52];
  assign P75[8] = IN1[22]&IN2[53];
  assign P76[7] = IN1[22]&IN2[54];
  assign P77[6] = IN1[22]&IN2[55];
  assign P78[5] = IN1[22]&IN2[56];
  assign P79[4] = IN1[22]&IN2[57];
  assign P80[3] = IN1[22]&IN2[58];
  assign P81[2] = IN1[22]&IN2[59];
  assign P82[1] = IN1[22]&IN2[60];
  assign P83[0] = IN1[22]&IN2[61];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[23] = IN1[23]&IN2[12];
  assign P36[23] = IN1[23]&IN2[13];
  assign P37[23] = IN1[23]&IN2[14];
  assign P38[23] = IN1[23]&IN2[15];
  assign P39[23] = IN1[23]&IN2[16];
  assign P40[23] = IN1[23]&IN2[17];
  assign P41[23] = IN1[23]&IN2[18];
  assign P42[23] = IN1[23]&IN2[19];
  assign P43[23] = IN1[23]&IN2[20];
  assign P44[23] = IN1[23]&IN2[21];
  assign P45[23] = IN1[23]&IN2[22];
  assign P46[23] = IN1[23]&IN2[23];
  assign P47[23] = IN1[23]&IN2[24];
  assign P48[23] = IN1[23]&IN2[25];
  assign P49[23] = IN1[23]&IN2[26];
  assign P50[23] = IN1[23]&IN2[27];
  assign P51[23] = IN1[23]&IN2[28];
  assign P52[23] = IN1[23]&IN2[29];
  assign P53[23] = IN1[23]&IN2[30];
  assign P54[23] = IN1[23]&IN2[31];
  assign P55[23] = IN1[23]&IN2[32];
  assign P56[23] = IN1[23]&IN2[33];
  assign P57[23] = IN1[23]&IN2[34];
  assign P58[23] = IN1[23]&IN2[35];
  assign P59[23] = IN1[23]&IN2[36];
  assign P60[23] = IN1[23]&IN2[37];
  assign P61[23] = IN1[23]&IN2[38];
  assign P62[22] = IN1[23]&IN2[39];
  assign P63[21] = IN1[23]&IN2[40];
  assign P64[20] = IN1[23]&IN2[41];
  assign P65[19] = IN1[23]&IN2[42];
  assign P66[18] = IN1[23]&IN2[43];
  assign P67[17] = IN1[23]&IN2[44];
  assign P68[16] = IN1[23]&IN2[45];
  assign P69[15] = IN1[23]&IN2[46];
  assign P70[14] = IN1[23]&IN2[47];
  assign P71[13] = IN1[23]&IN2[48];
  assign P72[12] = IN1[23]&IN2[49];
  assign P73[11] = IN1[23]&IN2[50];
  assign P74[10] = IN1[23]&IN2[51];
  assign P75[9] = IN1[23]&IN2[52];
  assign P76[8] = IN1[23]&IN2[53];
  assign P77[7] = IN1[23]&IN2[54];
  assign P78[6] = IN1[23]&IN2[55];
  assign P79[5] = IN1[23]&IN2[56];
  assign P80[4] = IN1[23]&IN2[57];
  assign P81[3] = IN1[23]&IN2[58];
  assign P82[2] = IN1[23]&IN2[59];
  assign P83[1] = IN1[23]&IN2[60];
  assign P84[0] = IN1[23]&IN2[61];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[24] = IN1[24]&IN2[11];
  assign P36[24] = IN1[24]&IN2[12];
  assign P37[24] = IN1[24]&IN2[13];
  assign P38[24] = IN1[24]&IN2[14];
  assign P39[24] = IN1[24]&IN2[15];
  assign P40[24] = IN1[24]&IN2[16];
  assign P41[24] = IN1[24]&IN2[17];
  assign P42[24] = IN1[24]&IN2[18];
  assign P43[24] = IN1[24]&IN2[19];
  assign P44[24] = IN1[24]&IN2[20];
  assign P45[24] = IN1[24]&IN2[21];
  assign P46[24] = IN1[24]&IN2[22];
  assign P47[24] = IN1[24]&IN2[23];
  assign P48[24] = IN1[24]&IN2[24];
  assign P49[24] = IN1[24]&IN2[25];
  assign P50[24] = IN1[24]&IN2[26];
  assign P51[24] = IN1[24]&IN2[27];
  assign P52[24] = IN1[24]&IN2[28];
  assign P53[24] = IN1[24]&IN2[29];
  assign P54[24] = IN1[24]&IN2[30];
  assign P55[24] = IN1[24]&IN2[31];
  assign P56[24] = IN1[24]&IN2[32];
  assign P57[24] = IN1[24]&IN2[33];
  assign P58[24] = IN1[24]&IN2[34];
  assign P59[24] = IN1[24]&IN2[35];
  assign P60[24] = IN1[24]&IN2[36];
  assign P61[24] = IN1[24]&IN2[37];
  assign P62[23] = IN1[24]&IN2[38];
  assign P63[22] = IN1[24]&IN2[39];
  assign P64[21] = IN1[24]&IN2[40];
  assign P65[20] = IN1[24]&IN2[41];
  assign P66[19] = IN1[24]&IN2[42];
  assign P67[18] = IN1[24]&IN2[43];
  assign P68[17] = IN1[24]&IN2[44];
  assign P69[16] = IN1[24]&IN2[45];
  assign P70[15] = IN1[24]&IN2[46];
  assign P71[14] = IN1[24]&IN2[47];
  assign P72[13] = IN1[24]&IN2[48];
  assign P73[12] = IN1[24]&IN2[49];
  assign P74[11] = IN1[24]&IN2[50];
  assign P75[10] = IN1[24]&IN2[51];
  assign P76[9] = IN1[24]&IN2[52];
  assign P77[8] = IN1[24]&IN2[53];
  assign P78[7] = IN1[24]&IN2[54];
  assign P79[6] = IN1[24]&IN2[55];
  assign P80[5] = IN1[24]&IN2[56];
  assign P81[4] = IN1[24]&IN2[57];
  assign P82[3] = IN1[24]&IN2[58];
  assign P83[2] = IN1[24]&IN2[59];
  assign P84[1] = IN1[24]&IN2[60];
  assign P85[0] = IN1[24]&IN2[61];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[25] = IN1[25]&IN2[10];
  assign P36[25] = IN1[25]&IN2[11];
  assign P37[25] = IN1[25]&IN2[12];
  assign P38[25] = IN1[25]&IN2[13];
  assign P39[25] = IN1[25]&IN2[14];
  assign P40[25] = IN1[25]&IN2[15];
  assign P41[25] = IN1[25]&IN2[16];
  assign P42[25] = IN1[25]&IN2[17];
  assign P43[25] = IN1[25]&IN2[18];
  assign P44[25] = IN1[25]&IN2[19];
  assign P45[25] = IN1[25]&IN2[20];
  assign P46[25] = IN1[25]&IN2[21];
  assign P47[25] = IN1[25]&IN2[22];
  assign P48[25] = IN1[25]&IN2[23];
  assign P49[25] = IN1[25]&IN2[24];
  assign P50[25] = IN1[25]&IN2[25];
  assign P51[25] = IN1[25]&IN2[26];
  assign P52[25] = IN1[25]&IN2[27];
  assign P53[25] = IN1[25]&IN2[28];
  assign P54[25] = IN1[25]&IN2[29];
  assign P55[25] = IN1[25]&IN2[30];
  assign P56[25] = IN1[25]&IN2[31];
  assign P57[25] = IN1[25]&IN2[32];
  assign P58[25] = IN1[25]&IN2[33];
  assign P59[25] = IN1[25]&IN2[34];
  assign P60[25] = IN1[25]&IN2[35];
  assign P61[25] = IN1[25]&IN2[36];
  assign P62[24] = IN1[25]&IN2[37];
  assign P63[23] = IN1[25]&IN2[38];
  assign P64[22] = IN1[25]&IN2[39];
  assign P65[21] = IN1[25]&IN2[40];
  assign P66[20] = IN1[25]&IN2[41];
  assign P67[19] = IN1[25]&IN2[42];
  assign P68[18] = IN1[25]&IN2[43];
  assign P69[17] = IN1[25]&IN2[44];
  assign P70[16] = IN1[25]&IN2[45];
  assign P71[15] = IN1[25]&IN2[46];
  assign P72[14] = IN1[25]&IN2[47];
  assign P73[13] = IN1[25]&IN2[48];
  assign P74[12] = IN1[25]&IN2[49];
  assign P75[11] = IN1[25]&IN2[50];
  assign P76[10] = IN1[25]&IN2[51];
  assign P77[9] = IN1[25]&IN2[52];
  assign P78[8] = IN1[25]&IN2[53];
  assign P79[7] = IN1[25]&IN2[54];
  assign P80[6] = IN1[25]&IN2[55];
  assign P81[5] = IN1[25]&IN2[56];
  assign P82[4] = IN1[25]&IN2[57];
  assign P83[3] = IN1[25]&IN2[58];
  assign P84[2] = IN1[25]&IN2[59];
  assign P85[1] = IN1[25]&IN2[60];
  assign P86[0] = IN1[25]&IN2[61];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[26] = IN1[26]&IN2[3];
  assign P30[26] = IN1[26]&IN2[4];
  assign P31[26] = IN1[26]&IN2[5];
  assign P32[26] = IN1[26]&IN2[6];
  assign P33[26] = IN1[26]&IN2[7];
  assign P34[26] = IN1[26]&IN2[8];
  assign P35[26] = IN1[26]&IN2[9];
  assign P36[26] = IN1[26]&IN2[10];
  assign P37[26] = IN1[26]&IN2[11];
  assign P38[26] = IN1[26]&IN2[12];
  assign P39[26] = IN1[26]&IN2[13];
  assign P40[26] = IN1[26]&IN2[14];
  assign P41[26] = IN1[26]&IN2[15];
  assign P42[26] = IN1[26]&IN2[16];
  assign P43[26] = IN1[26]&IN2[17];
  assign P44[26] = IN1[26]&IN2[18];
  assign P45[26] = IN1[26]&IN2[19];
  assign P46[26] = IN1[26]&IN2[20];
  assign P47[26] = IN1[26]&IN2[21];
  assign P48[26] = IN1[26]&IN2[22];
  assign P49[26] = IN1[26]&IN2[23];
  assign P50[26] = IN1[26]&IN2[24];
  assign P51[26] = IN1[26]&IN2[25];
  assign P52[26] = IN1[26]&IN2[26];
  assign P53[26] = IN1[26]&IN2[27];
  assign P54[26] = IN1[26]&IN2[28];
  assign P55[26] = IN1[26]&IN2[29];
  assign P56[26] = IN1[26]&IN2[30];
  assign P57[26] = IN1[26]&IN2[31];
  assign P58[26] = IN1[26]&IN2[32];
  assign P59[26] = IN1[26]&IN2[33];
  assign P60[26] = IN1[26]&IN2[34];
  assign P61[26] = IN1[26]&IN2[35];
  assign P62[25] = IN1[26]&IN2[36];
  assign P63[24] = IN1[26]&IN2[37];
  assign P64[23] = IN1[26]&IN2[38];
  assign P65[22] = IN1[26]&IN2[39];
  assign P66[21] = IN1[26]&IN2[40];
  assign P67[20] = IN1[26]&IN2[41];
  assign P68[19] = IN1[26]&IN2[42];
  assign P69[18] = IN1[26]&IN2[43];
  assign P70[17] = IN1[26]&IN2[44];
  assign P71[16] = IN1[26]&IN2[45];
  assign P72[15] = IN1[26]&IN2[46];
  assign P73[14] = IN1[26]&IN2[47];
  assign P74[13] = IN1[26]&IN2[48];
  assign P75[12] = IN1[26]&IN2[49];
  assign P76[11] = IN1[26]&IN2[50];
  assign P77[10] = IN1[26]&IN2[51];
  assign P78[9] = IN1[26]&IN2[52];
  assign P79[8] = IN1[26]&IN2[53];
  assign P80[7] = IN1[26]&IN2[54];
  assign P81[6] = IN1[26]&IN2[55];
  assign P82[5] = IN1[26]&IN2[56];
  assign P83[4] = IN1[26]&IN2[57];
  assign P84[3] = IN1[26]&IN2[58];
  assign P85[2] = IN1[26]&IN2[59];
  assign P86[1] = IN1[26]&IN2[60];
  assign P87[0] = IN1[26]&IN2[61];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[27] = IN1[27]&IN2[2];
  assign P30[27] = IN1[27]&IN2[3];
  assign P31[27] = IN1[27]&IN2[4];
  assign P32[27] = IN1[27]&IN2[5];
  assign P33[27] = IN1[27]&IN2[6];
  assign P34[27] = IN1[27]&IN2[7];
  assign P35[27] = IN1[27]&IN2[8];
  assign P36[27] = IN1[27]&IN2[9];
  assign P37[27] = IN1[27]&IN2[10];
  assign P38[27] = IN1[27]&IN2[11];
  assign P39[27] = IN1[27]&IN2[12];
  assign P40[27] = IN1[27]&IN2[13];
  assign P41[27] = IN1[27]&IN2[14];
  assign P42[27] = IN1[27]&IN2[15];
  assign P43[27] = IN1[27]&IN2[16];
  assign P44[27] = IN1[27]&IN2[17];
  assign P45[27] = IN1[27]&IN2[18];
  assign P46[27] = IN1[27]&IN2[19];
  assign P47[27] = IN1[27]&IN2[20];
  assign P48[27] = IN1[27]&IN2[21];
  assign P49[27] = IN1[27]&IN2[22];
  assign P50[27] = IN1[27]&IN2[23];
  assign P51[27] = IN1[27]&IN2[24];
  assign P52[27] = IN1[27]&IN2[25];
  assign P53[27] = IN1[27]&IN2[26];
  assign P54[27] = IN1[27]&IN2[27];
  assign P55[27] = IN1[27]&IN2[28];
  assign P56[27] = IN1[27]&IN2[29];
  assign P57[27] = IN1[27]&IN2[30];
  assign P58[27] = IN1[27]&IN2[31];
  assign P59[27] = IN1[27]&IN2[32];
  assign P60[27] = IN1[27]&IN2[33];
  assign P61[27] = IN1[27]&IN2[34];
  assign P62[26] = IN1[27]&IN2[35];
  assign P63[25] = IN1[27]&IN2[36];
  assign P64[24] = IN1[27]&IN2[37];
  assign P65[23] = IN1[27]&IN2[38];
  assign P66[22] = IN1[27]&IN2[39];
  assign P67[21] = IN1[27]&IN2[40];
  assign P68[20] = IN1[27]&IN2[41];
  assign P69[19] = IN1[27]&IN2[42];
  assign P70[18] = IN1[27]&IN2[43];
  assign P71[17] = IN1[27]&IN2[44];
  assign P72[16] = IN1[27]&IN2[45];
  assign P73[15] = IN1[27]&IN2[46];
  assign P74[14] = IN1[27]&IN2[47];
  assign P75[13] = IN1[27]&IN2[48];
  assign P76[12] = IN1[27]&IN2[49];
  assign P77[11] = IN1[27]&IN2[50];
  assign P78[10] = IN1[27]&IN2[51];
  assign P79[9] = IN1[27]&IN2[52];
  assign P80[8] = IN1[27]&IN2[53];
  assign P81[7] = IN1[27]&IN2[54];
  assign P82[6] = IN1[27]&IN2[55];
  assign P83[5] = IN1[27]&IN2[56];
  assign P84[4] = IN1[27]&IN2[57];
  assign P85[3] = IN1[27]&IN2[58];
  assign P86[2] = IN1[27]&IN2[59];
  assign P87[1] = IN1[27]&IN2[60];
  assign P88[0] = IN1[27]&IN2[61];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[28] = IN1[28]&IN2[1];
  assign P30[28] = IN1[28]&IN2[2];
  assign P31[28] = IN1[28]&IN2[3];
  assign P32[28] = IN1[28]&IN2[4];
  assign P33[28] = IN1[28]&IN2[5];
  assign P34[28] = IN1[28]&IN2[6];
  assign P35[28] = IN1[28]&IN2[7];
  assign P36[28] = IN1[28]&IN2[8];
  assign P37[28] = IN1[28]&IN2[9];
  assign P38[28] = IN1[28]&IN2[10];
  assign P39[28] = IN1[28]&IN2[11];
  assign P40[28] = IN1[28]&IN2[12];
  assign P41[28] = IN1[28]&IN2[13];
  assign P42[28] = IN1[28]&IN2[14];
  assign P43[28] = IN1[28]&IN2[15];
  assign P44[28] = IN1[28]&IN2[16];
  assign P45[28] = IN1[28]&IN2[17];
  assign P46[28] = IN1[28]&IN2[18];
  assign P47[28] = IN1[28]&IN2[19];
  assign P48[28] = IN1[28]&IN2[20];
  assign P49[28] = IN1[28]&IN2[21];
  assign P50[28] = IN1[28]&IN2[22];
  assign P51[28] = IN1[28]&IN2[23];
  assign P52[28] = IN1[28]&IN2[24];
  assign P53[28] = IN1[28]&IN2[25];
  assign P54[28] = IN1[28]&IN2[26];
  assign P55[28] = IN1[28]&IN2[27];
  assign P56[28] = IN1[28]&IN2[28];
  assign P57[28] = IN1[28]&IN2[29];
  assign P58[28] = IN1[28]&IN2[30];
  assign P59[28] = IN1[28]&IN2[31];
  assign P60[28] = IN1[28]&IN2[32];
  assign P61[28] = IN1[28]&IN2[33];
  assign P62[27] = IN1[28]&IN2[34];
  assign P63[26] = IN1[28]&IN2[35];
  assign P64[25] = IN1[28]&IN2[36];
  assign P65[24] = IN1[28]&IN2[37];
  assign P66[23] = IN1[28]&IN2[38];
  assign P67[22] = IN1[28]&IN2[39];
  assign P68[21] = IN1[28]&IN2[40];
  assign P69[20] = IN1[28]&IN2[41];
  assign P70[19] = IN1[28]&IN2[42];
  assign P71[18] = IN1[28]&IN2[43];
  assign P72[17] = IN1[28]&IN2[44];
  assign P73[16] = IN1[28]&IN2[45];
  assign P74[15] = IN1[28]&IN2[46];
  assign P75[14] = IN1[28]&IN2[47];
  assign P76[13] = IN1[28]&IN2[48];
  assign P77[12] = IN1[28]&IN2[49];
  assign P78[11] = IN1[28]&IN2[50];
  assign P79[10] = IN1[28]&IN2[51];
  assign P80[9] = IN1[28]&IN2[52];
  assign P81[8] = IN1[28]&IN2[53];
  assign P82[7] = IN1[28]&IN2[54];
  assign P83[6] = IN1[28]&IN2[55];
  assign P84[5] = IN1[28]&IN2[56];
  assign P85[4] = IN1[28]&IN2[57];
  assign P86[3] = IN1[28]&IN2[58];
  assign P87[2] = IN1[28]&IN2[59];
  assign P88[1] = IN1[28]&IN2[60];
  assign P89[0] = IN1[28]&IN2[61];
  assign P29[29] = IN1[29]&IN2[0];
  assign P30[29] = IN1[29]&IN2[1];
  assign P31[29] = IN1[29]&IN2[2];
  assign P32[29] = IN1[29]&IN2[3];
  assign P33[29] = IN1[29]&IN2[4];
  assign P34[29] = IN1[29]&IN2[5];
  assign P35[29] = IN1[29]&IN2[6];
  assign P36[29] = IN1[29]&IN2[7];
  assign P37[29] = IN1[29]&IN2[8];
  assign P38[29] = IN1[29]&IN2[9];
  assign P39[29] = IN1[29]&IN2[10];
  assign P40[29] = IN1[29]&IN2[11];
  assign P41[29] = IN1[29]&IN2[12];
  assign P42[29] = IN1[29]&IN2[13];
  assign P43[29] = IN1[29]&IN2[14];
  assign P44[29] = IN1[29]&IN2[15];
  assign P45[29] = IN1[29]&IN2[16];
  assign P46[29] = IN1[29]&IN2[17];
  assign P47[29] = IN1[29]&IN2[18];
  assign P48[29] = IN1[29]&IN2[19];
  assign P49[29] = IN1[29]&IN2[20];
  assign P50[29] = IN1[29]&IN2[21];
  assign P51[29] = IN1[29]&IN2[22];
  assign P52[29] = IN1[29]&IN2[23];
  assign P53[29] = IN1[29]&IN2[24];
  assign P54[29] = IN1[29]&IN2[25];
  assign P55[29] = IN1[29]&IN2[26];
  assign P56[29] = IN1[29]&IN2[27];
  assign P57[29] = IN1[29]&IN2[28];
  assign P58[29] = IN1[29]&IN2[29];
  assign P59[29] = IN1[29]&IN2[30];
  assign P60[29] = IN1[29]&IN2[31];
  assign P61[29] = IN1[29]&IN2[32];
  assign P62[28] = IN1[29]&IN2[33];
  assign P63[27] = IN1[29]&IN2[34];
  assign P64[26] = IN1[29]&IN2[35];
  assign P65[25] = IN1[29]&IN2[36];
  assign P66[24] = IN1[29]&IN2[37];
  assign P67[23] = IN1[29]&IN2[38];
  assign P68[22] = IN1[29]&IN2[39];
  assign P69[21] = IN1[29]&IN2[40];
  assign P70[20] = IN1[29]&IN2[41];
  assign P71[19] = IN1[29]&IN2[42];
  assign P72[18] = IN1[29]&IN2[43];
  assign P73[17] = IN1[29]&IN2[44];
  assign P74[16] = IN1[29]&IN2[45];
  assign P75[15] = IN1[29]&IN2[46];
  assign P76[14] = IN1[29]&IN2[47];
  assign P77[13] = IN1[29]&IN2[48];
  assign P78[12] = IN1[29]&IN2[49];
  assign P79[11] = IN1[29]&IN2[50];
  assign P80[10] = IN1[29]&IN2[51];
  assign P81[9] = IN1[29]&IN2[52];
  assign P82[8] = IN1[29]&IN2[53];
  assign P83[7] = IN1[29]&IN2[54];
  assign P84[6] = IN1[29]&IN2[55];
  assign P85[5] = IN1[29]&IN2[56];
  assign P86[4] = IN1[29]&IN2[57];
  assign P87[3] = IN1[29]&IN2[58];
  assign P88[2] = IN1[29]&IN2[59];
  assign P89[1] = IN1[29]&IN2[60];
  assign P90[0] = IN1[29]&IN2[61];
  assign P30[30] = IN1[30]&IN2[0];
  assign P31[30] = IN1[30]&IN2[1];
  assign P32[30] = IN1[30]&IN2[2];
  assign P33[30] = IN1[30]&IN2[3];
  assign P34[30] = IN1[30]&IN2[4];
  assign P35[30] = IN1[30]&IN2[5];
  assign P36[30] = IN1[30]&IN2[6];
  assign P37[30] = IN1[30]&IN2[7];
  assign P38[30] = IN1[30]&IN2[8];
  assign P39[30] = IN1[30]&IN2[9];
  assign P40[30] = IN1[30]&IN2[10];
  assign P41[30] = IN1[30]&IN2[11];
  assign P42[30] = IN1[30]&IN2[12];
  assign P43[30] = IN1[30]&IN2[13];
  assign P44[30] = IN1[30]&IN2[14];
  assign P45[30] = IN1[30]&IN2[15];
  assign P46[30] = IN1[30]&IN2[16];
  assign P47[30] = IN1[30]&IN2[17];
  assign P48[30] = IN1[30]&IN2[18];
  assign P49[30] = IN1[30]&IN2[19];
  assign P50[30] = IN1[30]&IN2[20];
  assign P51[30] = IN1[30]&IN2[21];
  assign P52[30] = IN1[30]&IN2[22];
  assign P53[30] = IN1[30]&IN2[23];
  assign P54[30] = IN1[30]&IN2[24];
  assign P55[30] = IN1[30]&IN2[25];
  assign P56[30] = IN1[30]&IN2[26];
  assign P57[30] = IN1[30]&IN2[27];
  assign P58[30] = IN1[30]&IN2[28];
  assign P59[30] = IN1[30]&IN2[29];
  assign P60[30] = IN1[30]&IN2[30];
  assign P61[30] = IN1[30]&IN2[31];
  assign P62[29] = IN1[30]&IN2[32];
  assign P63[28] = IN1[30]&IN2[33];
  assign P64[27] = IN1[30]&IN2[34];
  assign P65[26] = IN1[30]&IN2[35];
  assign P66[25] = IN1[30]&IN2[36];
  assign P67[24] = IN1[30]&IN2[37];
  assign P68[23] = IN1[30]&IN2[38];
  assign P69[22] = IN1[30]&IN2[39];
  assign P70[21] = IN1[30]&IN2[40];
  assign P71[20] = IN1[30]&IN2[41];
  assign P72[19] = IN1[30]&IN2[42];
  assign P73[18] = IN1[30]&IN2[43];
  assign P74[17] = IN1[30]&IN2[44];
  assign P75[16] = IN1[30]&IN2[45];
  assign P76[15] = IN1[30]&IN2[46];
  assign P77[14] = IN1[30]&IN2[47];
  assign P78[13] = IN1[30]&IN2[48];
  assign P79[12] = IN1[30]&IN2[49];
  assign P80[11] = IN1[30]&IN2[50];
  assign P81[10] = IN1[30]&IN2[51];
  assign P82[9] = IN1[30]&IN2[52];
  assign P83[8] = IN1[30]&IN2[53];
  assign P84[7] = IN1[30]&IN2[54];
  assign P85[6] = IN1[30]&IN2[55];
  assign P86[5] = IN1[30]&IN2[56];
  assign P87[4] = IN1[30]&IN2[57];
  assign P88[3] = IN1[30]&IN2[58];
  assign P89[2] = IN1[30]&IN2[59];
  assign P90[1] = IN1[30]&IN2[60];
  assign P91[0] = IN1[30]&IN2[61];
  assign P31[31] = IN1[31]&IN2[0];
  assign P32[31] = IN1[31]&IN2[1];
  assign P33[31] = IN1[31]&IN2[2];
  assign P34[31] = IN1[31]&IN2[3];
  assign P35[31] = IN1[31]&IN2[4];
  assign P36[31] = IN1[31]&IN2[5];
  assign P37[31] = IN1[31]&IN2[6];
  assign P38[31] = IN1[31]&IN2[7];
  assign P39[31] = IN1[31]&IN2[8];
  assign P40[31] = IN1[31]&IN2[9];
  assign P41[31] = IN1[31]&IN2[10];
  assign P42[31] = IN1[31]&IN2[11];
  assign P43[31] = IN1[31]&IN2[12];
  assign P44[31] = IN1[31]&IN2[13];
  assign P45[31] = IN1[31]&IN2[14];
  assign P46[31] = IN1[31]&IN2[15];
  assign P47[31] = IN1[31]&IN2[16];
  assign P48[31] = IN1[31]&IN2[17];
  assign P49[31] = IN1[31]&IN2[18];
  assign P50[31] = IN1[31]&IN2[19];
  assign P51[31] = IN1[31]&IN2[20];
  assign P52[31] = IN1[31]&IN2[21];
  assign P53[31] = IN1[31]&IN2[22];
  assign P54[31] = IN1[31]&IN2[23];
  assign P55[31] = IN1[31]&IN2[24];
  assign P56[31] = IN1[31]&IN2[25];
  assign P57[31] = IN1[31]&IN2[26];
  assign P58[31] = IN1[31]&IN2[27];
  assign P59[31] = IN1[31]&IN2[28];
  assign P60[31] = IN1[31]&IN2[29];
  assign P61[31] = IN1[31]&IN2[30];
  assign P62[30] = IN1[31]&IN2[31];
  assign P63[29] = IN1[31]&IN2[32];
  assign P64[28] = IN1[31]&IN2[33];
  assign P65[27] = IN1[31]&IN2[34];
  assign P66[26] = IN1[31]&IN2[35];
  assign P67[25] = IN1[31]&IN2[36];
  assign P68[24] = IN1[31]&IN2[37];
  assign P69[23] = IN1[31]&IN2[38];
  assign P70[22] = IN1[31]&IN2[39];
  assign P71[21] = IN1[31]&IN2[40];
  assign P72[20] = IN1[31]&IN2[41];
  assign P73[19] = IN1[31]&IN2[42];
  assign P74[18] = IN1[31]&IN2[43];
  assign P75[17] = IN1[31]&IN2[44];
  assign P76[16] = IN1[31]&IN2[45];
  assign P77[15] = IN1[31]&IN2[46];
  assign P78[14] = IN1[31]&IN2[47];
  assign P79[13] = IN1[31]&IN2[48];
  assign P80[12] = IN1[31]&IN2[49];
  assign P81[11] = IN1[31]&IN2[50];
  assign P82[10] = IN1[31]&IN2[51];
  assign P83[9] = IN1[31]&IN2[52];
  assign P84[8] = IN1[31]&IN2[53];
  assign P85[7] = IN1[31]&IN2[54];
  assign P86[6] = IN1[31]&IN2[55];
  assign P87[5] = IN1[31]&IN2[56];
  assign P88[4] = IN1[31]&IN2[57];
  assign P89[3] = IN1[31]&IN2[58];
  assign P90[2] = IN1[31]&IN2[59];
  assign P91[1] = IN1[31]&IN2[60];
  assign P92[0] = IN1[31]&IN2[61];
  assign P32[32] = IN1[32]&IN2[0];
  assign P33[32] = IN1[32]&IN2[1];
  assign P34[32] = IN1[32]&IN2[2];
  assign P35[32] = IN1[32]&IN2[3];
  assign P36[32] = IN1[32]&IN2[4];
  assign P37[32] = IN1[32]&IN2[5];
  assign P38[32] = IN1[32]&IN2[6];
  assign P39[32] = IN1[32]&IN2[7];
  assign P40[32] = IN1[32]&IN2[8];
  assign P41[32] = IN1[32]&IN2[9];
  assign P42[32] = IN1[32]&IN2[10];
  assign P43[32] = IN1[32]&IN2[11];
  assign P44[32] = IN1[32]&IN2[12];
  assign P45[32] = IN1[32]&IN2[13];
  assign P46[32] = IN1[32]&IN2[14];
  assign P47[32] = IN1[32]&IN2[15];
  assign P48[32] = IN1[32]&IN2[16];
  assign P49[32] = IN1[32]&IN2[17];
  assign P50[32] = IN1[32]&IN2[18];
  assign P51[32] = IN1[32]&IN2[19];
  assign P52[32] = IN1[32]&IN2[20];
  assign P53[32] = IN1[32]&IN2[21];
  assign P54[32] = IN1[32]&IN2[22];
  assign P55[32] = IN1[32]&IN2[23];
  assign P56[32] = IN1[32]&IN2[24];
  assign P57[32] = IN1[32]&IN2[25];
  assign P58[32] = IN1[32]&IN2[26];
  assign P59[32] = IN1[32]&IN2[27];
  assign P60[32] = IN1[32]&IN2[28];
  assign P61[32] = IN1[32]&IN2[29];
  assign P62[31] = IN1[32]&IN2[30];
  assign P63[30] = IN1[32]&IN2[31];
  assign P64[29] = IN1[32]&IN2[32];
  assign P65[28] = IN1[32]&IN2[33];
  assign P66[27] = IN1[32]&IN2[34];
  assign P67[26] = IN1[32]&IN2[35];
  assign P68[25] = IN1[32]&IN2[36];
  assign P69[24] = IN1[32]&IN2[37];
  assign P70[23] = IN1[32]&IN2[38];
  assign P71[22] = IN1[32]&IN2[39];
  assign P72[21] = IN1[32]&IN2[40];
  assign P73[20] = IN1[32]&IN2[41];
  assign P74[19] = IN1[32]&IN2[42];
  assign P75[18] = IN1[32]&IN2[43];
  assign P76[17] = IN1[32]&IN2[44];
  assign P77[16] = IN1[32]&IN2[45];
  assign P78[15] = IN1[32]&IN2[46];
  assign P79[14] = IN1[32]&IN2[47];
  assign P80[13] = IN1[32]&IN2[48];
  assign P81[12] = IN1[32]&IN2[49];
  assign P82[11] = IN1[32]&IN2[50];
  assign P83[10] = IN1[32]&IN2[51];
  assign P84[9] = IN1[32]&IN2[52];
  assign P85[8] = IN1[32]&IN2[53];
  assign P86[7] = IN1[32]&IN2[54];
  assign P87[6] = IN1[32]&IN2[55];
  assign P88[5] = IN1[32]&IN2[56];
  assign P89[4] = IN1[32]&IN2[57];
  assign P90[3] = IN1[32]&IN2[58];
  assign P91[2] = IN1[32]&IN2[59];
  assign P92[1] = IN1[32]&IN2[60];
  assign P93[0] = IN1[32]&IN2[61];
  assign P33[33] = IN1[33]&IN2[0];
  assign P34[33] = IN1[33]&IN2[1];
  assign P35[33] = IN1[33]&IN2[2];
  assign P36[33] = IN1[33]&IN2[3];
  assign P37[33] = IN1[33]&IN2[4];
  assign P38[33] = IN1[33]&IN2[5];
  assign P39[33] = IN1[33]&IN2[6];
  assign P40[33] = IN1[33]&IN2[7];
  assign P41[33] = IN1[33]&IN2[8];
  assign P42[33] = IN1[33]&IN2[9];
  assign P43[33] = IN1[33]&IN2[10];
  assign P44[33] = IN1[33]&IN2[11];
  assign P45[33] = IN1[33]&IN2[12];
  assign P46[33] = IN1[33]&IN2[13];
  assign P47[33] = IN1[33]&IN2[14];
  assign P48[33] = IN1[33]&IN2[15];
  assign P49[33] = IN1[33]&IN2[16];
  assign P50[33] = IN1[33]&IN2[17];
  assign P51[33] = IN1[33]&IN2[18];
  assign P52[33] = IN1[33]&IN2[19];
  assign P53[33] = IN1[33]&IN2[20];
  assign P54[33] = IN1[33]&IN2[21];
  assign P55[33] = IN1[33]&IN2[22];
  assign P56[33] = IN1[33]&IN2[23];
  assign P57[33] = IN1[33]&IN2[24];
  assign P58[33] = IN1[33]&IN2[25];
  assign P59[33] = IN1[33]&IN2[26];
  assign P60[33] = IN1[33]&IN2[27];
  assign P61[33] = IN1[33]&IN2[28];
  assign P62[32] = IN1[33]&IN2[29];
  assign P63[31] = IN1[33]&IN2[30];
  assign P64[30] = IN1[33]&IN2[31];
  assign P65[29] = IN1[33]&IN2[32];
  assign P66[28] = IN1[33]&IN2[33];
  assign P67[27] = IN1[33]&IN2[34];
  assign P68[26] = IN1[33]&IN2[35];
  assign P69[25] = IN1[33]&IN2[36];
  assign P70[24] = IN1[33]&IN2[37];
  assign P71[23] = IN1[33]&IN2[38];
  assign P72[22] = IN1[33]&IN2[39];
  assign P73[21] = IN1[33]&IN2[40];
  assign P74[20] = IN1[33]&IN2[41];
  assign P75[19] = IN1[33]&IN2[42];
  assign P76[18] = IN1[33]&IN2[43];
  assign P77[17] = IN1[33]&IN2[44];
  assign P78[16] = IN1[33]&IN2[45];
  assign P79[15] = IN1[33]&IN2[46];
  assign P80[14] = IN1[33]&IN2[47];
  assign P81[13] = IN1[33]&IN2[48];
  assign P82[12] = IN1[33]&IN2[49];
  assign P83[11] = IN1[33]&IN2[50];
  assign P84[10] = IN1[33]&IN2[51];
  assign P85[9] = IN1[33]&IN2[52];
  assign P86[8] = IN1[33]&IN2[53];
  assign P87[7] = IN1[33]&IN2[54];
  assign P88[6] = IN1[33]&IN2[55];
  assign P89[5] = IN1[33]&IN2[56];
  assign P90[4] = IN1[33]&IN2[57];
  assign P91[3] = IN1[33]&IN2[58];
  assign P92[2] = IN1[33]&IN2[59];
  assign P93[1] = IN1[33]&IN2[60];
  assign P94[0] = IN1[33]&IN2[61];
  assign P34[34] = IN1[34]&IN2[0];
  assign P35[34] = IN1[34]&IN2[1];
  assign P36[34] = IN1[34]&IN2[2];
  assign P37[34] = IN1[34]&IN2[3];
  assign P38[34] = IN1[34]&IN2[4];
  assign P39[34] = IN1[34]&IN2[5];
  assign P40[34] = IN1[34]&IN2[6];
  assign P41[34] = IN1[34]&IN2[7];
  assign P42[34] = IN1[34]&IN2[8];
  assign P43[34] = IN1[34]&IN2[9];
  assign P44[34] = IN1[34]&IN2[10];
  assign P45[34] = IN1[34]&IN2[11];
  assign P46[34] = IN1[34]&IN2[12];
  assign P47[34] = IN1[34]&IN2[13];
  assign P48[34] = IN1[34]&IN2[14];
  assign P49[34] = IN1[34]&IN2[15];
  assign P50[34] = IN1[34]&IN2[16];
  assign P51[34] = IN1[34]&IN2[17];
  assign P52[34] = IN1[34]&IN2[18];
  assign P53[34] = IN1[34]&IN2[19];
  assign P54[34] = IN1[34]&IN2[20];
  assign P55[34] = IN1[34]&IN2[21];
  assign P56[34] = IN1[34]&IN2[22];
  assign P57[34] = IN1[34]&IN2[23];
  assign P58[34] = IN1[34]&IN2[24];
  assign P59[34] = IN1[34]&IN2[25];
  assign P60[34] = IN1[34]&IN2[26];
  assign P61[34] = IN1[34]&IN2[27];
  assign P62[33] = IN1[34]&IN2[28];
  assign P63[32] = IN1[34]&IN2[29];
  assign P64[31] = IN1[34]&IN2[30];
  assign P65[30] = IN1[34]&IN2[31];
  assign P66[29] = IN1[34]&IN2[32];
  assign P67[28] = IN1[34]&IN2[33];
  assign P68[27] = IN1[34]&IN2[34];
  assign P69[26] = IN1[34]&IN2[35];
  assign P70[25] = IN1[34]&IN2[36];
  assign P71[24] = IN1[34]&IN2[37];
  assign P72[23] = IN1[34]&IN2[38];
  assign P73[22] = IN1[34]&IN2[39];
  assign P74[21] = IN1[34]&IN2[40];
  assign P75[20] = IN1[34]&IN2[41];
  assign P76[19] = IN1[34]&IN2[42];
  assign P77[18] = IN1[34]&IN2[43];
  assign P78[17] = IN1[34]&IN2[44];
  assign P79[16] = IN1[34]&IN2[45];
  assign P80[15] = IN1[34]&IN2[46];
  assign P81[14] = IN1[34]&IN2[47];
  assign P82[13] = IN1[34]&IN2[48];
  assign P83[12] = IN1[34]&IN2[49];
  assign P84[11] = IN1[34]&IN2[50];
  assign P85[10] = IN1[34]&IN2[51];
  assign P86[9] = IN1[34]&IN2[52];
  assign P87[8] = IN1[34]&IN2[53];
  assign P88[7] = IN1[34]&IN2[54];
  assign P89[6] = IN1[34]&IN2[55];
  assign P90[5] = IN1[34]&IN2[56];
  assign P91[4] = IN1[34]&IN2[57];
  assign P92[3] = IN1[34]&IN2[58];
  assign P93[2] = IN1[34]&IN2[59];
  assign P94[1] = IN1[34]&IN2[60];
  assign P95[0] = IN1[34]&IN2[61];
  assign P35[35] = IN1[35]&IN2[0];
  assign P36[35] = IN1[35]&IN2[1];
  assign P37[35] = IN1[35]&IN2[2];
  assign P38[35] = IN1[35]&IN2[3];
  assign P39[35] = IN1[35]&IN2[4];
  assign P40[35] = IN1[35]&IN2[5];
  assign P41[35] = IN1[35]&IN2[6];
  assign P42[35] = IN1[35]&IN2[7];
  assign P43[35] = IN1[35]&IN2[8];
  assign P44[35] = IN1[35]&IN2[9];
  assign P45[35] = IN1[35]&IN2[10];
  assign P46[35] = IN1[35]&IN2[11];
  assign P47[35] = IN1[35]&IN2[12];
  assign P48[35] = IN1[35]&IN2[13];
  assign P49[35] = IN1[35]&IN2[14];
  assign P50[35] = IN1[35]&IN2[15];
  assign P51[35] = IN1[35]&IN2[16];
  assign P52[35] = IN1[35]&IN2[17];
  assign P53[35] = IN1[35]&IN2[18];
  assign P54[35] = IN1[35]&IN2[19];
  assign P55[35] = IN1[35]&IN2[20];
  assign P56[35] = IN1[35]&IN2[21];
  assign P57[35] = IN1[35]&IN2[22];
  assign P58[35] = IN1[35]&IN2[23];
  assign P59[35] = IN1[35]&IN2[24];
  assign P60[35] = IN1[35]&IN2[25];
  assign P61[35] = IN1[35]&IN2[26];
  assign P62[34] = IN1[35]&IN2[27];
  assign P63[33] = IN1[35]&IN2[28];
  assign P64[32] = IN1[35]&IN2[29];
  assign P65[31] = IN1[35]&IN2[30];
  assign P66[30] = IN1[35]&IN2[31];
  assign P67[29] = IN1[35]&IN2[32];
  assign P68[28] = IN1[35]&IN2[33];
  assign P69[27] = IN1[35]&IN2[34];
  assign P70[26] = IN1[35]&IN2[35];
  assign P71[25] = IN1[35]&IN2[36];
  assign P72[24] = IN1[35]&IN2[37];
  assign P73[23] = IN1[35]&IN2[38];
  assign P74[22] = IN1[35]&IN2[39];
  assign P75[21] = IN1[35]&IN2[40];
  assign P76[20] = IN1[35]&IN2[41];
  assign P77[19] = IN1[35]&IN2[42];
  assign P78[18] = IN1[35]&IN2[43];
  assign P79[17] = IN1[35]&IN2[44];
  assign P80[16] = IN1[35]&IN2[45];
  assign P81[15] = IN1[35]&IN2[46];
  assign P82[14] = IN1[35]&IN2[47];
  assign P83[13] = IN1[35]&IN2[48];
  assign P84[12] = IN1[35]&IN2[49];
  assign P85[11] = IN1[35]&IN2[50];
  assign P86[10] = IN1[35]&IN2[51];
  assign P87[9] = IN1[35]&IN2[52];
  assign P88[8] = IN1[35]&IN2[53];
  assign P89[7] = IN1[35]&IN2[54];
  assign P90[6] = IN1[35]&IN2[55];
  assign P91[5] = IN1[35]&IN2[56];
  assign P92[4] = IN1[35]&IN2[57];
  assign P93[3] = IN1[35]&IN2[58];
  assign P94[2] = IN1[35]&IN2[59];
  assign P95[1] = IN1[35]&IN2[60];
  assign P96[0] = IN1[35]&IN2[61];
  assign P36[36] = IN1[36]&IN2[0];
  assign P37[36] = IN1[36]&IN2[1];
  assign P38[36] = IN1[36]&IN2[2];
  assign P39[36] = IN1[36]&IN2[3];
  assign P40[36] = IN1[36]&IN2[4];
  assign P41[36] = IN1[36]&IN2[5];
  assign P42[36] = IN1[36]&IN2[6];
  assign P43[36] = IN1[36]&IN2[7];
  assign P44[36] = IN1[36]&IN2[8];
  assign P45[36] = IN1[36]&IN2[9];
  assign P46[36] = IN1[36]&IN2[10];
  assign P47[36] = IN1[36]&IN2[11];
  assign P48[36] = IN1[36]&IN2[12];
  assign P49[36] = IN1[36]&IN2[13];
  assign P50[36] = IN1[36]&IN2[14];
  assign P51[36] = IN1[36]&IN2[15];
  assign P52[36] = IN1[36]&IN2[16];
  assign P53[36] = IN1[36]&IN2[17];
  assign P54[36] = IN1[36]&IN2[18];
  assign P55[36] = IN1[36]&IN2[19];
  assign P56[36] = IN1[36]&IN2[20];
  assign P57[36] = IN1[36]&IN2[21];
  assign P58[36] = IN1[36]&IN2[22];
  assign P59[36] = IN1[36]&IN2[23];
  assign P60[36] = IN1[36]&IN2[24];
  assign P61[36] = IN1[36]&IN2[25];
  assign P62[35] = IN1[36]&IN2[26];
  assign P63[34] = IN1[36]&IN2[27];
  assign P64[33] = IN1[36]&IN2[28];
  assign P65[32] = IN1[36]&IN2[29];
  assign P66[31] = IN1[36]&IN2[30];
  assign P67[30] = IN1[36]&IN2[31];
  assign P68[29] = IN1[36]&IN2[32];
  assign P69[28] = IN1[36]&IN2[33];
  assign P70[27] = IN1[36]&IN2[34];
  assign P71[26] = IN1[36]&IN2[35];
  assign P72[25] = IN1[36]&IN2[36];
  assign P73[24] = IN1[36]&IN2[37];
  assign P74[23] = IN1[36]&IN2[38];
  assign P75[22] = IN1[36]&IN2[39];
  assign P76[21] = IN1[36]&IN2[40];
  assign P77[20] = IN1[36]&IN2[41];
  assign P78[19] = IN1[36]&IN2[42];
  assign P79[18] = IN1[36]&IN2[43];
  assign P80[17] = IN1[36]&IN2[44];
  assign P81[16] = IN1[36]&IN2[45];
  assign P82[15] = IN1[36]&IN2[46];
  assign P83[14] = IN1[36]&IN2[47];
  assign P84[13] = IN1[36]&IN2[48];
  assign P85[12] = IN1[36]&IN2[49];
  assign P86[11] = IN1[36]&IN2[50];
  assign P87[10] = IN1[36]&IN2[51];
  assign P88[9] = IN1[36]&IN2[52];
  assign P89[8] = IN1[36]&IN2[53];
  assign P90[7] = IN1[36]&IN2[54];
  assign P91[6] = IN1[36]&IN2[55];
  assign P92[5] = IN1[36]&IN2[56];
  assign P93[4] = IN1[36]&IN2[57];
  assign P94[3] = IN1[36]&IN2[58];
  assign P95[2] = IN1[36]&IN2[59];
  assign P96[1] = IN1[36]&IN2[60];
  assign P97[0] = IN1[36]&IN2[61];
  assign P37[37] = IN1[37]&IN2[0];
  assign P38[37] = IN1[37]&IN2[1];
  assign P39[37] = IN1[37]&IN2[2];
  assign P40[37] = IN1[37]&IN2[3];
  assign P41[37] = IN1[37]&IN2[4];
  assign P42[37] = IN1[37]&IN2[5];
  assign P43[37] = IN1[37]&IN2[6];
  assign P44[37] = IN1[37]&IN2[7];
  assign P45[37] = IN1[37]&IN2[8];
  assign P46[37] = IN1[37]&IN2[9];
  assign P47[37] = IN1[37]&IN2[10];
  assign P48[37] = IN1[37]&IN2[11];
  assign P49[37] = IN1[37]&IN2[12];
  assign P50[37] = IN1[37]&IN2[13];
  assign P51[37] = IN1[37]&IN2[14];
  assign P52[37] = IN1[37]&IN2[15];
  assign P53[37] = IN1[37]&IN2[16];
  assign P54[37] = IN1[37]&IN2[17];
  assign P55[37] = IN1[37]&IN2[18];
  assign P56[37] = IN1[37]&IN2[19];
  assign P57[37] = IN1[37]&IN2[20];
  assign P58[37] = IN1[37]&IN2[21];
  assign P59[37] = IN1[37]&IN2[22];
  assign P60[37] = IN1[37]&IN2[23];
  assign P61[37] = IN1[37]&IN2[24];
  assign P62[36] = IN1[37]&IN2[25];
  assign P63[35] = IN1[37]&IN2[26];
  assign P64[34] = IN1[37]&IN2[27];
  assign P65[33] = IN1[37]&IN2[28];
  assign P66[32] = IN1[37]&IN2[29];
  assign P67[31] = IN1[37]&IN2[30];
  assign P68[30] = IN1[37]&IN2[31];
  assign P69[29] = IN1[37]&IN2[32];
  assign P70[28] = IN1[37]&IN2[33];
  assign P71[27] = IN1[37]&IN2[34];
  assign P72[26] = IN1[37]&IN2[35];
  assign P73[25] = IN1[37]&IN2[36];
  assign P74[24] = IN1[37]&IN2[37];
  assign P75[23] = IN1[37]&IN2[38];
  assign P76[22] = IN1[37]&IN2[39];
  assign P77[21] = IN1[37]&IN2[40];
  assign P78[20] = IN1[37]&IN2[41];
  assign P79[19] = IN1[37]&IN2[42];
  assign P80[18] = IN1[37]&IN2[43];
  assign P81[17] = IN1[37]&IN2[44];
  assign P82[16] = IN1[37]&IN2[45];
  assign P83[15] = IN1[37]&IN2[46];
  assign P84[14] = IN1[37]&IN2[47];
  assign P85[13] = IN1[37]&IN2[48];
  assign P86[12] = IN1[37]&IN2[49];
  assign P87[11] = IN1[37]&IN2[50];
  assign P88[10] = IN1[37]&IN2[51];
  assign P89[9] = IN1[37]&IN2[52];
  assign P90[8] = IN1[37]&IN2[53];
  assign P91[7] = IN1[37]&IN2[54];
  assign P92[6] = IN1[37]&IN2[55];
  assign P93[5] = IN1[37]&IN2[56];
  assign P94[4] = IN1[37]&IN2[57];
  assign P95[3] = IN1[37]&IN2[58];
  assign P96[2] = IN1[37]&IN2[59];
  assign P97[1] = IN1[37]&IN2[60];
  assign P98[0] = IN1[37]&IN2[61];
  assign P38[38] = IN1[38]&IN2[0];
  assign P39[38] = IN1[38]&IN2[1];
  assign P40[38] = IN1[38]&IN2[2];
  assign P41[38] = IN1[38]&IN2[3];
  assign P42[38] = IN1[38]&IN2[4];
  assign P43[38] = IN1[38]&IN2[5];
  assign P44[38] = IN1[38]&IN2[6];
  assign P45[38] = IN1[38]&IN2[7];
  assign P46[38] = IN1[38]&IN2[8];
  assign P47[38] = IN1[38]&IN2[9];
  assign P48[38] = IN1[38]&IN2[10];
  assign P49[38] = IN1[38]&IN2[11];
  assign P50[38] = IN1[38]&IN2[12];
  assign P51[38] = IN1[38]&IN2[13];
  assign P52[38] = IN1[38]&IN2[14];
  assign P53[38] = IN1[38]&IN2[15];
  assign P54[38] = IN1[38]&IN2[16];
  assign P55[38] = IN1[38]&IN2[17];
  assign P56[38] = IN1[38]&IN2[18];
  assign P57[38] = IN1[38]&IN2[19];
  assign P58[38] = IN1[38]&IN2[20];
  assign P59[38] = IN1[38]&IN2[21];
  assign P60[38] = IN1[38]&IN2[22];
  assign P61[38] = IN1[38]&IN2[23];
  assign P62[37] = IN1[38]&IN2[24];
  assign P63[36] = IN1[38]&IN2[25];
  assign P64[35] = IN1[38]&IN2[26];
  assign P65[34] = IN1[38]&IN2[27];
  assign P66[33] = IN1[38]&IN2[28];
  assign P67[32] = IN1[38]&IN2[29];
  assign P68[31] = IN1[38]&IN2[30];
  assign P69[30] = IN1[38]&IN2[31];
  assign P70[29] = IN1[38]&IN2[32];
  assign P71[28] = IN1[38]&IN2[33];
  assign P72[27] = IN1[38]&IN2[34];
  assign P73[26] = IN1[38]&IN2[35];
  assign P74[25] = IN1[38]&IN2[36];
  assign P75[24] = IN1[38]&IN2[37];
  assign P76[23] = IN1[38]&IN2[38];
  assign P77[22] = IN1[38]&IN2[39];
  assign P78[21] = IN1[38]&IN2[40];
  assign P79[20] = IN1[38]&IN2[41];
  assign P80[19] = IN1[38]&IN2[42];
  assign P81[18] = IN1[38]&IN2[43];
  assign P82[17] = IN1[38]&IN2[44];
  assign P83[16] = IN1[38]&IN2[45];
  assign P84[15] = IN1[38]&IN2[46];
  assign P85[14] = IN1[38]&IN2[47];
  assign P86[13] = IN1[38]&IN2[48];
  assign P87[12] = IN1[38]&IN2[49];
  assign P88[11] = IN1[38]&IN2[50];
  assign P89[10] = IN1[38]&IN2[51];
  assign P90[9] = IN1[38]&IN2[52];
  assign P91[8] = IN1[38]&IN2[53];
  assign P92[7] = IN1[38]&IN2[54];
  assign P93[6] = IN1[38]&IN2[55];
  assign P94[5] = IN1[38]&IN2[56];
  assign P95[4] = IN1[38]&IN2[57];
  assign P96[3] = IN1[38]&IN2[58];
  assign P97[2] = IN1[38]&IN2[59];
  assign P98[1] = IN1[38]&IN2[60];
  assign P99[0] = IN1[38]&IN2[61];
  assign P39[39] = IN1[39]&IN2[0];
  assign P40[39] = IN1[39]&IN2[1];
  assign P41[39] = IN1[39]&IN2[2];
  assign P42[39] = IN1[39]&IN2[3];
  assign P43[39] = IN1[39]&IN2[4];
  assign P44[39] = IN1[39]&IN2[5];
  assign P45[39] = IN1[39]&IN2[6];
  assign P46[39] = IN1[39]&IN2[7];
  assign P47[39] = IN1[39]&IN2[8];
  assign P48[39] = IN1[39]&IN2[9];
  assign P49[39] = IN1[39]&IN2[10];
  assign P50[39] = IN1[39]&IN2[11];
  assign P51[39] = IN1[39]&IN2[12];
  assign P52[39] = IN1[39]&IN2[13];
  assign P53[39] = IN1[39]&IN2[14];
  assign P54[39] = IN1[39]&IN2[15];
  assign P55[39] = IN1[39]&IN2[16];
  assign P56[39] = IN1[39]&IN2[17];
  assign P57[39] = IN1[39]&IN2[18];
  assign P58[39] = IN1[39]&IN2[19];
  assign P59[39] = IN1[39]&IN2[20];
  assign P60[39] = IN1[39]&IN2[21];
  assign P61[39] = IN1[39]&IN2[22];
  assign P62[38] = IN1[39]&IN2[23];
  assign P63[37] = IN1[39]&IN2[24];
  assign P64[36] = IN1[39]&IN2[25];
  assign P65[35] = IN1[39]&IN2[26];
  assign P66[34] = IN1[39]&IN2[27];
  assign P67[33] = IN1[39]&IN2[28];
  assign P68[32] = IN1[39]&IN2[29];
  assign P69[31] = IN1[39]&IN2[30];
  assign P70[30] = IN1[39]&IN2[31];
  assign P71[29] = IN1[39]&IN2[32];
  assign P72[28] = IN1[39]&IN2[33];
  assign P73[27] = IN1[39]&IN2[34];
  assign P74[26] = IN1[39]&IN2[35];
  assign P75[25] = IN1[39]&IN2[36];
  assign P76[24] = IN1[39]&IN2[37];
  assign P77[23] = IN1[39]&IN2[38];
  assign P78[22] = IN1[39]&IN2[39];
  assign P79[21] = IN1[39]&IN2[40];
  assign P80[20] = IN1[39]&IN2[41];
  assign P81[19] = IN1[39]&IN2[42];
  assign P82[18] = IN1[39]&IN2[43];
  assign P83[17] = IN1[39]&IN2[44];
  assign P84[16] = IN1[39]&IN2[45];
  assign P85[15] = IN1[39]&IN2[46];
  assign P86[14] = IN1[39]&IN2[47];
  assign P87[13] = IN1[39]&IN2[48];
  assign P88[12] = IN1[39]&IN2[49];
  assign P89[11] = IN1[39]&IN2[50];
  assign P90[10] = IN1[39]&IN2[51];
  assign P91[9] = IN1[39]&IN2[52];
  assign P92[8] = IN1[39]&IN2[53];
  assign P93[7] = IN1[39]&IN2[54];
  assign P94[6] = IN1[39]&IN2[55];
  assign P95[5] = IN1[39]&IN2[56];
  assign P96[4] = IN1[39]&IN2[57];
  assign P97[3] = IN1[39]&IN2[58];
  assign P98[2] = IN1[39]&IN2[59];
  assign P99[1] = IN1[39]&IN2[60];
  assign P100[0] = IN1[39]&IN2[61];
  assign P40[40] = IN1[40]&IN2[0];
  assign P41[40] = IN1[40]&IN2[1];
  assign P42[40] = IN1[40]&IN2[2];
  assign P43[40] = IN1[40]&IN2[3];
  assign P44[40] = IN1[40]&IN2[4];
  assign P45[40] = IN1[40]&IN2[5];
  assign P46[40] = IN1[40]&IN2[6];
  assign P47[40] = IN1[40]&IN2[7];
  assign P48[40] = IN1[40]&IN2[8];
  assign P49[40] = IN1[40]&IN2[9];
  assign P50[40] = IN1[40]&IN2[10];
  assign P51[40] = IN1[40]&IN2[11];
  assign P52[40] = IN1[40]&IN2[12];
  assign P53[40] = IN1[40]&IN2[13];
  assign P54[40] = IN1[40]&IN2[14];
  assign P55[40] = IN1[40]&IN2[15];
  assign P56[40] = IN1[40]&IN2[16];
  assign P57[40] = IN1[40]&IN2[17];
  assign P58[40] = IN1[40]&IN2[18];
  assign P59[40] = IN1[40]&IN2[19];
  assign P60[40] = IN1[40]&IN2[20];
  assign P61[40] = IN1[40]&IN2[21];
  assign P62[39] = IN1[40]&IN2[22];
  assign P63[38] = IN1[40]&IN2[23];
  assign P64[37] = IN1[40]&IN2[24];
  assign P65[36] = IN1[40]&IN2[25];
  assign P66[35] = IN1[40]&IN2[26];
  assign P67[34] = IN1[40]&IN2[27];
  assign P68[33] = IN1[40]&IN2[28];
  assign P69[32] = IN1[40]&IN2[29];
  assign P70[31] = IN1[40]&IN2[30];
  assign P71[30] = IN1[40]&IN2[31];
  assign P72[29] = IN1[40]&IN2[32];
  assign P73[28] = IN1[40]&IN2[33];
  assign P74[27] = IN1[40]&IN2[34];
  assign P75[26] = IN1[40]&IN2[35];
  assign P76[25] = IN1[40]&IN2[36];
  assign P77[24] = IN1[40]&IN2[37];
  assign P78[23] = IN1[40]&IN2[38];
  assign P79[22] = IN1[40]&IN2[39];
  assign P80[21] = IN1[40]&IN2[40];
  assign P81[20] = IN1[40]&IN2[41];
  assign P82[19] = IN1[40]&IN2[42];
  assign P83[18] = IN1[40]&IN2[43];
  assign P84[17] = IN1[40]&IN2[44];
  assign P85[16] = IN1[40]&IN2[45];
  assign P86[15] = IN1[40]&IN2[46];
  assign P87[14] = IN1[40]&IN2[47];
  assign P88[13] = IN1[40]&IN2[48];
  assign P89[12] = IN1[40]&IN2[49];
  assign P90[11] = IN1[40]&IN2[50];
  assign P91[10] = IN1[40]&IN2[51];
  assign P92[9] = IN1[40]&IN2[52];
  assign P93[8] = IN1[40]&IN2[53];
  assign P94[7] = IN1[40]&IN2[54];
  assign P95[6] = IN1[40]&IN2[55];
  assign P96[5] = IN1[40]&IN2[56];
  assign P97[4] = IN1[40]&IN2[57];
  assign P98[3] = IN1[40]&IN2[58];
  assign P99[2] = IN1[40]&IN2[59];
  assign P100[1] = IN1[40]&IN2[60];
  assign P101[0] = IN1[40]&IN2[61];
  assign P41[41] = IN1[41]&IN2[0];
  assign P42[41] = IN1[41]&IN2[1];
  assign P43[41] = IN1[41]&IN2[2];
  assign P44[41] = IN1[41]&IN2[3];
  assign P45[41] = IN1[41]&IN2[4];
  assign P46[41] = IN1[41]&IN2[5];
  assign P47[41] = IN1[41]&IN2[6];
  assign P48[41] = IN1[41]&IN2[7];
  assign P49[41] = IN1[41]&IN2[8];
  assign P50[41] = IN1[41]&IN2[9];
  assign P51[41] = IN1[41]&IN2[10];
  assign P52[41] = IN1[41]&IN2[11];
  assign P53[41] = IN1[41]&IN2[12];
  assign P54[41] = IN1[41]&IN2[13];
  assign P55[41] = IN1[41]&IN2[14];
  assign P56[41] = IN1[41]&IN2[15];
  assign P57[41] = IN1[41]&IN2[16];
  assign P58[41] = IN1[41]&IN2[17];
  assign P59[41] = IN1[41]&IN2[18];
  assign P60[41] = IN1[41]&IN2[19];
  assign P61[41] = IN1[41]&IN2[20];
  assign P62[40] = IN1[41]&IN2[21];
  assign P63[39] = IN1[41]&IN2[22];
  assign P64[38] = IN1[41]&IN2[23];
  assign P65[37] = IN1[41]&IN2[24];
  assign P66[36] = IN1[41]&IN2[25];
  assign P67[35] = IN1[41]&IN2[26];
  assign P68[34] = IN1[41]&IN2[27];
  assign P69[33] = IN1[41]&IN2[28];
  assign P70[32] = IN1[41]&IN2[29];
  assign P71[31] = IN1[41]&IN2[30];
  assign P72[30] = IN1[41]&IN2[31];
  assign P73[29] = IN1[41]&IN2[32];
  assign P74[28] = IN1[41]&IN2[33];
  assign P75[27] = IN1[41]&IN2[34];
  assign P76[26] = IN1[41]&IN2[35];
  assign P77[25] = IN1[41]&IN2[36];
  assign P78[24] = IN1[41]&IN2[37];
  assign P79[23] = IN1[41]&IN2[38];
  assign P80[22] = IN1[41]&IN2[39];
  assign P81[21] = IN1[41]&IN2[40];
  assign P82[20] = IN1[41]&IN2[41];
  assign P83[19] = IN1[41]&IN2[42];
  assign P84[18] = IN1[41]&IN2[43];
  assign P85[17] = IN1[41]&IN2[44];
  assign P86[16] = IN1[41]&IN2[45];
  assign P87[15] = IN1[41]&IN2[46];
  assign P88[14] = IN1[41]&IN2[47];
  assign P89[13] = IN1[41]&IN2[48];
  assign P90[12] = IN1[41]&IN2[49];
  assign P91[11] = IN1[41]&IN2[50];
  assign P92[10] = IN1[41]&IN2[51];
  assign P93[9] = IN1[41]&IN2[52];
  assign P94[8] = IN1[41]&IN2[53];
  assign P95[7] = IN1[41]&IN2[54];
  assign P96[6] = IN1[41]&IN2[55];
  assign P97[5] = IN1[41]&IN2[56];
  assign P98[4] = IN1[41]&IN2[57];
  assign P99[3] = IN1[41]&IN2[58];
  assign P100[2] = IN1[41]&IN2[59];
  assign P101[1] = IN1[41]&IN2[60];
  assign P102[0] = IN1[41]&IN2[61];
  assign P42[42] = IN1[42]&IN2[0];
  assign P43[42] = IN1[42]&IN2[1];
  assign P44[42] = IN1[42]&IN2[2];
  assign P45[42] = IN1[42]&IN2[3];
  assign P46[42] = IN1[42]&IN2[4];
  assign P47[42] = IN1[42]&IN2[5];
  assign P48[42] = IN1[42]&IN2[6];
  assign P49[42] = IN1[42]&IN2[7];
  assign P50[42] = IN1[42]&IN2[8];
  assign P51[42] = IN1[42]&IN2[9];
  assign P52[42] = IN1[42]&IN2[10];
  assign P53[42] = IN1[42]&IN2[11];
  assign P54[42] = IN1[42]&IN2[12];
  assign P55[42] = IN1[42]&IN2[13];
  assign P56[42] = IN1[42]&IN2[14];
  assign P57[42] = IN1[42]&IN2[15];
  assign P58[42] = IN1[42]&IN2[16];
  assign P59[42] = IN1[42]&IN2[17];
  assign P60[42] = IN1[42]&IN2[18];
  assign P61[42] = IN1[42]&IN2[19];
  assign P62[41] = IN1[42]&IN2[20];
  assign P63[40] = IN1[42]&IN2[21];
  assign P64[39] = IN1[42]&IN2[22];
  assign P65[38] = IN1[42]&IN2[23];
  assign P66[37] = IN1[42]&IN2[24];
  assign P67[36] = IN1[42]&IN2[25];
  assign P68[35] = IN1[42]&IN2[26];
  assign P69[34] = IN1[42]&IN2[27];
  assign P70[33] = IN1[42]&IN2[28];
  assign P71[32] = IN1[42]&IN2[29];
  assign P72[31] = IN1[42]&IN2[30];
  assign P73[30] = IN1[42]&IN2[31];
  assign P74[29] = IN1[42]&IN2[32];
  assign P75[28] = IN1[42]&IN2[33];
  assign P76[27] = IN1[42]&IN2[34];
  assign P77[26] = IN1[42]&IN2[35];
  assign P78[25] = IN1[42]&IN2[36];
  assign P79[24] = IN1[42]&IN2[37];
  assign P80[23] = IN1[42]&IN2[38];
  assign P81[22] = IN1[42]&IN2[39];
  assign P82[21] = IN1[42]&IN2[40];
  assign P83[20] = IN1[42]&IN2[41];
  assign P84[19] = IN1[42]&IN2[42];
  assign P85[18] = IN1[42]&IN2[43];
  assign P86[17] = IN1[42]&IN2[44];
  assign P87[16] = IN1[42]&IN2[45];
  assign P88[15] = IN1[42]&IN2[46];
  assign P89[14] = IN1[42]&IN2[47];
  assign P90[13] = IN1[42]&IN2[48];
  assign P91[12] = IN1[42]&IN2[49];
  assign P92[11] = IN1[42]&IN2[50];
  assign P93[10] = IN1[42]&IN2[51];
  assign P94[9] = IN1[42]&IN2[52];
  assign P95[8] = IN1[42]&IN2[53];
  assign P96[7] = IN1[42]&IN2[54];
  assign P97[6] = IN1[42]&IN2[55];
  assign P98[5] = IN1[42]&IN2[56];
  assign P99[4] = IN1[42]&IN2[57];
  assign P100[3] = IN1[42]&IN2[58];
  assign P101[2] = IN1[42]&IN2[59];
  assign P102[1] = IN1[42]&IN2[60];
  assign P103[0] = IN1[42]&IN2[61];
  assign P43[43] = IN1[43]&IN2[0];
  assign P44[43] = IN1[43]&IN2[1];
  assign P45[43] = IN1[43]&IN2[2];
  assign P46[43] = IN1[43]&IN2[3];
  assign P47[43] = IN1[43]&IN2[4];
  assign P48[43] = IN1[43]&IN2[5];
  assign P49[43] = IN1[43]&IN2[6];
  assign P50[43] = IN1[43]&IN2[7];
  assign P51[43] = IN1[43]&IN2[8];
  assign P52[43] = IN1[43]&IN2[9];
  assign P53[43] = IN1[43]&IN2[10];
  assign P54[43] = IN1[43]&IN2[11];
  assign P55[43] = IN1[43]&IN2[12];
  assign P56[43] = IN1[43]&IN2[13];
  assign P57[43] = IN1[43]&IN2[14];
  assign P58[43] = IN1[43]&IN2[15];
  assign P59[43] = IN1[43]&IN2[16];
  assign P60[43] = IN1[43]&IN2[17];
  assign P61[43] = IN1[43]&IN2[18];
  assign P62[42] = IN1[43]&IN2[19];
  assign P63[41] = IN1[43]&IN2[20];
  assign P64[40] = IN1[43]&IN2[21];
  assign P65[39] = IN1[43]&IN2[22];
  assign P66[38] = IN1[43]&IN2[23];
  assign P67[37] = IN1[43]&IN2[24];
  assign P68[36] = IN1[43]&IN2[25];
  assign P69[35] = IN1[43]&IN2[26];
  assign P70[34] = IN1[43]&IN2[27];
  assign P71[33] = IN1[43]&IN2[28];
  assign P72[32] = IN1[43]&IN2[29];
  assign P73[31] = IN1[43]&IN2[30];
  assign P74[30] = IN1[43]&IN2[31];
  assign P75[29] = IN1[43]&IN2[32];
  assign P76[28] = IN1[43]&IN2[33];
  assign P77[27] = IN1[43]&IN2[34];
  assign P78[26] = IN1[43]&IN2[35];
  assign P79[25] = IN1[43]&IN2[36];
  assign P80[24] = IN1[43]&IN2[37];
  assign P81[23] = IN1[43]&IN2[38];
  assign P82[22] = IN1[43]&IN2[39];
  assign P83[21] = IN1[43]&IN2[40];
  assign P84[20] = IN1[43]&IN2[41];
  assign P85[19] = IN1[43]&IN2[42];
  assign P86[18] = IN1[43]&IN2[43];
  assign P87[17] = IN1[43]&IN2[44];
  assign P88[16] = IN1[43]&IN2[45];
  assign P89[15] = IN1[43]&IN2[46];
  assign P90[14] = IN1[43]&IN2[47];
  assign P91[13] = IN1[43]&IN2[48];
  assign P92[12] = IN1[43]&IN2[49];
  assign P93[11] = IN1[43]&IN2[50];
  assign P94[10] = IN1[43]&IN2[51];
  assign P95[9] = IN1[43]&IN2[52];
  assign P96[8] = IN1[43]&IN2[53];
  assign P97[7] = IN1[43]&IN2[54];
  assign P98[6] = IN1[43]&IN2[55];
  assign P99[5] = IN1[43]&IN2[56];
  assign P100[4] = IN1[43]&IN2[57];
  assign P101[3] = IN1[43]&IN2[58];
  assign P102[2] = IN1[43]&IN2[59];
  assign P103[1] = IN1[43]&IN2[60];
  assign P104[0] = IN1[43]&IN2[61];
  assign P44[44] = IN1[44]&IN2[0];
  assign P45[44] = IN1[44]&IN2[1];
  assign P46[44] = IN1[44]&IN2[2];
  assign P47[44] = IN1[44]&IN2[3];
  assign P48[44] = IN1[44]&IN2[4];
  assign P49[44] = IN1[44]&IN2[5];
  assign P50[44] = IN1[44]&IN2[6];
  assign P51[44] = IN1[44]&IN2[7];
  assign P52[44] = IN1[44]&IN2[8];
  assign P53[44] = IN1[44]&IN2[9];
  assign P54[44] = IN1[44]&IN2[10];
  assign P55[44] = IN1[44]&IN2[11];
  assign P56[44] = IN1[44]&IN2[12];
  assign P57[44] = IN1[44]&IN2[13];
  assign P58[44] = IN1[44]&IN2[14];
  assign P59[44] = IN1[44]&IN2[15];
  assign P60[44] = IN1[44]&IN2[16];
  assign P61[44] = IN1[44]&IN2[17];
  assign P62[43] = IN1[44]&IN2[18];
  assign P63[42] = IN1[44]&IN2[19];
  assign P64[41] = IN1[44]&IN2[20];
  assign P65[40] = IN1[44]&IN2[21];
  assign P66[39] = IN1[44]&IN2[22];
  assign P67[38] = IN1[44]&IN2[23];
  assign P68[37] = IN1[44]&IN2[24];
  assign P69[36] = IN1[44]&IN2[25];
  assign P70[35] = IN1[44]&IN2[26];
  assign P71[34] = IN1[44]&IN2[27];
  assign P72[33] = IN1[44]&IN2[28];
  assign P73[32] = IN1[44]&IN2[29];
  assign P74[31] = IN1[44]&IN2[30];
  assign P75[30] = IN1[44]&IN2[31];
  assign P76[29] = IN1[44]&IN2[32];
  assign P77[28] = IN1[44]&IN2[33];
  assign P78[27] = IN1[44]&IN2[34];
  assign P79[26] = IN1[44]&IN2[35];
  assign P80[25] = IN1[44]&IN2[36];
  assign P81[24] = IN1[44]&IN2[37];
  assign P82[23] = IN1[44]&IN2[38];
  assign P83[22] = IN1[44]&IN2[39];
  assign P84[21] = IN1[44]&IN2[40];
  assign P85[20] = IN1[44]&IN2[41];
  assign P86[19] = IN1[44]&IN2[42];
  assign P87[18] = IN1[44]&IN2[43];
  assign P88[17] = IN1[44]&IN2[44];
  assign P89[16] = IN1[44]&IN2[45];
  assign P90[15] = IN1[44]&IN2[46];
  assign P91[14] = IN1[44]&IN2[47];
  assign P92[13] = IN1[44]&IN2[48];
  assign P93[12] = IN1[44]&IN2[49];
  assign P94[11] = IN1[44]&IN2[50];
  assign P95[10] = IN1[44]&IN2[51];
  assign P96[9] = IN1[44]&IN2[52];
  assign P97[8] = IN1[44]&IN2[53];
  assign P98[7] = IN1[44]&IN2[54];
  assign P99[6] = IN1[44]&IN2[55];
  assign P100[5] = IN1[44]&IN2[56];
  assign P101[4] = IN1[44]&IN2[57];
  assign P102[3] = IN1[44]&IN2[58];
  assign P103[2] = IN1[44]&IN2[59];
  assign P104[1] = IN1[44]&IN2[60];
  assign P105[0] = IN1[44]&IN2[61];
  assign P45[45] = IN1[45]&IN2[0];
  assign P46[45] = IN1[45]&IN2[1];
  assign P47[45] = IN1[45]&IN2[2];
  assign P48[45] = IN1[45]&IN2[3];
  assign P49[45] = IN1[45]&IN2[4];
  assign P50[45] = IN1[45]&IN2[5];
  assign P51[45] = IN1[45]&IN2[6];
  assign P52[45] = IN1[45]&IN2[7];
  assign P53[45] = IN1[45]&IN2[8];
  assign P54[45] = IN1[45]&IN2[9];
  assign P55[45] = IN1[45]&IN2[10];
  assign P56[45] = IN1[45]&IN2[11];
  assign P57[45] = IN1[45]&IN2[12];
  assign P58[45] = IN1[45]&IN2[13];
  assign P59[45] = IN1[45]&IN2[14];
  assign P60[45] = IN1[45]&IN2[15];
  assign P61[45] = IN1[45]&IN2[16];
  assign P62[44] = IN1[45]&IN2[17];
  assign P63[43] = IN1[45]&IN2[18];
  assign P64[42] = IN1[45]&IN2[19];
  assign P65[41] = IN1[45]&IN2[20];
  assign P66[40] = IN1[45]&IN2[21];
  assign P67[39] = IN1[45]&IN2[22];
  assign P68[38] = IN1[45]&IN2[23];
  assign P69[37] = IN1[45]&IN2[24];
  assign P70[36] = IN1[45]&IN2[25];
  assign P71[35] = IN1[45]&IN2[26];
  assign P72[34] = IN1[45]&IN2[27];
  assign P73[33] = IN1[45]&IN2[28];
  assign P74[32] = IN1[45]&IN2[29];
  assign P75[31] = IN1[45]&IN2[30];
  assign P76[30] = IN1[45]&IN2[31];
  assign P77[29] = IN1[45]&IN2[32];
  assign P78[28] = IN1[45]&IN2[33];
  assign P79[27] = IN1[45]&IN2[34];
  assign P80[26] = IN1[45]&IN2[35];
  assign P81[25] = IN1[45]&IN2[36];
  assign P82[24] = IN1[45]&IN2[37];
  assign P83[23] = IN1[45]&IN2[38];
  assign P84[22] = IN1[45]&IN2[39];
  assign P85[21] = IN1[45]&IN2[40];
  assign P86[20] = IN1[45]&IN2[41];
  assign P87[19] = IN1[45]&IN2[42];
  assign P88[18] = IN1[45]&IN2[43];
  assign P89[17] = IN1[45]&IN2[44];
  assign P90[16] = IN1[45]&IN2[45];
  assign P91[15] = IN1[45]&IN2[46];
  assign P92[14] = IN1[45]&IN2[47];
  assign P93[13] = IN1[45]&IN2[48];
  assign P94[12] = IN1[45]&IN2[49];
  assign P95[11] = IN1[45]&IN2[50];
  assign P96[10] = IN1[45]&IN2[51];
  assign P97[9] = IN1[45]&IN2[52];
  assign P98[8] = IN1[45]&IN2[53];
  assign P99[7] = IN1[45]&IN2[54];
  assign P100[6] = IN1[45]&IN2[55];
  assign P101[5] = IN1[45]&IN2[56];
  assign P102[4] = IN1[45]&IN2[57];
  assign P103[3] = IN1[45]&IN2[58];
  assign P104[2] = IN1[45]&IN2[59];
  assign P105[1] = IN1[45]&IN2[60];
  assign P106[0] = IN1[45]&IN2[61];
  assign P46[46] = IN1[46]&IN2[0];
  assign P47[46] = IN1[46]&IN2[1];
  assign P48[46] = IN1[46]&IN2[2];
  assign P49[46] = IN1[46]&IN2[3];
  assign P50[46] = IN1[46]&IN2[4];
  assign P51[46] = IN1[46]&IN2[5];
  assign P52[46] = IN1[46]&IN2[6];
  assign P53[46] = IN1[46]&IN2[7];
  assign P54[46] = IN1[46]&IN2[8];
  assign P55[46] = IN1[46]&IN2[9];
  assign P56[46] = IN1[46]&IN2[10];
  assign P57[46] = IN1[46]&IN2[11];
  assign P58[46] = IN1[46]&IN2[12];
  assign P59[46] = IN1[46]&IN2[13];
  assign P60[46] = IN1[46]&IN2[14];
  assign P61[46] = IN1[46]&IN2[15];
  assign P62[45] = IN1[46]&IN2[16];
  assign P63[44] = IN1[46]&IN2[17];
  assign P64[43] = IN1[46]&IN2[18];
  assign P65[42] = IN1[46]&IN2[19];
  assign P66[41] = IN1[46]&IN2[20];
  assign P67[40] = IN1[46]&IN2[21];
  assign P68[39] = IN1[46]&IN2[22];
  assign P69[38] = IN1[46]&IN2[23];
  assign P70[37] = IN1[46]&IN2[24];
  assign P71[36] = IN1[46]&IN2[25];
  assign P72[35] = IN1[46]&IN2[26];
  assign P73[34] = IN1[46]&IN2[27];
  assign P74[33] = IN1[46]&IN2[28];
  assign P75[32] = IN1[46]&IN2[29];
  assign P76[31] = IN1[46]&IN2[30];
  assign P77[30] = IN1[46]&IN2[31];
  assign P78[29] = IN1[46]&IN2[32];
  assign P79[28] = IN1[46]&IN2[33];
  assign P80[27] = IN1[46]&IN2[34];
  assign P81[26] = IN1[46]&IN2[35];
  assign P82[25] = IN1[46]&IN2[36];
  assign P83[24] = IN1[46]&IN2[37];
  assign P84[23] = IN1[46]&IN2[38];
  assign P85[22] = IN1[46]&IN2[39];
  assign P86[21] = IN1[46]&IN2[40];
  assign P87[20] = IN1[46]&IN2[41];
  assign P88[19] = IN1[46]&IN2[42];
  assign P89[18] = IN1[46]&IN2[43];
  assign P90[17] = IN1[46]&IN2[44];
  assign P91[16] = IN1[46]&IN2[45];
  assign P92[15] = IN1[46]&IN2[46];
  assign P93[14] = IN1[46]&IN2[47];
  assign P94[13] = IN1[46]&IN2[48];
  assign P95[12] = IN1[46]&IN2[49];
  assign P96[11] = IN1[46]&IN2[50];
  assign P97[10] = IN1[46]&IN2[51];
  assign P98[9] = IN1[46]&IN2[52];
  assign P99[8] = IN1[46]&IN2[53];
  assign P100[7] = IN1[46]&IN2[54];
  assign P101[6] = IN1[46]&IN2[55];
  assign P102[5] = IN1[46]&IN2[56];
  assign P103[4] = IN1[46]&IN2[57];
  assign P104[3] = IN1[46]&IN2[58];
  assign P105[2] = IN1[46]&IN2[59];
  assign P106[1] = IN1[46]&IN2[60];
  assign P107[0] = IN1[46]&IN2[61];
  assign P47[47] = IN1[47]&IN2[0];
  assign P48[47] = IN1[47]&IN2[1];
  assign P49[47] = IN1[47]&IN2[2];
  assign P50[47] = IN1[47]&IN2[3];
  assign P51[47] = IN1[47]&IN2[4];
  assign P52[47] = IN1[47]&IN2[5];
  assign P53[47] = IN1[47]&IN2[6];
  assign P54[47] = IN1[47]&IN2[7];
  assign P55[47] = IN1[47]&IN2[8];
  assign P56[47] = IN1[47]&IN2[9];
  assign P57[47] = IN1[47]&IN2[10];
  assign P58[47] = IN1[47]&IN2[11];
  assign P59[47] = IN1[47]&IN2[12];
  assign P60[47] = IN1[47]&IN2[13];
  assign P61[47] = IN1[47]&IN2[14];
  assign P62[46] = IN1[47]&IN2[15];
  assign P63[45] = IN1[47]&IN2[16];
  assign P64[44] = IN1[47]&IN2[17];
  assign P65[43] = IN1[47]&IN2[18];
  assign P66[42] = IN1[47]&IN2[19];
  assign P67[41] = IN1[47]&IN2[20];
  assign P68[40] = IN1[47]&IN2[21];
  assign P69[39] = IN1[47]&IN2[22];
  assign P70[38] = IN1[47]&IN2[23];
  assign P71[37] = IN1[47]&IN2[24];
  assign P72[36] = IN1[47]&IN2[25];
  assign P73[35] = IN1[47]&IN2[26];
  assign P74[34] = IN1[47]&IN2[27];
  assign P75[33] = IN1[47]&IN2[28];
  assign P76[32] = IN1[47]&IN2[29];
  assign P77[31] = IN1[47]&IN2[30];
  assign P78[30] = IN1[47]&IN2[31];
  assign P79[29] = IN1[47]&IN2[32];
  assign P80[28] = IN1[47]&IN2[33];
  assign P81[27] = IN1[47]&IN2[34];
  assign P82[26] = IN1[47]&IN2[35];
  assign P83[25] = IN1[47]&IN2[36];
  assign P84[24] = IN1[47]&IN2[37];
  assign P85[23] = IN1[47]&IN2[38];
  assign P86[22] = IN1[47]&IN2[39];
  assign P87[21] = IN1[47]&IN2[40];
  assign P88[20] = IN1[47]&IN2[41];
  assign P89[19] = IN1[47]&IN2[42];
  assign P90[18] = IN1[47]&IN2[43];
  assign P91[17] = IN1[47]&IN2[44];
  assign P92[16] = IN1[47]&IN2[45];
  assign P93[15] = IN1[47]&IN2[46];
  assign P94[14] = IN1[47]&IN2[47];
  assign P95[13] = IN1[47]&IN2[48];
  assign P96[12] = IN1[47]&IN2[49];
  assign P97[11] = IN1[47]&IN2[50];
  assign P98[10] = IN1[47]&IN2[51];
  assign P99[9] = IN1[47]&IN2[52];
  assign P100[8] = IN1[47]&IN2[53];
  assign P101[7] = IN1[47]&IN2[54];
  assign P102[6] = IN1[47]&IN2[55];
  assign P103[5] = IN1[47]&IN2[56];
  assign P104[4] = IN1[47]&IN2[57];
  assign P105[3] = IN1[47]&IN2[58];
  assign P106[2] = IN1[47]&IN2[59];
  assign P107[1] = IN1[47]&IN2[60];
  assign P108[0] = IN1[47]&IN2[61];
  assign P48[48] = IN1[48]&IN2[0];
  assign P49[48] = IN1[48]&IN2[1];
  assign P50[48] = IN1[48]&IN2[2];
  assign P51[48] = IN1[48]&IN2[3];
  assign P52[48] = IN1[48]&IN2[4];
  assign P53[48] = IN1[48]&IN2[5];
  assign P54[48] = IN1[48]&IN2[6];
  assign P55[48] = IN1[48]&IN2[7];
  assign P56[48] = IN1[48]&IN2[8];
  assign P57[48] = IN1[48]&IN2[9];
  assign P58[48] = IN1[48]&IN2[10];
  assign P59[48] = IN1[48]&IN2[11];
  assign P60[48] = IN1[48]&IN2[12];
  assign P61[48] = IN1[48]&IN2[13];
  assign P62[47] = IN1[48]&IN2[14];
  assign P63[46] = IN1[48]&IN2[15];
  assign P64[45] = IN1[48]&IN2[16];
  assign P65[44] = IN1[48]&IN2[17];
  assign P66[43] = IN1[48]&IN2[18];
  assign P67[42] = IN1[48]&IN2[19];
  assign P68[41] = IN1[48]&IN2[20];
  assign P69[40] = IN1[48]&IN2[21];
  assign P70[39] = IN1[48]&IN2[22];
  assign P71[38] = IN1[48]&IN2[23];
  assign P72[37] = IN1[48]&IN2[24];
  assign P73[36] = IN1[48]&IN2[25];
  assign P74[35] = IN1[48]&IN2[26];
  assign P75[34] = IN1[48]&IN2[27];
  assign P76[33] = IN1[48]&IN2[28];
  assign P77[32] = IN1[48]&IN2[29];
  assign P78[31] = IN1[48]&IN2[30];
  assign P79[30] = IN1[48]&IN2[31];
  assign P80[29] = IN1[48]&IN2[32];
  assign P81[28] = IN1[48]&IN2[33];
  assign P82[27] = IN1[48]&IN2[34];
  assign P83[26] = IN1[48]&IN2[35];
  assign P84[25] = IN1[48]&IN2[36];
  assign P85[24] = IN1[48]&IN2[37];
  assign P86[23] = IN1[48]&IN2[38];
  assign P87[22] = IN1[48]&IN2[39];
  assign P88[21] = IN1[48]&IN2[40];
  assign P89[20] = IN1[48]&IN2[41];
  assign P90[19] = IN1[48]&IN2[42];
  assign P91[18] = IN1[48]&IN2[43];
  assign P92[17] = IN1[48]&IN2[44];
  assign P93[16] = IN1[48]&IN2[45];
  assign P94[15] = IN1[48]&IN2[46];
  assign P95[14] = IN1[48]&IN2[47];
  assign P96[13] = IN1[48]&IN2[48];
  assign P97[12] = IN1[48]&IN2[49];
  assign P98[11] = IN1[48]&IN2[50];
  assign P99[10] = IN1[48]&IN2[51];
  assign P100[9] = IN1[48]&IN2[52];
  assign P101[8] = IN1[48]&IN2[53];
  assign P102[7] = IN1[48]&IN2[54];
  assign P103[6] = IN1[48]&IN2[55];
  assign P104[5] = IN1[48]&IN2[56];
  assign P105[4] = IN1[48]&IN2[57];
  assign P106[3] = IN1[48]&IN2[58];
  assign P107[2] = IN1[48]&IN2[59];
  assign P108[1] = IN1[48]&IN2[60];
  assign P109[0] = IN1[48]&IN2[61];
  assign P49[49] = IN1[49]&IN2[0];
  assign P50[49] = IN1[49]&IN2[1];
  assign P51[49] = IN1[49]&IN2[2];
  assign P52[49] = IN1[49]&IN2[3];
  assign P53[49] = IN1[49]&IN2[4];
  assign P54[49] = IN1[49]&IN2[5];
  assign P55[49] = IN1[49]&IN2[6];
  assign P56[49] = IN1[49]&IN2[7];
  assign P57[49] = IN1[49]&IN2[8];
  assign P58[49] = IN1[49]&IN2[9];
  assign P59[49] = IN1[49]&IN2[10];
  assign P60[49] = IN1[49]&IN2[11];
  assign P61[49] = IN1[49]&IN2[12];
  assign P62[48] = IN1[49]&IN2[13];
  assign P63[47] = IN1[49]&IN2[14];
  assign P64[46] = IN1[49]&IN2[15];
  assign P65[45] = IN1[49]&IN2[16];
  assign P66[44] = IN1[49]&IN2[17];
  assign P67[43] = IN1[49]&IN2[18];
  assign P68[42] = IN1[49]&IN2[19];
  assign P69[41] = IN1[49]&IN2[20];
  assign P70[40] = IN1[49]&IN2[21];
  assign P71[39] = IN1[49]&IN2[22];
  assign P72[38] = IN1[49]&IN2[23];
  assign P73[37] = IN1[49]&IN2[24];
  assign P74[36] = IN1[49]&IN2[25];
  assign P75[35] = IN1[49]&IN2[26];
  assign P76[34] = IN1[49]&IN2[27];
  assign P77[33] = IN1[49]&IN2[28];
  assign P78[32] = IN1[49]&IN2[29];
  assign P79[31] = IN1[49]&IN2[30];
  assign P80[30] = IN1[49]&IN2[31];
  assign P81[29] = IN1[49]&IN2[32];
  assign P82[28] = IN1[49]&IN2[33];
  assign P83[27] = IN1[49]&IN2[34];
  assign P84[26] = IN1[49]&IN2[35];
  assign P85[25] = IN1[49]&IN2[36];
  assign P86[24] = IN1[49]&IN2[37];
  assign P87[23] = IN1[49]&IN2[38];
  assign P88[22] = IN1[49]&IN2[39];
  assign P89[21] = IN1[49]&IN2[40];
  assign P90[20] = IN1[49]&IN2[41];
  assign P91[19] = IN1[49]&IN2[42];
  assign P92[18] = IN1[49]&IN2[43];
  assign P93[17] = IN1[49]&IN2[44];
  assign P94[16] = IN1[49]&IN2[45];
  assign P95[15] = IN1[49]&IN2[46];
  assign P96[14] = IN1[49]&IN2[47];
  assign P97[13] = IN1[49]&IN2[48];
  assign P98[12] = IN1[49]&IN2[49];
  assign P99[11] = IN1[49]&IN2[50];
  assign P100[10] = IN1[49]&IN2[51];
  assign P101[9] = IN1[49]&IN2[52];
  assign P102[8] = IN1[49]&IN2[53];
  assign P103[7] = IN1[49]&IN2[54];
  assign P104[6] = IN1[49]&IN2[55];
  assign P105[5] = IN1[49]&IN2[56];
  assign P106[4] = IN1[49]&IN2[57];
  assign P107[3] = IN1[49]&IN2[58];
  assign P108[2] = IN1[49]&IN2[59];
  assign P109[1] = IN1[49]&IN2[60];
  assign P110[0] = IN1[49]&IN2[61];
  assign P50[50] = IN1[50]&IN2[0];
  assign P51[50] = IN1[50]&IN2[1];
  assign P52[50] = IN1[50]&IN2[2];
  assign P53[50] = IN1[50]&IN2[3];
  assign P54[50] = IN1[50]&IN2[4];
  assign P55[50] = IN1[50]&IN2[5];
  assign P56[50] = IN1[50]&IN2[6];
  assign P57[50] = IN1[50]&IN2[7];
  assign P58[50] = IN1[50]&IN2[8];
  assign P59[50] = IN1[50]&IN2[9];
  assign P60[50] = IN1[50]&IN2[10];
  assign P61[50] = IN1[50]&IN2[11];
  assign P62[49] = IN1[50]&IN2[12];
  assign P63[48] = IN1[50]&IN2[13];
  assign P64[47] = IN1[50]&IN2[14];
  assign P65[46] = IN1[50]&IN2[15];
  assign P66[45] = IN1[50]&IN2[16];
  assign P67[44] = IN1[50]&IN2[17];
  assign P68[43] = IN1[50]&IN2[18];
  assign P69[42] = IN1[50]&IN2[19];
  assign P70[41] = IN1[50]&IN2[20];
  assign P71[40] = IN1[50]&IN2[21];
  assign P72[39] = IN1[50]&IN2[22];
  assign P73[38] = IN1[50]&IN2[23];
  assign P74[37] = IN1[50]&IN2[24];
  assign P75[36] = IN1[50]&IN2[25];
  assign P76[35] = IN1[50]&IN2[26];
  assign P77[34] = IN1[50]&IN2[27];
  assign P78[33] = IN1[50]&IN2[28];
  assign P79[32] = IN1[50]&IN2[29];
  assign P80[31] = IN1[50]&IN2[30];
  assign P81[30] = IN1[50]&IN2[31];
  assign P82[29] = IN1[50]&IN2[32];
  assign P83[28] = IN1[50]&IN2[33];
  assign P84[27] = IN1[50]&IN2[34];
  assign P85[26] = IN1[50]&IN2[35];
  assign P86[25] = IN1[50]&IN2[36];
  assign P87[24] = IN1[50]&IN2[37];
  assign P88[23] = IN1[50]&IN2[38];
  assign P89[22] = IN1[50]&IN2[39];
  assign P90[21] = IN1[50]&IN2[40];
  assign P91[20] = IN1[50]&IN2[41];
  assign P92[19] = IN1[50]&IN2[42];
  assign P93[18] = IN1[50]&IN2[43];
  assign P94[17] = IN1[50]&IN2[44];
  assign P95[16] = IN1[50]&IN2[45];
  assign P96[15] = IN1[50]&IN2[46];
  assign P97[14] = IN1[50]&IN2[47];
  assign P98[13] = IN1[50]&IN2[48];
  assign P99[12] = IN1[50]&IN2[49];
  assign P100[11] = IN1[50]&IN2[50];
  assign P101[10] = IN1[50]&IN2[51];
  assign P102[9] = IN1[50]&IN2[52];
  assign P103[8] = IN1[50]&IN2[53];
  assign P104[7] = IN1[50]&IN2[54];
  assign P105[6] = IN1[50]&IN2[55];
  assign P106[5] = IN1[50]&IN2[56];
  assign P107[4] = IN1[50]&IN2[57];
  assign P108[3] = IN1[50]&IN2[58];
  assign P109[2] = IN1[50]&IN2[59];
  assign P110[1] = IN1[50]&IN2[60];
  assign P111[0] = IN1[50]&IN2[61];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, IN79, IN80, IN81, IN82, IN83, IN84, IN85, IN86, IN87, IN88, IN89, IN90, IN91, IN92, IN93, IN94, IN95, IN96, IN97, IN98, IN99, IN100, IN101, IN102, IN103, IN104, IN105, IN106, IN107, IN108, IN109, IN110, IN111, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [29:0] IN29;
  input [30:0] IN30;
  input [31:0] IN31;
  input [32:0] IN32;
  input [33:0] IN33;
  input [34:0] IN34;
  input [35:0] IN35;
  input [36:0] IN36;
  input [37:0] IN37;
  input [38:0] IN38;
  input [39:0] IN39;
  input [40:0] IN40;
  input [41:0] IN41;
  input [42:0] IN42;
  input [43:0] IN43;
  input [44:0] IN44;
  input [45:0] IN45;
  input [46:0] IN46;
  input [47:0] IN47;
  input [48:0] IN48;
  input [49:0] IN49;
  input [50:0] IN50;
  input [50:0] IN51;
  input [50:0] IN52;
  input [50:0] IN53;
  input [50:0] IN54;
  input [50:0] IN55;
  input [50:0] IN56;
  input [50:0] IN57;
  input [50:0] IN58;
  input [50:0] IN59;
  input [50:0] IN60;
  input [50:0] IN61;
  input [49:0] IN62;
  input [48:0] IN63;
  input [47:0] IN64;
  input [46:0] IN65;
  input [45:0] IN66;
  input [44:0] IN67;
  input [43:0] IN68;
  input [42:0] IN69;
  input [41:0] IN70;
  input [40:0] IN71;
  input [39:0] IN72;
  input [38:0] IN73;
  input [37:0] IN74;
  input [36:0] IN75;
  input [35:0] IN76;
  input [34:0] IN77;
  input [33:0] IN78;
  input [32:0] IN79;
  input [31:0] IN80;
  input [30:0] IN81;
  input [29:0] IN82;
  input [28:0] IN83;
  input [27:0] IN84;
  input [26:0] IN85;
  input [25:0] IN86;
  input [24:0] IN87;
  input [23:0] IN88;
  input [22:0] IN89;
  input [21:0] IN90;
  input [20:0] IN91;
  input [19:0] IN92;
  input [18:0] IN93;
  input [17:0] IN94;
  input [16:0] IN95;
  input [15:0] IN96;
  input [14:0] IN97;
  input [13:0] IN98;
  input [12:0] IN99;
  input [11:0] IN100;
  input [10:0] IN101;
  input [9:0] IN102;
  input [8:0] IN103;
  input [7:0] IN104;
  input [6:0] IN105;
  input [5:0] IN106;
  input [4:0] IN107;
  input [3:0] IN108;
  input [2:0] IN109;
  input [1:0] IN110;
  input [0:0] IN111;
  output [111:0] Out1;
  output [60:0] Out2;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3225;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3254;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3272;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3285;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3327;
  wire w3328;
  wire w3329;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3334;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3366;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3385;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3414;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3433;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3443;
  wire w3444;
  wire w3445;
  wire w3446;
  wire w3447;
  wire w3448;
  wire w3449;
  wire w3450;
  wire w3451;
  wire w3452;
  wire w3453;
  wire w3454;
  wire w3455;
  wire w3456;
  wire w3457;
  wire w3458;
  wire w3459;
  wire w3460;
  wire w3461;
  wire w3463;
  wire w3464;
  wire w3465;
  wire w3466;
  wire w3467;
  wire w3468;
  wire w3469;
  wire w3470;
  wire w3471;
  wire w3472;
  wire w3473;
  wire w3474;
  wire w3475;
  wire w3476;
  wire w3477;
  wire w3478;
  wire w3479;
  wire w3480;
  wire w3481;
  wire w3482;
  wire w3483;
  wire w3484;
  wire w3485;
  wire w3486;
  wire w3487;
  wire w3488;
  wire w3489;
  wire w3490;
  wire w3491;
  wire w3492;
  wire w3493;
  wire w3494;
  wire w3495;
  wire w3496;
  wire w3497;
  wire w3498;
  wire w3499;
  wire w3500;
  wire w3501;
  wire w3502;
  wire w3503;
  wire w3504;
  wire w3505;
  wire w3506;
  wire w3507;
  wire w3508;
  wire w3509;
  wire w3510;
  wire w3511;
  wire w3512;
  wire w3513;
  wire w3514;
  wire w3515;
  wire w3516;
  wire w3517;
  wire w3518;
  wire w3519;
  wire w3520;
  wire w3521;
  wire w3522;
  wire w3523;
  wire w3524;
  wire w3525;
  wire w3526;
  wire w3527;
  wire w3528;
  wire w3529;
  wire w3530;
  wire w3531;
  wire w3532;
  wire w3533;
  wire w3534;
  wire w3535;
  wire w3536;
  wire w3537;
  wire w3538;
  wire w3539;
  wire w3540;
  wire w3541;
  wire w3542;
  wire w3543;
  wire w3544;
  wire w3545;
  wire w3546;
  wire w3547;
  wire w3548;
  wire w3549;
  wire w3550;
  wire w3551;
  wire w3552;
  wire w3553;
  wire w3554;
  wire w3555;
  wire w3556;
  wire w3557;
  wire w3558;
  wire w3559;
  wire w3560;
  wire w3561;
  wire w3563;
  wire w3564;
  wire w3565;
  wire w3566;
  wire w3567;
  wire w3568;
  wire w3569;
  wire w3570;
  wire w3571;
  wire w3572;
  wire w3573;
  wire w3574;
  wire w3575;
  wire w3576;
  wire w3577;
  wire w3578;
  wire w3579;
  wire w3580;
  wire w3581;
  wire w3582;
  wire w3583;
  wire w3584;
  wire w3585;
  wire w3586;
  wire w3587;
  wire w3588;
  wire w3589;
  wire w3590;
  wire w3591;
  wire w3592;
  wire w3593;
  wire w3594;
  wire w3595;
  wire w3596;
  wire w3597;
  wire w3598;
  wire w3599;
  wire w3600;
  wire w3601;
  wire w3602;
  wire w3603;
  wire w3604;
  wire w3605;
  wire w3606;
  wire w3607;
  wire w3608;
  wire w3609;
  wire w3610;
  wire w3611;
  wire w3612;
  wire w3613;
  wire w3614;
  wire w3615;
  wire w3616;
  wire w3617;
  wire w3618;
  wire w3619;
  wire w3620;
  wire w3621;
  wire w3622;
  wire w3623;
  wire w3624;
  wire w3625;
  wire w3626;
  wire w3627;
  wire w3628;
  wire w3629;
  wire w3630;
  wire w3631;
  wire w3632;
  wire w3633;
  wire w3634;
  wire w3635;
  wire w3636;
  wire w3637;
  wire w3638;
  wire w3639;
  wire w3640;
  wire w3641;
  wire w3642;
  wire w3643;
  wire w3644;
  wire w3645;
  wire w3646;
  wire w3647;
  wire w3648;
  wire w3649;
  wire w3650;
  wire w3651;
  wire w3652;
  wire w3653;
  wire w3654;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3685;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3734;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3742;
  wire w3743;
  wire w3744;
  wire w3745;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3768;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3785;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3814;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3836;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3849;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3882;
  wire w3883;
  wire w3884;
  wire w3885;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3894;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3930;
  wire w3931;
  wire w3932;
  wire w3933;
  wire w3934;
  wire w3935;
  wire w3936;
  wire w3937;
  wire w3938;
  wire w3939;
  wire w3940;
  wire w3941;
  wire w3942;
  wire w3943;
  wire w3944;
  wire w3945;
  wire w3946;
  wire w3947;
  wire w3948;
  wire w3949;
  wire w3950;
  wire w3951;
  wire w3952;
  wire w3953;
  wire w3954;
  wire w3955;
  wire w3956;
  wire w3957;
  wire w3958;
  wire w3959;
  wire w3960;
  wire w3961;
  wire w3963;
  wire w3964;
  wire w3965;
  wire w3966;
  wire w3967;
  wire w3968;
  wire w3969;
  wire w3970;
  wire w3971;
  wire w3972;
  wire w3973;
  wire w3974;
  wire w3975;
  wire w3976;
  wire w3977;
  wire w3978;
  wire w3979;
  wire w3980;
  wire w3981;
  wire w3982;
  wire w3983;
  wire w3984;
  wire w3985;
  wire w3986;
  wire w3987;
  wire w3988;
  wire w3989;
  wire w3990;
  wire w3991;
  wire w3992;
  wire w3993;
  wire w3994;
  wire w3995;
  wire w3996;
  wire w3997;
  wire w3998;
  wire w3999;
  wire w4000;
  wire w4001;
  wire w4002;
  wire w4003;
  wire w4004;
  wire w4005;
  wire w4006;
  wire w4007;
  wire w4008;
  wire w4009;
  wire w4010;
  wire w4011;
  wire w4012;
  wire w4013;
  wire w4014;
  wire w4015;
  wire w4016;
  wire w4017;
  wire w4018;
  wire w4019;
  wire w4020;
  wire w4021;
  wire w4022;
  wire w4023;
  wire w4024;
  wire w4025;
  wire w4026;
  wire w4027;
  wire w4028;
  wire w4029;
  wire w4030;
  wire w4031;
  wire w4032;
  wire w4033;
  wire w4034;
  wire w4035;
  wire w4036;
  wire w4037;
  wire w4038;
  wire w4039;
  wire w4040;
  wire w4041;
  wire w4042;
  wire w4043;
  wire w4044;
  wire w4045;
  wire w4046;
  wire w4047;
  wire w4048;
  wire w4049;
  wire w4050;
  wire w4051;
  wire w4052;
  wire w4053;
  wire w4054;
  wire w4055;
  wire w4056;
  wire w4057;
  wire w4058;
  wire w4059;
  wire w4060;
  wire w4061;
  wire w4063;
  wire w4064;
  wire w4065;
  wire w4066;
  wire w4067;
  wire w4068;
  wire w4069;
  wire w4070;
  wire w4071;
  wire w4072;
  wire w4073;
  wire w4074;
  wire w4075;
  wire w4076;
  wire w4077;
  wire w4078;
  wire w4079;
  wire w4080;
  wire w4081;
  wire w4082;
  wire w4083;
  wire w4084;
  wire w4085;
  wire w4086;
  wire w4087;
  wire w4088;
  wire w4089;
  wire w4090;
  wire w4091;
  wire w4092;
  wire w4093;
  wire w4094;
  wire w4095;
  wire w4096;
  wire w4097;
  wire w4098;
  wire w4099;
  wire w4100;
  wire w4101;
  wire w4102;
  wire w4103;
  wire w4104;
  wire w4105;
  wire w4106;
  wire w4107;
  wire w4108;
  wire w4109;
  wire w4110;
  wire w4111;
  wire w4112;
  wire w4113;
  wire w4114;
  wire w4115;
  wire w4116;
  wire w4117;
  wire w4118;
  wire w4119;
  wire w4120;
  wire w4121;
  wire w4122;
  wire w4123;
  wire w4124;
  wire w4125;
  wire w4126;
  wire w4127;
  wire w4128;
  wire w4129;
  wire w4130;
  wire w4131;
  wire w4132;
  wire w4133;
  wire w4134;
  wire w4135;
  wire w4136;
  wire w4137;
  wire w4138;
  wire w4139;
  wire w4140;
  wire w4141;
  wire w4142;
  wire w4143;
  wire w4144;
  wire w4145;
  wire w4146;
  wire w4147;
  wire w4148;
  wire w4149;
  wire w4150;
  wire w4151;
  wire w4152;
  wire w4153;
  wire w4154;
  wire w4155;
  wire w4156;
  wire w4157;
  wire w4158;
  wire w4159;
  wire w4160;
  wire w4161;
  wire w4163;
  wire w4164;
  wire w4165;
  wire w4166;
  wire w4167;
  wire w4168;
  wire w4169;
  wire w4170;
  wire w4171;
  wire w4172;
  wire w4173;
  wire w4174;
  wire w4175;
  wire w4176;
  wire w4177;
  wire w4178;
  wire w4179;
  wire w4180;
  wire w4181;
  wire w4182;
  wire w4183;
  wire w4184;
  wire w4185;
  wire w4186;
  wire w4187;
  wire w4188;
  wire w4189;
  wire w4190;
  wire w4191;
  wire w4192;
  wire w4193;
  wire w4194;
  wire w4195;
  wire w4196;
  wire w4197;
  wire w4198;
  wire w4199;
  wire w4200;
  wire w4201;
  wire w4202;
  wire w4203;
  wire w4204;
  wire w4205;
  wire w4206;
  wire w4207;
  wire w4208;
  wire w4209;
  wire w4210;
  wire w4211;
  wire w4212;
  wire w4213;
  wire w4214;
  wire w4215;
  wire w4216;
  wire w4217;
  wire w4218;
  wire w4219;
  wire w4220;
  wire w4221;
  wire w4222;
  wire w4223;
  wire w4224;
  wire w4225;
  wire w4226;
  wire w4227;
  wire w4228;
  wire w4229;
  wire w4230;
  wire w4231;
  wire w4232;
  wire w4233;
  wire w4234;
  wire w4235;
  wire w4236;
  wire w4237;
  wire w4238;
  wire w4239;
  wire w4240;
  wire w4241;
  wire w4242;
  wire w4243;
  wire w4244;
  wire w4245;
  wire w4246;
  wire w4247;
  wire w4248;
  wire w4249;
  wire w4250;
  wire w4251;
  wire w4252;
  wire w4253;
  wire w4254;
  wire w4255;
  wire w4256;
  wire w4257;
  wire w4258;
  wire w4259;
  wire w4260;
  wire w4261;
  wire w4263;
  wire w4264;
  wire w4265;
  wire w4266;
  wire w4267;
  wire w4268;
  wire w4269;
  wire w4270;
  wire w4271;
  wire w4272;
  wire w4273;
  wire w4274;
  wire w4275;
  wire w4276;
  wire w4277;
  wire w4278;
  wire w4279;
  wire w4280;
  wire w4281;
  wire w4282;
  wire w4283;
  wire w4284;
  wire w4285;
  wire w4286;
  wire w4287;
  wire w4288;
  wire w4289;
  wire w4290;
  wire w4291;
  wire w4292;
  wire w4293;
  wire w4294;
  wire w4295;
  wire w4296;
  wire w4297;
  wire w4298;
  wire w4299;
  wire w4300;
  wire w4301;
  wire w4302;
  wire w4303;
  wire w4304;
  wire w4305;
  wire w4306;
  wire w4307;
  wire w4308;
  wire w4309;
  wire w4310;
  wire w4311;
  wire w4312;
  wire w4313;
  wire w4314;
  wire w4315;
  wire w4316;
  wire w4317;
  wire w4318;
  wire w4319;
  wire w4320;
  wire w4321;
  wire w4322;
  wire w4323;
  wire w4324;
  wire w4325;
  wire w4326;
  wire w4327;
  wire w4328;
  wire w4329;
  wire w4330;
  wire w4331;
  wire w4332;
  wire w4333;
  wire w4334;
  wire w4335;
  wire w4336;
  wire w4337;
  wire w4338;
  wire w4339;
  wire w4340;
  wire w4341;
  wire w4342;
  wire w4343;
  wire w4344;
  wire w4345;
  wire w4346;
  wire w4347;
  wire w4348;
  wire w4349;
  wire w4350;
  wire w4351;
  wire w4352;
  wire w4353;
  wire w4354;
  wire w4355;
  wire w4356;
  wire w4357;
  wire w4358;
  wire w4359;
  wire w4360;
  wire w4361;
  wire w4363;
  wire w4364;
  wire w4365;
  wire w4366;
  wire w4367;
  wire w4368;
  wire w4369;
  wire w4370;
  wire w4371;
  wire w4372;
  wire w4373;
  wire w4374;
  wire w4375;
  wire w4376;
  wire w4377;
  wire w4378;
  wire w4379;
  wire w4380;
  wire w4381;
  wire w4382;
  wire w4383;
  wire w4384;
  wire w4385;
  wire w4386;
  wire w4387;
  wire w4388;
  wire w4389;
  wire w4390;
  wire w4391;
  wire w4392;
  wire w4393;
  wire w4394;
  wire w4395;
  wire w4396;
  wire w4397;
  wire w4398;
  wire w4399;
  wire w4400;
  wire w4401;
  wire w4402;
  wire w4403;
  wire w4404;
  wire w4405;
  wire w4406;
  wire w4407;
  wire w4408;
  wire w4409;
  wire w4410;
  wire w4411;
  wire w4412;
  wire w4413;
  wire w4414;
  wire w4415;
  wire w4416;
  wire w4417;
  wire w4418;
  wire w4419;
  wire w4420;
  wire w4421;
  wire w4422;
  wire w4423;
  wire w4424;
  wire w4425;
  wire w4426;
  wire w4427;
  wire w4428;
  wire w4429;
  wire w4430;
  wire w4431;
  wire w4432;
  wire w4433;
  wire w4434;
  wire w4435;
  wire w4436;
  wire w4437;
  wire w4438;
  wire w4439;
  wire w4440;
  wire w4441;
  wire w4442;
  wire w4443;
  wire w4444;
  wire w4445;
  wire w4446;
  wire w4447;
  wire w4448;
  wire w4449;
  wire w4450;
  wire w4451;
  wire w4452;
  wire w4453;
  wire w4454;
  wire w4455;
  wire w4456;
  wire w4457;
  wire w4458;
  wire w4459;
  wire w4460;
  wire w4461;
  wire w4463;
  wire w4464;
  wire w4465;
  wire w4466;
  wire w4467;
  wire w4468;
  wire w4469;
  wire w4470;
  wire w4471;
  wire w4472;
  wire w4473;
  wire w4474;
  wire w4475;
  wire w4476;
  wire w4477;
  wire w4478;
  wire w4479;
  wire w4480;
  wire w4481;
  wire w4482;
  wire w4483;
  wire w4484;
  wire w4485;
  wire w4486;
  wire w4487;
  wire w4488;
  wire w4489;
  wire w4490;
  wire w4491;
  wire w4492;
  wire w4493;
  wire w4494;
  wire w4495;
  wire w4496;
  wire w4497;
  wire w4498;
  wire w4499;
  wire w4500;
  wire w4501;
  wire w4502;
  wire w4503;
  wire w4504;
  wire w4505;
  wire w4506;
  wire w4507;
  wire w4508;
  wire w4509;
  wire w4510;
  wire w4511;
  wire w4512;
  wire w4513;
  wire w4514;
  wire w4515;
  wire w4516;
  wire w4517;
  wire w4518;
  wire w4519;
  wire w4520;
  wire w4521;
  wire w4522;
  wire w4523;
  wire w4524;
  wire w4525;
  wire w4526;
  wire w4527;
  wire w4528;
  wire w4529;
  wire w4530;
  wire w4531;
  wire w4532;
  wire w4533;
  wire w4534;
  wire w4535;
  wire w4536;
  wire w4537;
  wire w4538;
  wire w4539;
  wire w4540;
  wire w4541;
  wire w4542;
  wire w4543;
  wire w4544;
  wire w4545;
  wire w4546;
  wire w4547;
  wire w4548;
  wire w4549;
  wire w4550;
  wire w4551;
  wire w4552;
  wire w4553;
  wire w4554;
  wire w4555;
  wire w4556;
  wire w4557;
  wire w4558;
  wire w4559;
  wire w4560;
  wire w4561;
  wire w4563;
  wire w4564;
  wire w4565;
  wire w4566;
  wire w4567;
  wire w4568;
  wire w4569;
  wire w4570;
  wire w4571;
  wire w4572;
  wire w4573;
  wire w4574;
  wire w4575;
  wire w4576;
  wire w4577;
  wire w4578;
  wire w4579;
  wire w4580;
  wire w4581;
  wire w4582;
  wire w4583;
  wire w4584;
  wire w4585;
  wire w4586;
  wire w4587;
  wire w4588;
  wire w4589;
  wire w4590;
  wire w4591;
  wire w4592;
  wire w4593;
  wire w4594;
  wire w4595;
  wire w4596;
  wire w4597;
  wire w4598;
  wire w4599;
  wire w4600;
  wire w4601;
  wire w4602;
  wire w4603;
  wire w4604;
  wire w4605;
  wire w4606;
  wire w4607;
  wire w4608;
  wire w4609;
  wire w4610;
  wire w4611;
  wire w4612;
  wire w4613;
  wire w4614;
  wire w4615;
  wire w4616;
  wire w4617;
  wire w4618;
  wire w4619;
  wire w4620;
  wire w4621;
  wire w4622;
  wire w4623;
  wire w4624;
  wire w4625;
  wire w4626;
  wire w4627;
  wire w4628;
  wire w4629;
  wire w4630;
  wire w4631;
  wire w4632;
  wire w4633;
  wire w4634;
  wire w4635;
  wire w4636;
  wire w4637;
  wire w4638;
  wire w4639;
  wire w4640;
  wire w4641;
  wire w4642;
  wire w4643;
  wire w4644;
  wire w4645;
  wire w4646;
  wire w4647;
  wire w4648;
  wire w4649;
  wire w4650;
  wire w4651;
  wire w4652;
  wire w4653;
  wire w4654;
  wire w4655;
  wire w4656;
  wire w4657;
  wire w4658;
  wire w4659;
  wire w4660;
  wire w4661;
  wire w4663;
  wire w4664;
  wire w4665;
  wire w4666;
  wire w4667;
  wire w4668;
  wire w4669;
  wire w4670;
  wire w4671;
  wire w4672;
  wire w4673;
  wire w4674;
  wire w4675;
  wire w4676;
  wire w4677;
  wire w4678;
  wire w4679;
  wire w4680;
  wire w4681;
  wire w4682;
  wire w4683;
  wire w4684;
  wire w4685;
  wire w4686;
  wire w4687;
  wire w4688;
  wire w4689;
  wire w4690;
  wire w4691;
  wire w4692;
  wire w4693;
  wire w4694;
  wire w4695;
  wire w4696;
  wire w4697;
  wire w4698;
  wire w4699;
  wire w4700;
  wire w4701;
  wire w4702;
  wire w4703;
  wire w4704;
  wire w4705;
  wire w4706;
  wire w4707;
  wire w4708;
  wire w4709;
  wire w4710;
  wire w4711;
  wire w4712;
  wire w4713;
  wire w4714;
  wire w4715;
  wire w4716;
  wire w4717;
  wire w4718;
  wire w4719;
  wire w4720;
  wire w4721;
  wire w4722;
  wire w4723;
  wire w4724;
  wire w4725;
  wire w4726;
  wire w4727;
  wire w4728;
  wire w4729;
  wire w4730;
  wire w4731;
  wire w4732;
  wire w4733;
  wire w4734;
  wire w4735;
  wire w4736;
  wire w4737;
  wire w4738;
  wire w4739;
  wire w4740;
  wire w4741;
  wire w4742;
  wire w4743;
  wire w4744;
  wire w4745;
  wire w4746;
  wire w4747;
  wire w4748;
  wire w4749;
  wire w4750;
  wire w4751;
  wire w4752;
  wire w4753;
  wire w4754;
  wire w4755;
  wire w4756;
  wire w4757;
  wire w4758;
  wire w4759;
  wire w4760;
  wire w4761;
  wire w4763;
  wire w4764;
  wire w4765;
  wire w4766;
  wire w4767;
  wire w4768;
  wire w4769;
  wire w4770;
  wire w4771;
  wire w4772;
  wire w4773;
  wire w4774;
  wire w4775;
  wire w4776;
  wire w4777;
  wire w4778;
  wire w4779;
  wire w4780;
  wire w4781;
  wire w4782;
  wire w4783;
  wire w4784;
  wire w4785;
  wire w4786;
  wire w4787;
  wire w4788;
  wire w4789;
  wire w4790;
  wire w4791;
  wire w4792;
  wire w4793;
  wire w4794;
  wire w4795;
  wire w4796;
  wire w4797;
  wire w4798;
  wire w4799;
  wire w4800;
  wire w4801;
  wire w4802;
  wire w4803;
  wire w4804;
  wire w4805;
  wire w4806;
  wire w4807;
  wire w4808;
  wire w4809;
  wire w4810;
  wire w4811;
  wire w4812;
  wire w4813;
  wire w4814;
  wire w4815;
  wire w4816;
  wire w4817;
  wire w4818;
  wire w4819;
  wire w4820;
  wire w4821;
  wire w4822;
  wire w4823;
  wire w4824;
  wire w4825;
  wire w4826;
  wire w4827;
  wire w4828;
  wire w4829;
  wire w4830;
  wire w4831;
  wire w4832;
  wire w4833;
  wire w4834;
  wire w4835;
  wire w4836;
  wire w4837;
  wire w4838;
  wire w4839;
  wire w4840;
  wire w4841;
  wire w4842;
  wire w4843;
  wire w4844;
  wire w4845;
  wire w4846;
  wire w4847;
  wire w4848;
  wire w4849;
  wire w4850;
  wire w4851;
  wire w4852;
  wire w4853;
  wire w4854;
  wire w4855;
  wire w4856;
  wire w4857;
  wire w4858;
  wire w4859;
  wire w4860;
  wire w4861;
  wire w4863;
  wire w4864;
  wire w4865;
  wire w4866;
  wire w4867;
  wire w4868;
  wire w4869;
  wire w4870;
  wire w4871;
  wire w4872;
  wire w4873;
  wire w4874;
  wire w4875;
  wire w4876;
  wire w4877;
  wire w4878;
  wire w4879;
  wire w4880;
  wire w4881;
  wire w4882;
  wire w4883;
  wire w4884;
  wire w4885;
  wire w4886;
  wire w4887;
  wire w4888;
  wire w4889;
  wire w4890;
  wire w4891;
  wire w4892;
  wire w4893;
  wire w4894;
  wire w4895;
  wire w4896;
  wire w4897;
  wire w4898;
  wire w4899;
  wire w4900;
  wire w4901;
  wire w4902;
  wire w4903;
  wire w4904;
  wire w4905;
  wire w4906;
  wire w4907;
  wire w4908;
  wire w4909;
  wire w4910;
  wire w4911;
  wire w4912;
  wire w4913;
  wire w4914;
  wire w4915;
  wire w4916;
  wire w4917;
  wire w4918;
  wire w4919;
  wire w4920;
  wire w4921;
  wire w4922;
  wire w4923;
  wire w4924;
  wire w4925;
  wire w4926;
  wire w4927;
  wire w4928;
  wire w4929;
  wire w4930;
  wire w4931;
  wire w4932;
  wire w4933;
  wire w4934;
  wire w4935;
  wire w4936;
  wire w4937;
  wire w4938;
  wire w4939;
  wire w4940;
  wire w4941;
  wire w4942;
  wire w4943;
  wire w4944;
  wire w4945;
  wire w4946;
  wire w4947;
  wire w4948;
  wire w4949;
  wire w4950;
  wire w4951;
  wire w4952;
  wire w4953;
  wire w4954;
  wire w4955;
  wire w4956;
  wire w4957;
  wire w4958;
  wire w4959;
  wire w4960;
  wire w4961;
  wire w4963;
  wire w4964;
  wire w4965;
  wire w4966;
  wire w4967;
  wire w4968;
  wire w4969;
  wire w4970;
  wire w4971;
  wire w4972;
  wire w4973;
  wire w4974;
  wire w4975;
  wire w4976;
  wire w4977;
  wire w4978;
  wire w4979;
  wire w4980;
  wire w4981;
  wire w4982;
  wire w4983;
  wire w4984;
  wire w4985;
  wire w4986;
  wire w4987;
  wire w4988;
  wire w4989;
  wire w4990;
  wire w4991;
  wire w4992;
  wire w4993;
  wire w4994;
  wire w4995;
  wire w4996;
  wire w4997;
  wire w4998;
  wire w4999;
  wire w5000;
  wire w5001;
  wire w5002;
  wire w5003;
  wire w5004;
  wire w5005;
  wire w5006;
  wire w5007;
  wire w5008;
  wire w5009;
  wire w5010;
  wire w5011;
  wire w5012;
  wire w5013;
  wire w5014;
  wire w5015;
  wire w5016;
  wire w5017;
  wire w5018;
  wire w5019;
  wire w5020;
  wire w5021;
  wire w5022;
  wire w5023;
  wire w5024;
  wire w5025;
  wire w5026;
  wire w5027;
  wire w5028;
  wire w5029;
  wire w5030;
  wire w5031;
  wire w5032;
  wire w5033;
  wire w5034;
  wire w5035;
  wire w5036;
  wire w5037;
  wire w5038;
  wire w5039;
  wire w5040;
  wire w5041;
  wire w5042;
  wire w5043;
  wire w5044;
  wire w5045;
  wire w5046;
  wire w5047;
  wire w5048;
  wire w5049;
  wire w5050;
  wire w5051;
  wire w5052;
  wire w5053;
  wire w5054;
  wire w5055;
  wire w5056;
  wire w5057;
  wire w5058;
  wire w5059;
  wire w5060;
  wire w5061;
  wire w5063;
  wire w5064;
  wire w5065;
  wire w5066;
  wire w5067;
  wire w5068;
  wire w5069;
  wire w5070;
  wire w5071;
  wire w5072;
  wire w5073;
  wire w5074;
  wire w5075;
  wire w5076;
  wire w5077;
  wire w5078;
  wire w5079;
  wire w5080;
  wire w5081;
  wire w5082;
  wire w5083;
  wire w5084;
  wire w5085;
  wire w5086;
  wire w5087;
  wire w5088;
  wire w5089;
  wire w5090;
  wire w5091;
  wire w5092;
  wire w5093;
  wire w5094;
  wire w5095;
  wire w5096;
  wire w5097;
  wire w5098;
  wire w5099;
  wire w5100;
  wire w5101;
  wire w5102;
  wire w5103;
  wire w5104;
  wire w5105;
  wire w5106;
  wire w5107;
  wire w5108;
  wire w5109;
  wire w5110;
  wire w5111;
  wire w5112;
  wire w5113;
  wire w5114;
  wire w5115;
  wire w5116;
  wire w5117;
  wire w5118;
  wire w5119;
  wire w5120;
  wire w5121;
  wire w5122;
  wire w5123;
  wire w5124;
  wire w5125;
  wire w5126;
  wire w5127;
  wire w5128;
  wire w5129;
  wire w5130;
  wire w5131;
  wire w5132;
  wire w5133;
  wire w5134;
  wire w5135;
  wire w5136;
  wire w5137;
  wire w5138;
  wire w5139;
  wire w5140;
  wire w5141;
  wire w5142;
  wire w5143;
  wire w5144;
  wire w5145;
  wire w5146;
  wire w5147;
  wire w5148;
  wire w5149;
  wire w5150;
  wire w5151;
  wire w5152;
  wire w5153;
  wire w5154;
  wire w5155;
  wire w5156;
  wire w5157;
  wire w5158;
  wire w5159;
  wire w5160;
  wire w5161;
  wire w5163;
  wire w5164;
  wire w5165;
  wire w5166;
  wire w5167;
  wire w5168;
  wire w5169;
  wire w5170;
  wire w5171;
  wire w5172;
  wire w5173;
  wire w5174;
  wire w5175;
  wire w5176;
  wire w5177;
  wire w5178;
  wire w5179;
  wire w5180;
  wire w5181;
  wire w5182;
  wire w5183;
  wire w5184;
  wire w5185;
  wire w5186;
  wire w5187;
  wire w5188;
  wire w5189;
  wire w5190;
  wire w5191;
  wire w5192;
  wire w5193;
  wire w5194;
  wire w5195;
  wire w5196;
  wire w5197;
  wire w5198;
  wire w5199;
  wire w5200;
  wire w5201;
  wire w5202;
  wire w5203;
  wire w5204;
  wire w5205;
  wire w5206;
  wire w5207;
  wire w5208;
  wire w5209;
  wire w5210;
  wire w5211;
  wire w5212;
  wire w5213;
  wire w5214;
  wire w5215;
  wire w5216;
  wire w5217;
  wire w5218;
  wire w5219;
  wire w5220;
  wire w5221;
  wire w5222;
  wire w5223;
  wire w5224;
  wire w5225;
  wire w5226;
  wire w5227;
  wire w5228;
  wire w5229;
  wire w5230;
  wire w5231;
  wire w5232;
  wire w5233;
  wire w5234;
  wire w5235;
  wire w5236;
  wire w5237;
  wire w5238;
  wire w5239;
  wire w5240;
  wire w5241;
  wire w5242;
  wire w5243;
  wire w5244;
  wire w5245;
  wire w5246;
  wire w5247;
  wire w5248;
  wire w5249;
  wire w5250;
  wire w5251;
  wire w5252;
  wire w5253;
  wire w5254;
  wire w5255;
  wire w5256;
  wire w5257;
  wire w5258;
  wire w5259;
  wire w5260;
  wire w5261;
  wire w5263;
  wire w5264;
  wire w5265;
  wire w5266;
  wire w5267;
  wire w5268;
  wire w5269;
  wire w5270;
  wire w5271;
  wire w5272;
  wire w5273;
  wire w5274;
  wire w5275;
  wire w5276;
  wire w5277;
  wire w5278;
  wire w5279;
  wire w5280;
  wire w5281;
  wire w5282;
  wire w5283;
  wire w5284;
  wire w5285;
  wire w5286;
  wire w5287;
  wire w5288;
  wire w5289;
  wire w5290;
  wire w5291;
  wire w5292;
  wire w5293;
  wire w5294;
  wire w5295;
  wire w5296;
  wire w5297;
  wire w5298;
  wire w5299;
  wire w5300;
  wire w5301;
  wire w5302;
  wire w5303;
  wire w5304;
  wire w5305;
  wire w5306;
  wire w5307;
  wire w5308;
  wire w5309;
  wire w5310;
  wire w5311;
  wire w5312;
  wire w5313;
  wire w5314;
  wire w5315;
  wire w5316;
  wire w5317;
  wire w5318;
  wire w5319;
  wire w5320;
  wire w5321;
  wire w5322;
  wire w5323;
  wire w5324;
  wire w5325;
  wire w5326;
  wire w5327;
  wire w5328;
  wire w5329;
  wire w5330;
  wire w5331;
  wire w5332;
  wire w5333;
  wire w5334;
  wire w5335;
  wire w5336;
  wire w5337;
  wire w5338;
  wire w5339;
  wire w5340;
  wire w5341;
  wire w5342;
  wire w5343;
  wire w5344;
  wire w5345;
  wire w5346;
  wire w5347;
  wire w5348;
  wire w5349;
  wire w5350;
  wire w5351;
  wire w5352;
  wire w5353;
  wire w5354;
  wire w5355;
  wire w5356;
  wire w5357;
  wire w5358;
  wire w5359;
  wire w5360;
  wire w5361;
  wire w5363;
  wire w5364;
  wire w5365;
  wire w5366;
  wire w5367;
  wire w5368;
  wire w5369;
  wire w5370;
  wire w5371;
  wire w5372;
  wire w5373;
  wire w5374;
  wire w5375;
  wire w5376;
  wire w5377;
  wire w5378;
  wire w5379;
  wire w5380;
  wire w5381;
  wire w5382;
  wire w5383;
  wire w5384;
  wire w5385;
  wire w5386;
  wire w5387;
  wire w5388;
  wire w5389;
  wire w5390;
  wire w5391;
  wire w5392;
  wire w5393;
  wire w5394;
  wire w5395;
  wire w5396;
  wire w5397;
  wire w5398;
  wire w5399;
  wire w5400;
  wire w5401;
  wire w5402;
  wire w5403;
  wire w5404;
  wire w5405;
  wire w5406;
  wire w5407;
  wire w5408;
  wire w5409;
  wire w5410;
  wire w5411;
  wire w5412;
  wire w5413;
  wire w5414;
  wire w5415;
  wire w5416;
  wire w5417;
  wire w5418;
  wire w5419;
  wire w5420;
  wire w5421;
  wire w5422;
  wire w5423;
  wire w5424;
  wire w5425;
  wire w5426;
  wire w5427;
  wire w5428;
  wire w5429;
  wire w5430;
  wire w5431;
  wire w5432;
  wire w5433;
  wire w5434;
  wire w5435;
  wire w5436;
  wire w5437;
  wire w5438;
  wire w5439;
  wire w5440;
  wire w5441;
  wire w5442;
  wire w5443;
  wire w5444;
  wire w5445;
  wire w5446;
  wire w5447;
  wire w5448;
  wire w5449;
  wire w5450;
  wire w5451;
  wire w5452;
  wire w5453;
  wire w5454;
  wire w5455;
  wire w5456;
  wire w5457;
  wire w5458;
  wire w5459;
  wire w5460;
  wire w5461;
  wire w5463;
  wire w5464;
  wire w5465;
  wire w5466;
  wire w5467;
  wire w5468;
  wire w5469;
  wire w5470;
  wire w5471;
  wire w5472;
  wire w5473;
  wire w5474;
  wire w5475;
  wire w5476;
  wire w5477;
  wire w5478;
  wire w5479;
  wire w5480;
  wire w5481;
  wire w5482;
  wire w5483;
  wire w5484;
  wire w5485;
  wire w5486;
  wire w5487;
  wire w5488;
  wire w5489;
  wire w5490;
  wire w5491;
  wire w5492;
  wire w5493;
  wire w5494;
  wire w5495;
  wire w5496;
  wire w5497;
  wire w5498;
  wire w5499;
  wire w5500;
  wire w5501;
  wire w5502;
  wire w5503;
  wire w5504;
  wire w5505;
  wire w5506;
  wire w5507;
  wire w5508;
  wire w5509;
  wire w5510;
  wire w5511;
  wire w5512;
  wire w5513;
  wire w5514;
  wire w5515;
  wire w5516;
  wire w5517;
  wire w5518;
  wire w5519;
  wire w5520;
  wire w5521;
  wire w5522;
  wire w5523;
  wire w5524;
  wire w5525;
  wire w5526;
  wire w5527;
  wire w5528;
  wire w5529;
  wire w5530;
  wire w5531;
  wire w5532;
  wire w5533;
  wire w5534;
  wire w5535;
  wire w5536;
  wire w5537;
  wire w5538;
  wire w5539;
  wire w5540;
  wire w5541;
  wire w5542;
  wire w5543;
  wire w5544;
  wire w5545;
  wire w5546;
  wire w5547;
  wire w5548;
  wire w5549;
  wire w5550;
  wire w5551;
  wire w5552;
  wire w5553;
  wire w5554;
  wire w5555;
  wire w5556;
  wire w5557;
  wire w5558;
  wire w5559;
  wire w5560;
  wire w5561;
  wire w5563;
  wire w5564;
  wire w5565;
  wire w5566;
  wire w5567;
  wire w5568;
  wire w5569;
  wire w5570;
  wire w5571;
  wire w5572;
  wire w5573;
  wire w5574;
  wire w5575;
  wire w5576;
  wire w5577;
  wire w5578;
  wire w5579;
  wire w5580;
  wire w5581;
  wire w5582;
  wire w5583;
  wire w5584;
  wire w5585;
  wire w5586;
  wire w5587;
  wire w5588;
  wire w5589;
  wire w5590;
  wire w5591;
  wire w5592;
  wire w5593;
  wire w5594;
  wire w5595;
  wire w5596;
  wire w5597;
  wire w5598;
  wire w5599;
  wire w5600;
  wire w5601;
  wire w5602;
  wire w5603;
  wire w5604;
  wire w5605;
  wire w5606;
  wire w5607;
  wire w5608;
  wire w5609;
  wire w5610;
  wire w5611;
  wire w5612;
  wire w5613;
  wire w5614;
  wire w5615;
  wire w5616;
  wire w5617;
  wire w5618;
  wire w5619;
  wire w5620;
  wire w5621;
  wire w5622;
  wire w5623;
  wire w5624;
  wire w5625;
  wire w5626;
  wire w5627;
  wire w5628;
  wire w5629;
  wire w5630;
  wire w5631;
  wire w5632;
  wire w5633;
  wire w5634;
  wire w5635;
  wire w5636;
  wire w5637;
  wire w5638;
  wire w5639;
  wire w5640;
  wire w5641;
  wire w5642;
  wire w5643;
  wire w5644;
  wire w5645;
  wire w5646;
  wire w5647;
  wire w5648;
  wire w5649;
  wire w5650;
  wire w5651;
  wire w5652;
  wire w5653;
  wire w5654;
  wire w5655;
  wire w5656;
  wire w5657;
  wire w5658;
  wire w5659;
  wire w5660;
  wire w5661;
  wire w5663;
  wire w5664;
  wire w5665;
  wire w5666;
  wire w5667;
  wire w5668;
  wire w5669;
  wire w5670;
  wire w5671;
  wire w5672;
  wire w5673;
  wire w5674;
  wire w5675;
  wire w5676;
  wire w5677;
  wire w5678;
  wire w5679;
  wire w5680;
  wire w5681;
  wire w5682;
  wire w5683;
  wire w5684;
  wire w5685;
  wire w5686;
  wire w5687;
  wire w5688;
  wire w5689;
  wire w5690;
  wire w5691;
  wire w5692;
  wire w5693;
  wire w5694;
  wire w5695;
  wire w5696;
  wire w5697;
  wire w5698;
  wire w5699;
  wire w5700;
  wire w5701;
  wire w5702;
  wire w5703;
  wire w5704;
  wire w5705;
  wire w5706;
  wire w5707;
  wire w5708;
  wire w5709;
  wire w5710;
  wire w5711;
  wire w5712;
  wire w5713;
  wire w5714;
  wire w5715;
  wire w5716;
  wire w5717;
  wire w5718;
  wire w5719;
  wire w5720;
  wire w5721;
  wire w5722;
  wire w5723;
  wire w5724;
  wire w5725;
  wire w5726;
  wire w5727;
  wire w5728;
  wire w5729;
  wire w5730;
  wire w5731;
  wire w5732;
  wire w5733;
  wire w5734;
  wire w5735;
  wire w5736;
  wire w5737;
  wire w5738;
  wire w5739;
  wire w5740;
  wire w5741;
  wire w5742;
  wire w5743;
  wire w5744;
  wire w5745;
  wire w5746;
  wire w5747;
  wire w5748;
  wire w5749;
  wire w5750;
  wire w5751;
  wire w5752;
  wire w5753;
  wire w5754;
  wire w5755;
  wire w5756;
  wire w5757;
  wire w5758;
  wire w5759;
  wire w5760;
  wire w5761;
  wire w5763;
  wire w5764;
  wire w5765;
  wire w5766;
  wire w5767;
  wire w5768;
  wire w5769;
  wire w5770;
  wire w5771;
  wire w5772;
  wire w5773;
  wire w5774;
  wire w5775;
  wire w5776;
  wire w5777;
  wire w5778;
  wire w5779;
  wire w5780;
  wire w5781;
  wire w5782;
  wire w5783;
  wire w5784;
  wire w5785;
  wire w5786;
  wire w5787;
  wire w5788;
  wire w5789;
  wire w5790;
  wire w5791;
  wire w5792;
  wire w5793;
  wire w5794;
  wire w5795;
  wire w5796;
  wire w5797;
  wire w5798;
  wire w5799;
  wire w5800;
  wire w5801;
  wire w5802;
  wire w5803;
  wire w5804;
  wire w5805;
  wire w5806;
  wire w5807;
  wire w5808;
  wire w5809;
  wire w5810;
  wire w5811;
  wire w5812;
  wire w5813;
  wire w5814;
  wire w5815;
  wire w5816;
  wire w5817;
  wire w5818;
  wire w5819;
  wire w5820;
  wire w5821;
  wire w5822;
  wire w5823;
  wire w5824;
  wire w5825;
  wire w5826;
  wire w5827;
  wire w5828;
  wire w5829;
  wire w5830;
  wire w5831;
  wire w5832;
  wire w5833;
  wire w5834;
  wire w5835;
  wire w5836;
  wire w5837;
  wire w5838;
  wire w5839;
  wire w5840;
  wire w5841;
  wire w5842;
  wire w5843;
  wire w5844;
  wire w5845;
  wire w5846;
  wire w5847;
  wire w5848;
  wire w5849;
  wire w5850;
  wire w5851;
  wire w5852;
  wire w5853;
  wire w5854;
  wire w5855;
  wire w5856;
  wire w5857;
  wire w5858;
  wire w5859;
  wire w5860;
  wire w5861;
  wire w5863;
  wire w5864;
  wire w5865;
  wire w5866;
  wire w5867;
  wire w5868;
  wire w5869;
  wire w5870;
  wire w5871;
  wire w5872;
  wire w5873;
  wire w5874;
  wire w5875;
  wire w5876;
  wire w5877;
  wire w5878;
  wire w5879;
  wire w5880;
  wire w5881;
  wire w5882;
  wire w5883;
  wire w5884;
  wire w5885;
  wire w5886;
  wire w5887;
  wire w5888;
  wire w5889;
  wire w5890;
  wire w5891;
  wire w5892;
  wire w5893;
  wire w5894;
  wire w5895;
  wire w5896;
  wire w5897;
  wire w5898;
  wire w5899;
  wire w5900;
  wire w5901;
  wire w5902;
  wire w5903;
  wire w5904;
  wire w5905;
  wire w5906;
  wire w5907;
  wire w5908;
  wire w5909;
  wire w5910;
  wire w5911;
  wire w5912;
  wire w5913;
  wire w5914;
  wire w5915;
  wire w5916;
  wire w5917;
  wire w5918;
  wire w5919;
  wire w5920;
  wire w5921;
  wire w5922;
  wire w5923;
  wire w5924;
  wire w5925;
  wire w5926;
  wire w5927;
  wire w5928;
  wire w5929;
  wire w5930;
  wire w5931;
  wire w5932;
  wire w5933;
  wire w5934;
  wire w5935;
  wire w5936;
  wire w5937;
  wire w5938;
  wire w5939;
  wire w5940;
  wire w5941;
  wire w5942;
  wire w5943;
  wire w5944;
  wire w5945;
  wire w5946;
  wire w5947;
  wire w5948;
  wire w5949;
  wire w5950;
  wire w5951;
  wire w5952;
  wire w5953;
  wire w5954;
  wire w5955;
  wire w5956;
  wire w5957;
  wire w5958;
  wire w5959;
  wire w5960;
  wire w5961;
  wire w5963;
  wire w5964;
  wire w5965;
  wire w5966;
  wire w5967;
  wire w5968;
  wire w5969;
  wire w5970;
  wire w5971;
  wire w5972;
  wire w5973;
  wire w5974;
  wire w5975;
  wire w5976;
  wire w5977;
  wire w5978;
  wire w5979;
  wire w5980;
  wire w5981;
  wire w5982;
  wire w5983;
  wire w5984;
  wire w5985;
  wire w5986;
  wire w5987;
  wire w5988;
  wire w5989;
  wire w5990;
  wire w5991;
  wire w5992;
  wire w5993;
  wire w5994;
  wire w5995;
  wire w5996;
  wire w5997;
  wire w5998;
  wire w5999;
  wire w6000;
  wire w6001;
  wire w6002;
  wire w6003;
  wire w6004;
  wire w6005;
  wire w6006;
  wire w6007;
  wire w6008;
  wire w6009;
  wire w6010;
  wire w6011;
  wire w6012;
  wire w6013;
  wire w6014;
  wire w6015;
  wire w6016;
  wire w6017;
  wire w6018;
  wire w6019;
  wire w6020;
  wire w6021;
  wire w6022;
  wire w6023;
  wire w6024;
  wire w6025;
  wire w6026;
  wire w6027;
  wire w6028;
  wire w6029;
  wire w6030;
  wire w6031;
  wire w6032;
  wire w6033;
  wire w6034;
  wire w6035;
  wire w6036;
  wire w6037;
  wire w6038;
  wire w6039;
  wire w6040;
  wire w6041;
  wire w6042;
  wire w6043;
  wire w6044;
  wire w6045;
  wire w6046;
  wire w6047;
  wire w6048;
  wire w6049;
  wire w6050;
  wire w6051;
  wire w6052;
  wire w6053;
  wire w6054;
  wire w6055;
  wire w6056;
  wire w6057;
  wire w6058;
  wire w6059;
  wire w6060;
  wire w6061;
  wire w6063;
  wire w6064;
  wire w6065;
  wire w6066;
  wire w6067;
  wire w6068;
  wire w6069;
  wire w6070;
  wire w6071;
  wire w6072;
  wire w6073;
  wire w6074;
  wire w6075;
  wire w6076;
  wire w6077;
  wire w6078;
  wire w6079;
  wire w6080;
  wire w6081;
  wire w6082;
  wire w6083;
  wire w6084;
  wire w6085;
  wire w6086;
  wire w6087;
  wire w6088;
  wire w6089;
  wire w6090;
  wire w6091;
  wire w6092;
  wire w6093;
  wire w6094;
  wire w6095;
  wire w6096;
  wire w6097;
  wire w6098;
  wire w6099;
  wire w6100;
  wire w6101;
  wire w6102;
  wire w6103;
  wire w6104;
  wire w6105;
  wire w6106;
  wire w6107;
  wire w6108;
  wire w6109;
  wire w6110;
  wire w6111;
  wire w6112;
  wire w6113;
  wire w6114;
  wire w6115;
  wire w6116;
  wire w6117;
  wire w6118;
  wire w6119;
  wire w6120;
  wire w6121;
  wire w6122;
  wire w6123;
  wire w6124;
  wire w6125;
  wire w6126;
  wire w6127;
  wire w6128;
  wire w6129;
  wire w6130;
  wire w6131;
  wire w6132;
  wire w6133;
  wire w6134;
  wire w6135;
  wire w6136;
  wire w6137;
  wire w6138;
  wire w6139;
  wire w6140;
  wire w6141;
  wire w6142;
  wire w6143;
  wire w6144;
  wire w6145;
  wire w6146;
  wire w6147;
  wire w6148;
  wire w6149;
  wire w6150;
  wire w6151;
  wire w6152;
  wire w6153;
  wire w6154;
  wire w6155;
  wire w6156;
  wire w6157;
  wire w6158;
  wire w6159;
  wire w6160;
  wire w6161;
  wire w6163;
  wire w6164;
  wire w6165;
  wire w6166;
  wire w6167;
  wire w6168;
  wire w6169;
  wire w6170;
  wire w6171;
  wire w6172;
  wire w6173;
  wire w6174;
  wire w6175;
  wire w6176;
  wire w6177;
  wire w6178;
  wire w6179;
  wire w6180;
  wire w6181;
  wire w6182;
  wire w6183;
  wire w6184;
  wire w6185;
  wire w6186;
  wire w6187;
  wire w6188;
  wire w6189;
  wire w6190;
  wire w6191;
  wire w6192;
  wire w6193;
  wire w6194;
  wire w6195;
  wire w6196;
  wire w6197;
  wire w6198;
  wire w6199;
  wire w6200;
  wire w6201;
  wire w6202;
  wire w6203;
  wire w6204;
  wire w6205;
  wire w6206;
  wire w6207;
  wire w6208;
  wire w6209;
  wire w6210;
  wire w6211;
  wire w6212;
  wire w6213;
  wire w6214;
  wire w6215;
  wire w6216;
  wire w6217;
  wire w6218;
  wire w6219;
  wire w6220;
  wire w6221;
  wire w6222;
  wire w6223;
  wire w6224;
  wire w6225;
  wire w6226;
  wire w6227;
  wire w6228;
  wire w6229;
  wire w6230;
  wire w6231;
  wire w6232;
  wire w6233;
  wire w6234;
  wire w6235;
  wire w6236;
  wire w6237;
  wire w6238;
  wire w6239;
  wire w6240;
  wire w6241;
  wire w6242;
  wire w6243;
  wire w6244;
  wire w6245;
  wire w6246;
  wire w6247;
  wire w6248;
  wire w6249;
  wire w6250;
  wire w6251;
  wire w6252;
  wire w6253;
  wire w6254;
  wire w6255;
  wire w6256;
  wire w6257;
  wire w6258;
  wire w6259;
  wire w6260;
  wire w6261;
  wire w6263;
  wire w6264;
  wire w6265;
  wire w6266;
  wire w6267;
  wire w6268;
  wire w6269;
  wire w6270;
  wire w6271;
  wire w6272;
  wire w6273;
  wire w6274;
  wire w6275;
  wire w6276;
  wire w6277;
  wire w6278;
  wire w6279;
  wire w6280;
  wire w6281;
  wire w6282;
  wire w6283;
  wire w6284;
  wire w6285;
  wire w6286;
  wire w6287;
  wire w6288;
  wire w6289;
  wire w6290;
  wire w6291;
  wire w6292;
  wire w6293;
  wire w6294;
  wire w6295;
  wire w6296;
  wire w6297;
  wire w6298;
  wire w6299;
  wire w6300;
  wire w6301;
  wire w6302;
  wire w6303;
  wire w6304;
  wire w6305;
  wire w6306;
  wire w6307;
  wire w6308;
  wire w6309;
  wire w6310;
  wire w6311;
  wire w6312;
  wire w6313;
  wire w6314;
  wire w6315;
  wire w6316;
  wire w6317;
  wire w6318;
  wire w6319;
  wire w6320;
  wire w6321;
  wire w6322;
  wire w6323;
  wire w6324;
  wire w6325;
  wire w6326;
  wire w6327;
  wire w6328;
  wire w6329;
  wire w6330;
  wire w6331;
  wire w6332;
  wire w6333;
  wire w6334;
  wire w6335;
  wire w6336;
  wire w6337;
  wire w6338;
  wire w6339;
  wire w6340;
  wire w6341;
  wire w6342;
  wire w6343;
  wire w6344;
  wire w6345;
  wire w6346;
  wire w6347;
  wire w6348;
  wire w6349;
  wire w6350;
  wire w6351;
  wire w6352;
  wire w6353;
  wire w6354;
  wire w6355;
  wire w6356;
  wire w6357;
  wire w6358;
  wire w6359;
  wire w6360;
  wire w6361;
  wire w6363;
  wire w6364;
  wire w6365;
  wire w6366;
  wire w6367;
  wire w6368;
  wire w6369;
  wire w6370;
  wire w6371;
  wire w6372;
  wire w6373;
  wire w6374;
  wire w6375;
  wire w6376;
  wire w6377;
  wire w6378;
  wire w6379;
  wire w6380;
  wire w6381;
  wire w6382;
  wire w6383;
  wire w6384;
  wire w6385;
  wire w6386;
  wire w6387;
  wire w6388;
  wire w6389;
  wire w6390;
  wire w6391;
  wire w6392;
  wire w6393;
  wire w6394;
  wire w6395;
  wire w6396;
  wire w6397;
  wire w6398;
  wire w6399;
  wire w6400;
  wire w6401;
  wire w6402;
  wire w6403;
  wire w6404;
  wire w6405;
  wire w6406;
  wire w6407;
  wire w6408;
  wire w6409;
  wire w6410;
  wire w6411;
  wire w6412;
  wire w6413;
  wire w6414;
  wire w6415;
  wire w6416;
  wire w6417;
  wire w6418;
  wire w6419;
  wire w6420;
  wire w6421;
  wire w6422;
  wire w6423;
  wire w6424;
  wire w6425;
  wire w6426;
  wire w6427;
  wire w6428;
  wire w6429;
  wire w6430;
  wire w6431;
  wire w6432;
  wire w6433;
  wire w6434;
  wire w6435;
  wire w6436;
  wire w6437;
  wire w6438;
  wire w6439;
  wire w6440;
  wire w6441;
  wire w6442;
  wire w6443;
  wire w6444;
  wire w6445;
  wire w6446;
  wire w6447;
  wire w6448;
  wire w6449;
  wire w6450;
  wire w6451;
  wire w6452;
  wire w6453;
  wire w6454;
  wire w6455;
  wire w6456;
  wire w6457;
  wire w6458;
  wire w6459;
  wire w6460;
  wire w6461;
  wire w6463;
  wire w6464;
  wire w6465;
  wire w6466;
  wire w6467;
  wire w6468;
  wire w6469;
  wire w6470;
  wire w6471;
  wire w6472;
  wire w6473;
  wire w6474;
  wire w6475;
  wire w6476;
  wire w6477;
  wire w6478;
  wire w6479;
  wire w6480;
  wire w6481;
  wire w6482;
  wire w6483;
  wire w6484;
  wire w6485;
  wire w6486;
  wire w6487;
  wire w6488;
  wire w6489;
  wire w6490;
  wire w6491;
  wire w6492;
  wire w6493;
  wire w6494;
  wire w6495;
  wire w6496;
  wire w6497;
  wire w6498;
  wire w6499;
  wire w6500;
  wire w6501;
  wire w6502;
  wire w6503;
  wire w6504;
  wire w6505;
  wire w6506;
  wire w6507;
  wire w6508;
  wire w6509;
  wire w6510;
  wire w6511;
  wire w6512;
  wire w6513;
  wire w6514;
  wire w6515;
  wire w6516;
  wire w6517;
  wire w6518;
  wire w6519;
  wire w6520;
  wire w6521;
  wire w6522;
  wire w6523;
  wire w6524;
  wire w6525;
  wire w6526;
  wire w6527;
  wire w6528;
  wire w6529;
  wire w6530;
  wire w6531;
  wire w6532;
  wire w6533;
  wire w6534;
  wire w6535;
  wire w6536;
  wire w6537;
  wire w6538;
  wire w6539;
  wire w6540;
  wire w6541;
  wire w6542;
  wire w6543;
  wire w6544;
  wire w6545;
  wire w6546;
  wire w6547;
  wire w6548;
  wire w6549;
  wire w6550;
  wire w6551;
  wire w6552;
  wire w6553;
  wire w6554;
  wire w6555;
  wire w6556;
  wire w6557;
  wire w6558;
  wire w6559;
  wire w6560;
  wire w6561;
  wire w6563;
  wire w6564;
  wire w6565;
  wire w6566;
  wire w6567;
  wire w6568;
  wire w6569;
  wire w6570;
  wire w6571;
  wire w6572;
  wire w6573;
  wire w6574;
  wire w6575;
  wire w6576;
  wire w6577;
  wire w6578;
  wire w6579;
  wire w6580;
  wire w6581;
  wire w6582;
  wire w6583;
  wire w6584;
  wire w6585;
  wire w6586;
  wire w6587;
  wire w6588;
  wire w6589;
  wire w6590;
  wire w6591;
  wire w6592;
  wire w6593;
  wire w6594;
  wire w6595;
  wire w6596;
  wire w6597;
  wire w6598;
  wire w6599;
  wire w6600;
  wire w6601;
  wire w6602;
  wire w6603;
  wire w6604;
  wire w6605;
  wire w6606;
  wire w6607;
  wire w6608;
  wire w6609;
  wire w6610;
  wire w6611;
  wire w6612;
  wire w6613;
  wire w6614;
  wire w6615;
  wire w6616;
  wire w6617;
  wire w6618;
  wire w6619;
  wire w6620;
  wire w6621;
  wire w6622;
  wire w6623;
  wire w6624;
  wire w6625;
  wire w6626;
  wire w6627;
  wire w6628;
  wire w6629;
  wire w6630;
  wire w6631;
  wire w6632;
  wire w6633;
  wire w6634;
  wire w6635;
  wire w6636;
  wire w6637;
  wire w6638;
  wire w6639;
  wire w6640;
  wire w6641;
  wire w6642;
  wire w6643;
  wire w6644;
  wire w6645;
  wire w6646;
  wire w6647;
  wire w6648;
  wire w6649;
  wire w6650;
  wire w6651;
  wire w6652;
  wire w6653;
  wire w6654;
  wire w6655;
  wire w6656;
  wire w6657;
  wire w6658;
  wire w6659;
  wire w6660;
  wire w6661;
  wire w6663;
  wire w6664;
  wire w6665;
  wire w6666;
  wire w6667;
  wire w6668;
  wire w6669;
  wire w6670;
  wire w6671;
  wire w6672;
  wire w6673;
  wire w6674;
  wire w6675;
  wire w6676;
  wire w6677;
  wire w6678;
  wire w6679;
  wire w6680;
  wire w6681;
  wire w6682;
  wire w6683;
  wire w6684;
  wire w6685;
  wire w6686;
  wire w6687;
  wire w6688;
  wire w6689;
  wire w6690;
  wire w6691;
  wire w6692;
  wire w6693;
  wire w6694;
  wire w6695;
  wire w6696;
  wire w6697;
  wire w6698;
  wire w6699;
  wire w6700;
  wire w6701;
  wire w6702;
  wire w6703;
  wire w6704;
  wire w6705;
  wire w6706;
  wire w6707;
  wire w6708;
  wire w6709;
  wire w6710;
  wire w6711;
  wire w6712;
  wire w6713;
  wire w6714;
  wire w6715;
  wire w6716;
  wire w6717;
  wire w6718;
  wire w6719;
  wire w6720;
  wire w6721;
  wire w6722;
  wire w6723;
  wire w6724;
  wire w6725;
  wire w6726;
  wire w6727;
  wire w6728;
  wire w6729;
  wire w6730;
  wire w6731;
  wire w6732;
  wire w6733;
  wire w6734;
  wire w6735;
  wire w6736;
  wire w6737;
  wire w6738;
  wire w6739;
  wire w6740;
  wire w6741;
  wire w6742;
  wire w6743;
  wire w6744;
  wire w6745;
  wire w6746;
  wire w6747;
  wire w6748;
  wire w6749;
  wire w6750;
  wire w6751;
  wire w6752;
  wire w6753;
  wire w6754;
  wire w6755;
  wire w6756;
  wire w6757;
  wire w6758;
  wire w6759;
  wire w6760;
  wire w6761;
  wire w6763;
  wire w6764;
  wire w6765;
  wire w6766;
  wire w6767;
  wire w6768;
  wire w6769;
  wire w6770;
  wire w6771;
  wire w6772;
  wire w6773;
  wire w6774;
  wire w6775;
  wire w6776;
  wire w6777;
  wire w6778;
  wire w6779;
  wire w6780;
  wire w6781;
  wire w6782;
  wire w6783;
  wire w6784;
  wire w6785;
  wire w6786;
  wire w6787;
  wire w6788;
  wire w6789;
  wire w6790;
  wire w6791;
  wire w6792;
  wire w6793;
  wire w6794;
  wire w6795;
  wire w6796;
  wire w6797;
  wire w6798;
  wire w6799;
  wire w6800;
  wire w6801;
  wire w6802;
  wire w6803;
  wire w6804;
  wire w6805;
  wire w6806;
  wire w6807;
  wire w6808;
  wire w6809;
  wire w6810;
  wire w6811;
  wire w6812;
  wire w6813;
  wire w6814;
  wire w6815;
  wire w6816;
  wire w6817;
  wire w6818;
  wire w6819;
  wire w6820;
  wire w6821;
  wire w6822;
  wire w6823;
  wire w6824;
  wire w6825;
  wire w6826;
  wire w6827;
  wire w6828;
  wire w6829;
  wire w6830;
  wire w6831;
  wire w6832;
  wire w6833;
  wire w6834;
  wire w6835;
  wire w6836;
  wire w6837;
  wire w6838;
  wire w6839;
  wire w6840;
  wire w6841;
  wire w6842;
  wire w6843;
  wire w6844;
  wire w6845;
  wire w6846;
  wire w6847;
  wire w6848;
  wire w6849;
  wire w6850;
  wire w6851;
  wire w6852;
  wire w6853;
  wire w6854;
  wire w6855;
  wire w6856;
  wire w6857;
  wire w6858;
  wire w6859;
  wire w6860;
  wire w6861;
  wire w6863;
  wire w6864;
  wire w6865;
  wire w6866;
  wire w6867;
  wire w6868;
  wire w6869;
  wire w6870;
  wire w6871;
  wire w6872;
  wire w6873;
  wire w6874;
  wire w6875;
  wire w6876;
  wire w6877;
  wire w6878;
  wire w6879;
  wire w6880;
  wire w6881;
  wire w6882;
  wire w6883;
  wire w6884;
  wire w6885;
  wire w6886;
  wire w6887;
  wire w6888;
  wire w6889;
  wire w6890;
  wire w6891;
  wire w6892;
  wire w6893;
  wire w6894;
  wire w6895;
  wire w6896;
  wire w6897;
  wire w6898;
  wire w6899;
  wire w6900;
  wire w6901;
  wire w6902;
  wire w6903;
  wire w6904;
  wire w6905;
  wire w6906;
  wire w6907;
  wire w6908;
  wire w6909;
  wire w6910;
  wire w6911;
  wire w6912;
  wire w6913;
  wire w6914;
  wire w6915;
  wire w6916;
  wire w6917;
  wire w6918;
  wire w6919;
  wire w6920;
  wire w6921;
  wire w6922;
  wire w6923;
  wire w6924;
  wire w6925;
  wire w6926;
  wire w6927;
  wire w6928;
  wire w6929;
  wire w6930;
  wire w6931;
  wire w6932;
  wire w6933;
  wire w6934;
  wire w6935;
  wire w6936;
  wire w6937;
  wire w6938;
  wire w6939;
  wire w6940;
  wire w6941;
  wire w6942;
  wire w6943;
  wire w6944;
  wire w6945;
  wire w6946;
  wire w6947;
  wire w6948;
  wire w6949;
  wire w6950;
  wire w6951;
  wire w6952;
  wire w6953;
  wire w6954;
  wire w6955;
  wire w6956;
  wire w6957;
  wire w6958;
  wire w6959;
  wire w6960;
  wire w6961;
  wire w6963;
  wire w6964;
  wire w6965;
  wire w6966;
  wire w6967;
  wire w6968;
  wire w6969;
  wire w6970;
  wire w6971;
  wire w6972;
  wire w6973;
  wire w6974;
  wire w6975;
  wire w6976;
  wire w6977;
  wire w6978;
  wire w6979;
  wire w6980;
  wire w6981;
  wire w6982;
  wire w6983;
  wire w6984;
  wire w6985;
  wire w6986;
  wire w6987;
  wire w6988;
  wire w6989;
  wire w6990;
  wire w6991;
  wire w6992;
  wire w6993;
  wire w6994;
  wire w6995;
  wire w6996;
  wire w6997;
  wire w6998;
  wire w6999;
  wire w7000;
  wire w7001;
  wire w7002;
  wire w7003;
  wire w7004;
  wire w7005;
  wire w7006;
  wire w7007;
  wire w7008;
  wire w7009;
  wire w7010;
  wire w7011;
  wire w7012;
  wire w7013;
  wire w7014;
  wire w7015;
  wire w7016;
  wire w7017;
  wire w7018;
  wire w7019;
  wire w7020;
  wire w7021;
  wire w7022;
  wire w7023;
  wire w7024;
  wire w7025;
  wire w7026;
  wire w7027;
  wire w7028;
  wire w7029;
  wire w7030;
  wire w7031;
  wire w7032;
  wire w7033;
  wire w7034;
  wire w7035;
  wire w7036;
  wire w7037;
  wire w7038;
  wire w7039;
  wire w7040;
  wire w7041;
  wire w7042;
  wire w7043;
  wire w7044;
  wire w7045;
  wire w7046;
  wire w7047;
  wire w7048;
  wire w7049;
  wire w7050;
  wire w7051;
  wire w7052;
  wire w7053;
  wire w7054;
  wire w7055;
  wire w7056;
  wire w7057;
  wire w7058;
  wire w7059;
  wire w7060;
  wire w7061;
  wire w7063;
  wire w7064;
  wire w7065;
  wire w7066;
  wire w7067;
  wire w7068;
  wire w7069;
  wire w7070;
  wire w7071;
  wire w7072;
  wire w7073;
  wire w7074;
  wire w7075;
  wire w7076;
  wire w7077;
  wire w7078;
  wire w7079;
  wire w7080;
  wire w7081;
  wire w7082;
  wire w7083;
  wire w7084;
  wire w7085;
  wire w7086;
  wire w7087;
  wire w7088;
  wire w7089;
  wire w7090;
  wire w7091;
  wire w7092;
  wire w7093;
  wire w7094;
  wire w7095;
  wire w7096;
  wire w7097;
  wire w7098;
  wire w7099;
  wire w7100;
  wire w7101;
  wire w7102;
  wire w7103;
  wire w7104;
  wire w7105;
  wire w7106;
  wire w7107;
  wire w7108;
  wire w7109;
  wire w7110;
  wire w7111;
  wire w7112;
  wire w7113;
  wire w7114;
  wire w7115;
  wire w7116;
  wire w7117;
  wire w7118;
  wire w7119;
  wire w7120;
  wire w7121;
  wire w7122;
  wire w7123;
  wire w7124;
  wire w7125;
  wire w7126;
  wire w7127;
  wire w7128;
  wire w7129;
  wire w7130;
  wire w7131;
  wire w7132;
  wire w7133;
  wire w7134;
  wire w7135;
  wire w7136;
  wire w7137;
  wire w7138;
  wire w7139;
  wire w7140;
  wire w7141;
  wire w7142;
  wire w7143;
  wire w7144;
  wire w7145;
  wire w7146;
  wire w7147;
  wire w7148;
  wire w7149;
  wire w7150;
  wire w7151;
  wire w7152;
  wire w7153;
  wire w7154;
  wire w7155;
  wire w7156;
  wire w7157;
  wire w7158;
  wire w7159;
  wire w7160;
  wire w7161;
  wire w7163;
  wire w7164;
  wire w7165;
  wire w7166;
  wire w7167;
  wire w7168;
  wire w7169;
  wire w7170;
  wire w7171;
  wire w7172;
  wire w7173;
  wire w7174;
  wire w7175;
  wire w7176;
  wire w7177;
  wire w7178;
  wire w7179;
  wire w7180;
  wire w7181;
  wire w7182;
  wire w7183;
  wire w7184;
  wire w7185;
  wire w7186;
  wire w7187;
  wire w7188;
  wire w7189;
  wire w7190;
  wire w7191;
  wire w7192;
  wire w7193;
  wire w7194;
  wire w7195;
  wire w7196;
  wire w7197;
  wire w7198;
  wire w7199;
  wire w7200;
  wire w7201;
  wire w7202;
  wire w7203;
  wire w7204;
  wire w7205;
  wire w7206;
  wire w7207;
  wire w7208;
  wire w7209;
  wire w7210;
  wire w7211;
  wire w7212;
  wire w7213;
  wire w7214;
  wire w7215;
  wire w7216;
  wire w7217;
  wire w7218;
  wire w7219;
  wire w7220;
  wire w7221;
  wire w7222;
  wire w7223;
  wire w7224;
  wire w7225;
  wire w7226;
  wire w7227;
  wire w7228;
  wire w7229;
  wire w7230;
  wire w7231;
  wire w7232;
  wire w7233;
  wire w7234;
  wire w7235;
  wire w7236;
  wire w7237;
  wire w7238;
  wire w7239;
  wire w7240;
  wire w7241;
  wire w7242;
  wire w7243;
  wire w7244;
  wire w7245;
  wire w7246;
  wire w7247;
  wire w7248;
  wire w7249;
  wire w7250;
  wire w7251;
  wire w7252;
  wire w7253;
  wire w7254;
  wire w7255;
  wire w7256;
  wire w7257;
  wire w7258;
  wire w7259;
  wire w7260;
  wire w7261;
  wire w7263;
  wire w7264;
  wire w7265;
  wire w7266;
  wire w7267;
  wire w7268;
  wire w7269;
  wire w7270;
  wire w7271;
  wire w7272;
  wire w7273;
  wire w7274;
  wire w7275;
  wire w7276;
  wire w7277;
  wire w7278;
  wire w7279;
  wire w7280;
  wire w7281;
  wire w7282;
  wire w7283;
  wire w7284;
  wire w7285;
  wire w7286;
  wire w7287;
  wire w7288;
  wire w7289;
  wire w7290;
  wire w7291;
  wire w7292;
  wire w7293;
  wire w7294;
  wire w7295;
  wire w7296;
  wire w7297;
  wire w7298;
  wire w7299;
  wire w7300;
  wire w7301;
  wire w7302;
  wire w7303;
  wire w7304;
  wire w7305;
  wire w7306;
  wire w7307;
  wire w7308;
  wire w7309;
  wire w7310;
  wire w7311;
  wire w7312;
  wire w7313;
  wire w7314;
  wire w7315;
  wire w7316;
  wire w7317;
  wire w7318;
  wire w7319;
  wire w7320;
  wire w7321;
  wire w7322;
  wire w7323;
  wire w7324;
  wire w7325;
  wire w7326;
  wire w7327;
  wire w7328;
  wire w7329;
  wire w7330;
  wire w7331;
  wire w7332;
  wire w7333;
  wire w7334;
  wire w7335;
  wire w7336;
  wire w7337;
  wire w7338;
  wire w7339;
  wire w7340;
  wire w7341;
  wire w7342;
  wire w7343;
  wire w7344;
  wire w7345;
  wire w7346;
  wire w7347;
  wire w7348;
  wire w7349;
  wire w7350;
  wire w7351;
  wire w7352;
  wire w7353;
  wire w7354;
  wire w7355;
  wire w7356;
  wire w7357;
  wire w7358;
  wire w7359;
  wire w7360;
  wire w7361;
  wire w7363;
  wire w7364;
  wire w7365;
  wire w7366;
  wire w7367;
  wire w7368;
  wire w7369;
  wire w7370;
  wire w7371;
  wire w7372;
  wire w7373;
  wire w7374;
  wire w7375;
  wire w7376;
  wire w7377;
  wire w7378;
  wire w7379;
  wire w7380;
  wire w7381;
  wire w7382;
  wire w7383;
  wire w7384;
  wire w7385;
  wire w7386;
  wire w7387;
  wire w7388;
  wire w7389;
  wire w7390;
  wire w7391;
  wire w7392;
  wire w7393;
  wire w7394;
  wire w7395;
  wire w7396;
  wire w7397;
  wire w7398;
  wire w7399;
  wire w7400;
  wire w7401;
  wire w7402;
  wire w7403;
  wire w7404;
  wire w7405;
  wire w7406;
  wire w7407;
  wire w7408;
  wire w7409;
  wire w7410;
  wire w7411;
  wire w7412;
  wire w7413;
  wire w7414;
  wire w7415;
  wire w7416;
  wire w7417;
  wire w7418;
  wire w7419;
  wire w7420;
  wire w7421;
  wire w7422;
  wire w7423;
  wire w7424;
  wire w7425;
  wire w7426;
  wire w7427;
  wire w7428;
  wire w7429;
  wire w7430;
  wire w7431;
  wire w7432;
  wire w7433;
  wire w7434;
  wire w7435;
  wire w7436;
  wire w7437;
  wire w7438;
  wire w7439;
  wire w7440;
  wire w7441;
  wire w7442;
  wire w7443;
  wire w7444;
  wire w7445;
  wire w7446;
  wire w7447;
  wire w7448;
  wire w7449;
  wire w7450;
  wire w7451;
  wire w7452;
  wire w7453;
  wire w7454;
  wire w7455;
  wire w7456;
  wire w7457;
  wire w7458;
  wire w7459;
  wire w7460;
  wire w7461;
  wire w7463;
  wire w7464;
  wire w7465;
  wire w7466;
  wire w7467;
  wire w7468;
  wire w7469;
  wire w7470;
  wire w7471;
  wire w7472;
  wire w7473;
  wire w7474;
  wire w7475;
  wire w7476;
  wire w7477;
  wire w7478;
  wire w7479;
  wire w7480;
  wire w7481;
  wire w7482;
  wire w7483;
  wire w7484;
  wire w7485;
  wire w7486;
  wire w7487;
  wire w7488;
  wire w7489;
  wire w7490;
  wire w7491;
  wire w7492;
  wire w7493;
  wire w7494;
  wire w7495;
  wire w7496;
  wire w7497;
  wire w7498;
  wire w7499;
  wire w7500;
  wire w7501;
  wire w7502;
  wire w7503;
  wire w7504;
  wire w7505;
  wire w7506;
  wire w7507;
  wire w7508;
  wire w7509;
  wire w7510;
  wire w7511;
  wire w7512;
  wire w7513;
  wire w7514;
  wire w7515;
  wire w7516;
  wire w7517;
  wire w7518;
  wire w7519;
  wire w7520;
  wire w7521;
  wire w7522;
  wire w7523;
  wire w7524;
  wire w7525;
  wire w7526;
  wire w7527;
  wire w7528;
  wire w7529;
  wire w7530;
  wire w7531;
  wire w7532;
  wire w7533;
  wire w7534;
  wire w7535;
  wire w7536;
  wire w7537;
  wire w7538;
  wire w7539;
  wire w7540;
  wire w7541;
  wire w7542;
  wire w7543;
  wire w7544;
  wire w7545;
  wire w7546;
  wire w7547;
  wire w7548;
  wire w7549;
  wire w7550;
  wire w7551;
  wire w7552;
  wire w7553;
  wire w7554;
  wire w7555;
  wire w7556;
  wire w7557;
  wire w7558;
  wire w7559;
  wire w7560;
  wire w7561;
  wire w7563;
  wire w7564;
  wire w7565;
  wire w7566;
  wire w7567;
  wire w7568;
  wire w7569;
  wire w7570;
  wire w7571;
  wire w7572;
  wire w7573;
  wire w7574;
  wire w7575;
  wire w7576;
  wire w7577;
  wire w7578;
  wire w7579;
  wire w7580;
  wire w7581;
  wire w7582;
  wire w7583;
  wire w7584;
  wire w7585;
  wire w7586;
  wire w7587;
  wire w7588;
  wire w7589;
  wire w7590;
  wire w7591;
  wire w7592;
  wire w7593;
  wire w7594;
  wire w7595;
  wire w7596;
  wire w7597;
  wire w7598;
  wire w7599;
  wire w7600;
  wire w7601;
  wire w7602;
  wire w7603;
  wire w7604;
  wire w7605;
  wire w7606;
  wire w7607;
  wire w7608;
  wire w7609;
  wire w7610;
  wire w7611;
  wire w7612;
  wire w7613;
  wire w7614;
  wire w7615;
  wire w7616;
  wire w7617;
  wire w7618;
  wire w7619;
  wire w7620;
  wire w7621;
  wire w7622;
  wire w7623;
  wire w7624;
  wire w7625;
  wire w7626;
  wire w7627;
  wire w7628;
  wire w7629;
  wire w7630;
  wire w7631;
  wire w7632;
  wire w7633;
  wire w7634;
  wire w7635;
  wire w7636;
  wire w7637;
  wire w7638;
  wire w7639;
  wire w7640;
  wire w7641;
  wire w7642;
  wire w7643;
  wire w7644;
  wire w7645;
  wire w7646;
  wire w7647;
  wire w7648;
  wire w7649;
  wire w7650;
  wire w7651;
  wire w7652;
  wire w7653;
  wire w7654;
  wire w7655;
  wire w7656;
  wire w7657;
  wire w7658;
  wire w7659;
  wire w7660;
  wire w7661;
  wire w7663;
  wire w7664;
  wire w7665;
  wire w7666;
  wire w7667;
  wire w7668;
  wire w7669;
  wire w7670;
  wire w7671;
  wire w7672;
  wire w7673;
  wire w7674;
  wire w7675;
  wire w7676;
  wire w7677;
  wire w7678;
  wire w7679;
  wire w7680;
  wire w7681;
  wire w7682;
  wire w7683;
  wire w7684;
  wire w7685;
  wire w7686;
  wire w7687;
  wire w7688;
  wire w7689;
  wire w7690;
  wire w7691;
  wire w7692;
  wire w7693;
  wire w7694;
  wire w7695;
  wire w7696;
  wire w7697;
  wire w7698;
  wire w7699;
  wire w7700;
  wire w7701;
  wire w7702;
  wire w7703;
  wire w7704;
  wire w7705;
  wire w7706;
  wire w7707;
  wire w7708;
  wire w7709;
  wire w7710;
  wire w7711;
  wire w7712;
  wire w7713;
  wire w7714;
  wire w7715;
  wire w7716;
  wire w7717;
  wire w7718;
  wire w7719;
  wire w7720;
  wire w7721;
  wire w7722;
  wire w7723;
  wire w7724;
  wire w7725;
  wire w7726;
  wire w7727;
  wire w7728;
  wire w7729;
  wire w7730;
  wire w7731;
  wire w7732;
  wire w7733;
  wire w7734;
  wire w7735;
  wire w7736;
  wire w7737;
  wire w7738;
  wire w7739;
  wire w7740;
  wire w7741;
  wire w7742;
  wire w7743;
  wire w7744;
  wire w7745;
  wire w7746;
  wire w7747;
  wire w7748;
  wire w7749;
  wire w7750;
  wire w7751;
  wire w7752;
  wire w7753;
  wire w7754;
  wire w7755;
  wire w7756;
  wire w7757;
  wire w7758;
  wire w7759;
  wire w7760;
  wire w7761;
  wire w7763;
  wire w7764;
  wire w7765;
  wire w7766;
  wire w7767;
  wire w7768;
  wire w7769;
  wire w7770;
  wire w7771;
  wire w7772;
  wire w7773;
  wire w7774;
  wire w7775;
  wire w7776;
  wire w7777;
  wire w7778;
  wire w7779;
  wire w7780;
  wire w7781;
  wire w7782;
  wire w7783;
  wire w7784;
  wire w7785;
  wire w7786;
  wire w7787;
  wire w7788;
  wire w7789;
  wire w7790;
  wire w7791;
  wire w7792;
  wire w7793;
  wire w7794;
  wire w7795;
  wire w7796;
  wire w7797;
  wire w7798;
  wire w7799;
  wire w7800;
  wire w7801;
  wire w7802;
  wire w7803;
  wire w7804;
  wire w7805;
  wire w7806;
  wire w7807;
  wire w7808;
  wire w7809;
  wire w7810;
  wire w7811;
  wire w7812;
  wire w7813;
  wire w7814;
  wire w7815;
  wire w7816;
  wire w7817;
  wire w7818;
  wire w7819;
  wire w7820;
  wire w7821;
  wire w7822;
  wire w7823;
  wire w7824;
  wire w7825;
  wire w7826;
  wire w7827;
  wire w7828;
  wire w7829;
  wire w7830;
  wire w7831;
  wire w7832;
  wire w7833;
  wire w7834;
  wire w7835;
  wire w7836;
  wire w7837;
  wire w7838;
  wire w7839;
  wire w7840;
  wire w7841;
  wire w7842;
  wire w7843;
  wire w7844;
  wire w7845;
  wire w7846;
  wire w7847;
  wire w7848;
  wire w7849;
  wire w7850;
  wire w7851;
  wire w7852;
  wire w7853;
  wire w7854;
  wire w7855;
  wire w7856;
  wire w7857;
  wire w7858;
  wire w7859;
  wire w7860;
  wire w7861;
  wire w7863;
  wire w7864;
  wire w7865;
  wire w7866;
  wire w7867;
  wire w7868;
  wire w7869;
  wire w7870;
  wire w7871;
  wire w7872;
  wire w7873;
  wire w7874;
  wire w7875;
  wire w7876;
  wire w7877;
  wire w7878;
  wire w7879;
  wire w7880;
  wire w7881;
  wire w7882;
  wire w7883;
  wire w7884;
  wire w7885;
  wire w7886;
  wire w7887;
  wire w7888;
  wire w7889;
  wire w7890;
  wire w7891;
  wire w7892;
  wire w7893;
  wire w7894;
  wire w7895;
  wire w7896;
  wire w7897;
  wire w7898;
  wire w7899;
  wire w7900;
  wire w7901;
  wire w7902;
  wire w7903;
  wire w7904;
  wire w7905;
  wire w7906;
  wire w7907;
  wire w7908;
  wire w7909;
  wire w7910;
  wire w7911;
  wire w7912;
  wire w7913;
  wire w7914;
  wire w7915;
  wire w7916;
  wire w7917;
  wire w7918;
  wire w7919;
  wire w7920;
  wire w7921;
  wire w7922;
  wire w7923;
  wire w7924;
  wire w7925;
  wire w7926;
  wire w7927;
  wire w7928;
  wire w7929;
  wire w7930;
  wire w7931;
  wire w7932;
  wire w7933;
  wire w7934;
  wire w7935;
  wire w7936;
  wire w7937;
  wire w7938;
  wire w7939;
  wire w7940;
  wire w7941;
  wire w7942;
  wire w7943;
  wire w7944;
  wire w7945;
  wire w7946;
  wire w7947;
  wire w7948;
  wire w7949;
  wire w7950;
  wire w7951;
  wire w7952;
  wire w7953;
  wire w7954;
  wire w7955;
  wire w7956;
  wire w7957;
  wire w7958;
  wire w7959;
  wire w7960;
  wire w7961;
  wire w7963;
  wire w7964;
  wire w7965;
  wire w7966;
  wire w7967;
  wire w7968;
  wire w7969;
  wire w7970;
  wire w7971;
  wire w7972;
  wire w7973;
  wire w7974;
  wire w7975;
  wire w7976;
  wire w7977;
  wire w7978;
  wire w7979;
  wire w7980;
  wire w7981;
  wire w7982;
  wire w7983;
  wire w7984;
  wire w7985;
  wire w7986;
  wire w7987;
  wire w7988;
  wire w7989;
  wire w7990;
  wire w7991;
  wire w7992;
  wire w7993;
  wire w7994;
  wire w7995;
  wire w7996;
  wire w7997;
  wire w7998;
  wire w7999;
  wire w8000;
  wire w8001;
  wire w8002;
  wire w8003;
  wire w8004;
  wire w8005;
  wire w8006;
  wire w8007;
  wire w8008;
  wire w8009;
  wire w8010;
  wire w8011;
  wire w8012;
  wire w8013;
  wire w8014;
  wire w8015;
  wire w8016;
  wire w8017;
  wire w8018;
  wire w8019;
  wire w8020;
  wire w8021;
  wire w8022;
  wire w8023;
  wire w8024;
  wire w8025;
  wire w8026;
  wire w8027;
  wire w8028;
  wire w8029;
  wire w8030;
  wire w8031;
  wire w8032;
  wire w8033;
  wire w8034;
  wire w8035;
  wire w8036;
  wire w8037;
  wire w8038;
  wire w8039;
  wire w8040;
  wire w8041;
  wire w8042;
  wire w8043;
  wire w8044;
  wire w8045;
  wire w8046;
  wire w8047;
  wire w8048;
  wire w8049;
  wire w8050;
  wire w8051;
  wire w8052;
  wire w8053;
  wire w8054;
  wire w8055;
  wire w8056;
  wire w8057;
  wire w8058;
  wire w8059;
  wire w8060;
  wire w8061;
  wire w8063;
  wire w8064;
  wire w8065;
  wire w8066;
  wire w8067;
  wire w8068;
  wire w8069;
  wire w8070;
  wire w8071;
  wire w8072;
  wire w8073;
  wire w8074;
  wire w8075;
  wire w8076;
  wire w8077;
  wire w8078;
  wire w8079;
  wire w8080;
  wire w8081;
  wire w8082;
  wire w8083;
  wire w8084;
  wire w8085;
  wire w8086;
  wire w8087;
  wire w8088;
  wire w8089;
  wire w8090;
  wire w8091;
  wire w8092;
  wire w8093;
  wire w8094;
  wire w8095;
  wire w8096;
  wire w8097;
  wire w8098;
  wire w8099;
  wire w8100;
  wire w8101;
  wire w8102;
  wire w8103;
  wire w8104;
  wire w8105;
  wire w8106;
  wire w8107;
  wire w8108;
  wire w8109;
  wire w8110;
  wire w8111;
  wire w8112;
  wire w8113;
  wire w8114;
  wire w8115;
  wire w8116;
  wire w8117;
  wire w8118;
  wire w8119;
  wire w8120;
  wire w8121;
  wire w8122;
  wire w8123;
  wire w8124;
  wire w8125;
  wire w8126;
  wire w8127;
  wire w8128;
  wire w8129;
  wire w8130;
  wire w8131;
  wire w8132;
  wire w8133;
  wire w8134;
  wire w8135;
  wire w8136;
  wire w8137;
  wire w8138;
  wire w8139;
  wire w8140;
  wire w8141;
  wire w8142;
  wire w8143;
  wire w8144;
  wire w8145;
  wire w8146;
  wire w8147;
  wire w8148;
  wire w8149;
  wire w8150;
  wire w8151;
  wire w8152;
  wire w8153;
  wire w8154;
  wire w8155;
  wire w8156;
  wire w8157;
  wire w8158;
  wire w8159;
  wire w8160;
  wire w8161;
  wire w8163;
  wire w8164;
  wire w8165;
  wire w8166;
  wire w8167;
  wire w8168;
  wire w8169;
  wire w8170;
  wire w8171;
  wire w8172;
  wire w8173;
  wire w8174;
  wire w8175;
  wire w8176;
  wire w8177;
  wire w8178;
  wire w8179;
  wire w8180;
  wire w8181;
  wire w8182;
  wire w8183;
  wire w8184;
  wire w8185;
  wire w8186;
  wire w8187;
  wire w8188;
  wire w8189;
  wire w8190;
  wire w8191;
  wire w8192;
  wire w8193;
  wire w8194;
  wire w8195;
  wire w8196;
  wire w8197;
  wire w8198;
  wire w8199;
  wire w8200;
  wire w8201;
  wire w8202;
  wire w8203;
  wire w8204;
  wire w8205;
  wire w8206;
  wire w8207;
  wire w8208;
  wire w8209;
  wire w8210;
  wire w8211;
  wire w8212;
  wire w8213;
  wire w8214;
  wire w8215;
  wire w8216;
  wire w8217;
  wire w8218;
  wire w8219;
  wire w8220;
  wire w8221;
  wire w8222;
  wire w8223;
  wire w8224;
  wire w8225;
  wire w8226;
  wire w8227;
  wire w8228;
  wire w8229;
  wire w8230;
  wire w8231;
  wire w8232;
  wire w8233;
  wire w8234;
  wire w8235;
  wire w8236;
  wire w8237;
  wire w8238;
  wire w8239;
  wire w8240;
  wire w8241;
  wire w8242;
  wire w8243;
  wire w8244;
  wire w8245;
  wire w8246;
  wire w8247;
  wire w8248;
  wire w8249;
  wire w8250;
  wire w8251;
  wire w8252;
  wire w8253;
  wire w8254;
  wire w8255;
  wire w8256;
  wire w8257;
  wire w8258;
  wire w8259;
  wire w8260;
  wire w8261;
  wire w8263;
  wire w8264;
  wire w8265;
  wire w8266;
  wire w8267;
  wire w8268;
  wire w8269;
  wire w8270;
  wire w8271;
  wire w8272;
  wire w8273;
  wire w8274;
  wire w8275;
  wire w8276;
  wire w8277;
  wire w8278;
  wire w8279;
  wire w8280;
  wire w8281;
  wire w8282;
  wire w8283;
  wire w8284;
  wire w8285;
  wire w8286;
  wire w8287;
  wire w8288;
  wire w8289;
  wire w8290;
  wire w8291;
  wire w8292;
  wire w8293;
  wire w8294;
  wire w8295;
  wire w8296;
  wire w8297;
  wire w8298;
  wire w8299;
  wire w8300;
  wire w8301;
  wire w8302;
  wire w8303;
  wire w8304;
  wire w8305;
  wire w8306;
  wire w8307;
  wire w8308;
  wire w8309;
  wire w8310;
  wire w8311;
  wire w8312;
  wire w8313;
  wire w8314;
  wire w8315;
  wire w8316;
  wire w8317;
  wire w8318;
  wire w8319;
  wire w8320;
  wire w8321;
  wire w8322;
  wire w8323;
  wire w8324;
  wire w8325;
  wire w8326;
  wire w8327;
  wire w8328;
  wire w8329;
  wire w8330;
  wire w8331;
  wire w8332;
  wire w8333;
  wire w8334;
  wire w8335;
  wire w8336;
  wire w8337;
  wire w8338;
  wire w8339;
  wire w8340;
  wire w8341;
  wire w8342;
  wire w8343;
  wire w8344;
  wire w8345;
  wire w8346;
  wire w8347;
  wire w8348;
  wire w8349;
  wire w8350;
  wire w8351;
  wire w8352;
  wire w8353;
  wire w8354;
  wire w8355;
  wire w8356;
  wire w8357;
  wire w8358;
  wire w8359;
  wire w8360;
  wire w8361;
  wire w8363;
  wire w8364;
  wire w8365;
  wire w8366;
  wire w8367;
  wire w8368;
  wire w8369;
  wire w8370;
  wire w8371;
  wire w8372;
  wire w8373;
  wire w8374;
  wire w8375;
  wire w8376;
  wire w8377;
  wire w8378;
  wire w8379;
  wire w8380;
  wire w8381;
  wire w8382;
  wire w8383;
  wire w8384;
  wire w8385;
  wire w8386;
  wire w8387;
  wire w8388;
  wire w8389;
  wire w8390;
  wire w8391;
  wire w8392;
  wire w8393;
  wire w8394;
  wire w8395;
  wire w8396;
  wire w8397;
  wire w8398;
  wire w8399;
  wire w8400;
  wire w8401;
  wire w8402;
  wire w8403;
  wire w8404;
  wire w8405;
  wire w8406;
  wire w8407;
  wire w8408;
  wire w8409;
  wire w8410;
  wire w8411;
  wire w8412;
  wire w8413;
  wire w8414;
  wire w8415;
  wire w8416;
  wire w8417;
  wire w8418;
  wire w8419;
  wire w8420;
  wire w8421;
  wire w8422;
  wire w8423;
  wire w8424;
  wire w8425;
  wire w8426;
  wire w8427;
  wire w8428;
  wire w8429;
  wire w8430;
  wire w8431;
  wire w8432;
  wire w8433;
  wire w8434;
  wire w8435;
  wire w8436;
  wire w8437;
  wire w8438;
  wire w8439;
  wire w8440;
  wire w8441;
  wire w8442;
  wire w8443;
  wire w8444;
  wire w8445;
  wire w8446;
  wire w8447;
  wire w8448;
  wire w8449;
  wire w8450;
  wire w8451;
  wire w8452;
  wire w8453;
  wire w8454;
  wire w8455;
  wire w8456;
  wire w8457;
  wire w8458;
  wire w8459;
  wire w8460;
  wire w8461;
  wire w8463;
  wire w8464;
  wire w8465;
  wire w8466;
  wire w8467;
  wire w8468;
  wire w8469;
  wire w8470;
  wire w8471;
  wire w8472;
  wire w8473;
  wire w8474;
  wire w8475;
  wire w8476;
  wire w8477;
  wire w8478;
  wire w8479;
  wire w8480;
  wire w8481;
  wire w8482;
  wire w8483;
  wire w8484;
  wire w8485;
  wire w8486;
  wire w8487;
  wire w8488;
  wire w8489;
  wire w8490;
  wire w8491;
  wire w8492;
  wire w8493;
  wire w8494;
  wire w8495;
  wire w8496;
  wire w8497;
  wire w8498;
  wire w8499;
  wire w8500;
  wire w8501;
  wire w8502;
  wire w8503;
  wire w8504;
  wire w8505;
  wire w8506;
  wire w8507;
  wire w8508;
  wire w8509;
  wire w8510;
  wire w8511;
  wire w8512;
  wire w8513;
  wire w8514;
  wire w8515;
  wire w8516;
  wire w8517;
  wire w8518;
  wire w8519;
  wire w8520;
  wire w8521;
  wire w8522;
  wire w8523;
  wire w8524;
  wire w8525;
  wire w8526;
  wire w8527;
  wire w8528;
  wire w8529;
  wire w8530;
  wire w8531;
  wire w8532;
  wire w8533;
  wire w8534;
  wire w8535;
  wire w8536;
  wire w8537;
  wire w8538;
  wire w8539;
  wire w8540;
  wire w8541;
  wire w8542;
  wire w8543;
  wire w8544;
  wire w8545;
  wire w8546;
  wire w8547;
  wire w8548;
  wire w8549;
  wire w8550;
  wire w8551;
  wire w8552;
  wire w8553;
  wire w8554;
  wire w8555;
  wire w8556;
  wire w8557;
  wire w8558;
  wire w8559;
  wire w8560;
  wire w8561;
  wire w8563;
  wire w8564;
  wire w8565;
  wire w8566;
  wire w8567;
  wire w8568;
  wire w8569;
  wire w8570;
  wire w8571;
  wire w8572;
  wire w8573;
  wire w8574;
  wire w8575;
  wire w8576;
  wire w8577;
  wire w8578;
  wire w8579;
  wire w8580;
  wire w8581;
  wire w8582;
  wire w8583;
  wire w8584;
  wire w8585;
  wire w8586;
  wire w8587;
  wire w8588;
  wire w8589;
  wire w8590;
  wire w8591;
  wire w8592;
  wire w8593;
  wire w8594;
  wire w8595;
  wire w8596;
  wire w8597;
  wire w8598;
  wire w8599;
  wire w8600;
  wire w8601;
  wire w8602;
  wire w8603;
  wire w8604;
  wire w8605;
  wire w8606;
  wire w8607;
  wire w8608;
  wire w8609;
  wire w8610;
  wire w8611;
  wire w8612;
  wire w8613;
  wire w8614;
  wire w8615;
  wire w8616;
  wire w8617;
  wire w8618;
  wire w8619;
  wire w8620;
  wire w8621;
  wire w8622;
  wire w8623;
  wire w8624;
  wire w8625;
  wire w8626;
  wire w8627;
  wire w8628;
  wire w8629;
  wire w8630;
  wire w8631;
  wire w8632;
  wire w8633;
  wire w8634;
  wire w8635;
  wire w8636;
  wire w8637;
  wire w8638;
  wire w8639;
  wire w8640;
  wire w8641;
  wire w8642;
  wire w8643;
  wire w8644;
  wire w8645;
  wire w8646;
  wire w8647;
  wire w8648;
  wire w8649;
  wire w8650;
  wire w8651;
  wire w8652;
  wire w8653;
  wire w8654;
  wire w8655;
  wire w8656;
  wire w8657;
  wire w8658;
  wire w8659;
  wire w8660;
  wire w8661;
  wire w8663;
  wire w8664;
  wire w8665;
  wire w8666;
  wire w8667;
  wire w8668;
  wire w8669;
  wire w8670;
  wire w8671;
  wire w8672;
  wire w8673;
  wire w8674;
  wire w8675;
  wire w8676;
  wire w8677;
  wire w8678;
  wire w8679;
  wire w8680;
  wire w8681;
  wire w8682;
  wire w8683;
  wire w8684;
  wire w8685;
  wire w8686;
  wire w8687;
  wire w8688;
  wire w8689;
  wire w8690;
  wire w8691;
  wire w8692;
  wire w8693;
  wire w8694;
  wire w8695;
  wire w8696;
  wire w8697;
  wire w8698;
  wire w8699;
  wire w8700;
  wire w8701;
  wire w8702;
  wire w8703;
  wire w8704;
  wire w8705;
  wire w8706;
  wire w8707;
  wire w8708;
  wire w8709;
  wire w8710;
  wire w8711;
  wire w8712;
  wire w8713;
  wire w8714;
  wire w8715;
  wire w8716;
  wire w8717;
  wire w8718;
  wire w8719;
  wire w8720;
  wire w8721;
  wire w8722;
  wire w8723;
  wire w8724;
  wire w8725;
  wire w8726;
  wire w8727;
  wire w8728;
  wire w8729;
  wire w8730;
  wire w8731;
  wire w8732;
  wire w8733;
  wire w8734;
  wire w8735;
  wire w8736;
  wire w8737;
  wire w8738;
  wire w8739;
  wire w8740;
  wire w8741;
  wire w8742;
  wire w8743;
  wire w8744;
  wire w8745;
  wire w8746;
  wire w8747;
  wire w8748;
  wire w8749;
  wire w8750;
  wire w8751;
  wire w8752;
  wire w8753;
  wire w8754;
  wire w8755;
  wire w8756;
  wire w8757;
  wire w8758;
  wire w8759;
  wire w8760;
  wire w8761;
  wire w8763;
  wire w8764;
  wire w8765;
  wire w8766;
  wire w8767;
  wire w8768;
  wire w8769;
  wire w8770;
  wire w8771;
  wire w8772;
  wire w8773;
  wire w8774;
  wire w8775;
  wire w8776;
  wire w8777;
  wire w8778;
  wire w8779;
  wire w8780;
  wire w8781;
  wire w8782;
  wire w8783;
  wire w8784;
  wire w8785;
  wire w8786;
  wire w8787;
  wire w8788;
  wire w8789;
  wire w8790;
  wire w8791;
  wire w8792;
  wire w8793;
  wire w8794;
  wire w8795;
  wire w8796;
  wire w8797;
  wire w8798;
  wire w8799;
  wire w8800;
  wire w8801;
  wire w8802;
  wire w8803;
  wire w8804;
  wire w8805;
  wire w8806;
  wire w8807;
  wire w8808;
  wire w8809;
  wire w8810;
  wire w8811;
  wire w8812;
  wire w8813;
  wire w8814;
  wire w8815;
  wire w8816;
  wire w8817;
  wire w8818;
  wire w8819;
  wire w8820;
  wire w8821;
  wire w8822;
  wire w8823;
  wire w8824;
  wire w8825;
  wire w8826;
  wire w8827;
  wire w8828;
  wire w8829;
  wire w8830;
  wire w8831;
  wire w8832;
  wire w8833;
  wire w8834;
  wire w8835;
  wire w8836;
  wire w8837;
  wire w8838;
  wire w8839;
  wire w8840;
  wire w8841;
  wire w8842;
  wire w8843;
  wire w8844;
  wire w8845;
  wire w8846;
  wire w8847;
  wire w8848;
  wire w8849;
  wire w8850;
  wire w8851;
  wire w8852;
  wire w8853;
  wire w8854;
  wire w8855;
  wire w8856;
  wire w8857;
  wire w8858;
  wire w8859;
  wire w8860;
  wire w8861;
  wire w8863;
  wire w8864;
  wire w8865;
  wire w8866;
  wire w8867;
  wire w8868;
  wire w8869;
  wire w8870;
  wire w8871;
  wire w8872;
  wire w8873;
  wire w8874;
  wire w8875;
  wire w8876;
  wire w8877;
  wire w8878;
  wire w8879;
  wire w8880;
  wire w8881;
  wire w8882;
  wire w8883;
  wire w8884;
  wire w8885;
  wire w8886;
  wire w8887;
  wire w8888;
  wire w8889;
  wire w8890;
  wire w8891;
  wire w8892;
  wire w8893;
  wire w8894;
  wire w8895;
  wire w8896;
  wire w8897;
  wire w8898;
  wire w8899;
  wire w8900;
  wire w8901;
  wire w8902;
  wire w8903;
  wire w8904;
  wire w8905;
  wire w8906;
  wire w8907;
  wire w8908;
  wire w8909;
  wire w8910;
  wire w8911;
  wire w8912;
  wire w8913;
  wire w8914;
  wire w8915;
  wire w8916;
  wire w8917;
  wire w8918;
  wire w8919;
  wire w8920;
  wire w8921;
  wire w8922;
  wire w8923;
  wire w8924;
  wire w8925;
  wire w8926;
  wire w8927;
  wire w8928;
  wire w8929;
  wire w8930;
  wire w8931;
  wire w8932;
  wire w8933;
  wire w8934;
  wire w8935;
  wire w8936;
  wire w8937;
  wire w8938;
  wire w8939;
  wire w8940;
  wire w8941;
  wire w8942;
  wire w8943;
  wire w8944;
  wire w8945;
  wire w8946;
  wire w8947;
  wire w8948;
  wire w8949;
  wire w8950;
  wire w8951;
  wire w8952;
  wire w8953;
  wire w8954;
  wire w8955;
  wire w8956;
  wire w8957;
  wire w8958;
  wire w8959;
  wire w8960;
  wire w8961;
  wire w8963;
  wire w8964;
  wire w8965;
  wire w8966;
  wire w8967;
  wire w8968;
  wire w8969;
  wire w8970;
  wire w8971;
  wire w8972;
  wire w8973;
  wire w8974;
  wire w8975;
  wire w8976;
  wire w8977;
  wire w8978;
  wire w8979;
  wire w8980;
  wire w8981;
  wire w8982;
  wire w8983;
  wire w8984;
  wire w8985;
  wire w8986;
  wire w8987;
  wire w8988;
  wire w8989;
  wire w8990;
  wire w8991;
  wire w8992;
  wire w8993;
  wire w8994;
  wire w8995;
  wire w8996;
  wire w8997;
  wire w8998;
  wire w8999;
  wire w9000;
  wire w9001;
  wire w9002;
  wire w9003;
  wire w9004;
  wire w9005;
  wire w9006;
  wire w9007;
  wire w9008;
  wire w9009;
  wire w9010;
  wire w9011;
  wire w9012;
  wire w9013;
  wire w9014;
  wire w9015;
  wire w9016;
  wire w9017;
  wire w9018;
  wire w9019;
  wire w9020;
  wire w9021;
  wire w9022;
  wire w9023;
  wire w9024;
  wire w9025;
  wire w9026;
  wire w9027;
  wire w9028;
  wire w9029;
  wire w9030;
  wire w9031;
  wire w9032;
  wire w9033;
  wire w9034;
  wire w9035;
  wire w9036;
  wire w9037;
  wire w9038;
  wire w9039;
  wire w9040;
  wire w9041;
  wire w9042;
  wire w9043;
  wire w9044;
  wire w9045;
  wire w9046;
  wire w9047;
  wire w9048;
  wire w9049;
  wire w9050;
  wire w9051;
  wire w9052;
  wire w9053;
  wire w9054;
  wire w9055;
  wire w9056;
  wire w9057;
  wire w9058;
  wire w9059;
  wire w9060;
  wire w9061;
  wire w9063;
  wire w9064;
  wire w9065;
  wire w9066;
  wire w9067;
  wire w9068;
  wire w9069;
  wire w9070;
  wire w9071;
  wire w9072;
  wire w9073;
  wire w9074;
  wire w9075;
  wire w9076;
  wire w9077;
  wire w9078;
  wire w9079;
  wire w9080;
  wire w9081;
  wire w9082;
  wire w9083;
  wire w9084;
  wire w9085;
  wire w9086;
  wire w9087;
  wire w9088;
  wire w9089;
  wire w9090;
  wire w9091;
  wire w9092;
  wire w9093;
  wire w9094;
  wire w9095;
  wire w9096;
  wire w9097;
  wire w9098;
  wire w9099;
  wire w9100;
  wire w9101;
  wire w9102;
  wire w9103;
  wire w9104;
  wire w9105;
  wire w9106;
  wire w9107;
  wire w9108;
  wire w9109;
  wire w9110;
  wire w9111;
  wire w9112;
  wire w9113;
  wire w9114;
  wire w9115;
  wire w9116;
  wire w9117;
  wire w9118;
  wire w9119;
  wire w9120;
  wire w9121;
  wire w9122;
  wire w9123;
  wire w9124;
  wire w9125;
  wire w9126;
  wire w9127;
  wire w9128;
  wire w9129;
  wire w9130;
  wire w9131;
  wire w9132;
  wire w9133;
  wire w9134;
  wire w9135;
  wire w9136;
  wire w9137;
  wire w9138;
  wire w9139;
  wire w9140;
  wire w9141;
  wire w9142;
  wire w9143;
  wire w9144;
  wire w9145;
  wire w9146;
  wire w9147;
  wire w9148;
  wire w9149;
  wire w9150;
  wire w9151;
  wire w9152;
  wire w9153;
  wire w9154;
  wire w9155;
  wire w9156;
  wire w9157;
  wire w9158;
  wire w9159;
  wire w9160;
  wire w9161;
  wire w9163;
  wire w9165;
  wire w9167;
  wire w9169;
  wire w9171;
  wire w9173;
  wire w9175;
  wire w9177;
  wire w9179;
  wire w9181;
  wire w9183;
  wire w9185;
  wire w9187;
  wire w9189;
  wire w9191;
  wire w9193;
  wire w9195;
  wire w9197;
  wire w9199;
  wire w9201;
  wire w9203;
  wire w9205;
  wire w9207;
  wire w9209;
  wire w9211;
  wire w9213;
  wire w9215;
  wire w9217;
  wire w9219;
  wire w9221;
  wire w9223;
  wire w9225;
  wire w9227;
  wire w9229;
  wire w9231;
  wire w9233;
  wire w9235;
  wire w9237;
  wire w9239;
  wire w9241;
  wire w9243;
  wire w9245;
  wire w9247;
  wire w9249;
  wire w9251;
  wire w9253;
  wire w9255;
  wire w9257;
  wire w9259;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w3163);
  FullAdder U1 (w3163, IN2[0], IN2[1], w3164, w3165);
  FullAdder U2 (w3165, IN3[0], IN3[1], w3166, w3167);
  FullAdder U3 (w3167, IN4[0], IN4[1], w3168, w3169);
  FullAdder U4 (w3169, IN5[0], IN5[1], w3170, w3171);
  FullAdder U5 (w3171, IN6[0], IN6[1], w3172, w3173);
  FullAdder U6 (w3173, IN7[0], IN7[1], w3174, w3175);
  FullAdder U7 (w3175, IN8[0], IN8[1], w3176, w3177);
  FullAdder U8 (w3177, IN9[0], IN9[1], w3178, w3179);
  FullAdder U9 (w3179, IN10[0], IN10[1], w3180, w3181);
  FullAdder U10 (w3181, IN11[0], IN11[1], w3182, w3183);
  FullAdder U11 (w3183, IN12[0], IN12[1], w3184, w3185);
  FullAdder U12 (w3185, IN13[0], IN13[1], w3186, w3187);
  FullAdder U13 (w3187, IN14[0], IN14[1], w3188, w3189);
  FullAdder U14 (w3189, IN15[0], IN15[1], w3190, w3191);
  FullAdder U15 (w3191, IN16[0], IN16[1], w3192, w3193);
  FullAdder U16 (w3193, IN17[0], IN17[1], w3194, w3195);
  FullAdder U17 (w3195, IN18[0], IN18[1], w3196, w3197);
  FullAdder U18 (w3197, IN19[0], IN19[1], w3198, w3199);
  FullAdder U19 (w3199, IN20[0], IN20[1], w3200, w3201);
  FullAdder U20 (w3201, IN21[0], IN21[1], w3202, w3203);
  FullAdder U21 (w3203, IN22[0], IN22[1], w3204, w3205);
  FullAdder U22 (w3205, IN23[0], IN23[1], w3206, w3207);
  FullAdder U23 (w3207, IN24[0], IN24[1], w3208, w3209);
  FullAdder U24 (w3209, IN25[0], IN25[1], w3210, w3211);
  FullAdder U25 (w3211, IN26[0], IN26[1], w3212, w3213);
  FullAdder U26 (w3213, IN27[0], IN27[1], w3214, w3215);
  FullAdder U27 (w3215, IN28[0], IN28[1], w3216, w3217);
  FullAdder U28 (w3217, IN29[0], IN29[1], w3218, w3219);
  FullAdder U29 (w3219, IN30[0], IN30[1], w3220, w3221);
  FullAdder U30 (w3221, IN31[0], IN31[1], w3222, w3223);
  FullAdder U31 (w3223, IN32[0], IN32[1], w3224, w3225);
  FullAdder U32 (w3225, IN33[0], IN33[1], w3226, w3227);
  FullAdder U33 (w3227, IN34[0], IN34[1], w3228, w3229);
  FullAdder U34 (w3229, IN35[0], IN35[1], w3230, w3231);
  FullAdder U35 (w3231, IN36[0], IN36[1], w3232, w3233);
  FullAdder U36 (w3233, IN37[0], IN37[1], w3234, w3235);
  FullAdder U37 (w3235, IN38[0], IN38[1], w3236, w3237);
  FullAdder U38 (w3237, IN39[0], IN39[1], w3238, w3239);
  FullAdder U39 (w3239, IN40[0], IN40[1], w3240, w3241);
  FullAdder U40 (w3241, IN41[0], IN41[1], w3242, w3243);
  FullAdder U41 (w3243, IN42[0], IN42[1], w3244, w3245);
  FullAdder U42 (w3245, IN43[0], IN43[1], w3246, w3247);
  FullAdder U43 (w3247, IN44[0], IN44[1], w3248, w3249);
  FullAdder U44 (w3249, IN45[0], IN45[1], w3250, w3251);
  FullAdder U45 (w3251, IN46[0], IN46[1], w3252, w3253);
  FullAdder U46 (w3253, IN47[0], IN47[1], w3254, w3255);
  FullAdder U47 (w3255, IN48[0], IN48[1], w3256, w3257);
  FullAdder U48 (w3257, IN49[0], IN49[1], w3258, w3259);
  FullAdder U49 (w3259, IN50[0], IN50[1], w3260, w3261);
  HalfAdder U50 (w3164, IN2[2], Out1[2], w3263);
  FullAdder U51 (w3263, w3166, IN3[2], w3264, w3265);
  FullAdder U52 (w3265, w3168, IN4[2], w3266, w3267);
  FullAdder U53 (w3267, w3170, IN5[2], w3268, w3269);
  FullAdder U54 (w3269, w3172, IN6[2], w3270, w3271);
  FullAdder U55 (w3271, w3174, IN7[2], w3272, w3273);
  FullAdder U56 (w3273, w3176, IN8[2], w3274, w3275);
  FullAdder U57 (w3275, w3178, IN9[2], w3276, w3277);
  FullAdder U58 (w3277, w3180, IN10[2], w3278, w3279);
  FullAdder U59 (w3279, w3182, IN11[2], w3280, w3281);
  FullAdder U60 (w3281, w3184, IN12[2], w3282, w3283);
  FullAdder U61 (w3283, w3186, IN13[2], w3284, w3285);
  FullAdder U62 (w3285, w3188, IN14[2], w3286, w3287);
  FullAdder U63 (w3287, w3190, IN15[2], w3288, w3289);
  FullAdder U64 (w3289, w3192, IN16[2], w3290, w3291);
  FullAdder U65 (w3291, w3194, IN17[2], w3292, w3293);
  FullAdder U66 (w3293, w3196, IN18[2], w3294, w3295);
  FullAdder U67 (w3295, w3198, IN19[2], w3296, w3297);
  FullAdder U68 (w3297, w3200, IN20[2], w3298, w3299);
  FullAdder U69 (w3299, w3202, IN21[2], w3300, w3301);
  FullAdder U70 (w3301, w3204, IN22[2], w3302, w3303);
  FullAdder U71 (w3303, w3206, IN23[2], w3304, w3305);
  FullAdder U72 (w3305, w3208, IN24[2], w3306, w3307);
  FullAdder U73 (w3307, w3210, IN25[2], w3308, w3309);
  FullAdder U74 (w3309, w3212, IN26[2], w3310, w3311);
  FullAdder U75 (w3311, w3214, IN27[2], w3312, w3313);
  FullAdder U76 (w3313, w3216, IN28[2], w3314, w3315);
  FullAdder U77 (w3315, w3218, IN29[2], w3316, w3317);
  FullAdder U78 (w3317, w3220, IN30[2], w3318, w3319);
  FullAdder U79 (w3319, w3222, IN31[2], w3320, w3321);
  FullAdder U80 (w3321, w3224, IN32[2], w3322, w3323);
  FullAdder U81 (w3323, w3226, IN33[2], w3324, w3325);
  FullAdder U82 (w3325, w3228, IN34[2], w3326, w3327);
  FullAdder U83 (w3327, w3230, IN35[2], w3328, w3329);
  FullAdder U84 (w3329, w3232, IN36[2], w3330, w3331);
  FullAdder U85 (w3331, w3234, IN37[2], w3332, w3333);
  FullAdder U86 (w3333, w3236, IN38[2], w3334, w3335);
  FullAdder U87 (w3335, w3238, IN39[2], w3336, w3337);
  FullAdder U88 (w3337, w3240, IN40[2], w3338, w3339);
  FullAdder U89 (w3339, w3242, IN41[2], w3340, w3341);
  FullAdder U90 (w3341, w3244, IN42[2], w3342, w3343);
  FullAdder U91 (w3343, w3246, IN43[2], w3344, w3345);
  FullAdder U92 (w3345, w3248, IN44[2], w3346, w3347);
  FullAdder U93 (w3347, w3250, IN45[2], w3348, w3349);
  FullAdder U94 (w3349, w3252, IN46[2], w3350, w3351);
  FullAdder U95 (w3351, w3254, IN47[2], w3352, w3353);
  FullAdder U96 (w3353, w3256, IN48[2], w3354, w3355);
  FullAdder U97 (w3355, w3258, IN49[2], w3356, w3357);
  FullAdder U98 (w3357, w3260, IN50[2], w3358, w3359);
  FullAdder U99 (w3359, w3261, IN51[0], w3360, w3361);
  HalfAdder U100 (w3264, IN3[3], Out1[3], w3363);
  FullAdder U101 (w3363, w3266, IN4[3], w3364, w3365);
  FullAdder U102 (w3365, w3268, IN5[3], w3366, w3367);
  FullAdder U103 (w3367, w3270, IN6[3], w3368, w3369);
  FullAdder U104 (w3369, w3272, IN7[3], w3370, w3371);
  FullAdder U105 (w3371, w3274, IN8[3], w3372, w3373);
  FullAdder U106 (w3373, w3276, IN9[3], w3374, w3375);
  FullAdder U107 (w3375, w3278, IN10[3], w3376, w3377);
  FullAdder U108 (w3377, w3280, IN11[3], w3378, w3379);
  FullAdder U109 (w3379, w3282, IN12[3], w3380, w3381);
  FullAdder U110 (w3381, w3284, IN13[3], w3382, w3383);
  FullAdder U111 (w3383, w3286, IN14[3], w3384, w3385);
  FullAdder U112 (w3385, w3288, IN15[3], w3386, w3387);
  FullAdder U113 (w3387, w3290, IN16[3], w3388, w3389);
  FullAdder U114 (w3389, w3292, IN17[3], w3390, w3391);
  FullAdder U115 (w3391, w3294, IN18[3], w3392, w3393);
  FullAdder U116 (w3393, w3296, IN19[3], w3394, w3395);
  FullAdder U117 (w3395, w3298, IN20[3], w3396, w3397);
  FullAdder U118 (w3397, w3300, IN21[3], w3398, w3399);
  FullAdder U119 (w3399, w3302, IN22[3], w3400, w3401);
  FullAdder U120 (w3401, w3304, IN23[3], w3402, w3403);
  FullAdder U121 (w3403, w3306, IN24[3], w3404, w3405);
  FullAdder U122 (w3405, w3308, IN25[3], w3406, w3407);
  FullAdder U123 (w3407, w3310, IN26[3], w3408, w3409);
  FullAdder U124 (w3409, w3312, IN27[3], w3410, w3411);
  FullAdder U125 (w3411, w3314, IN28[3], w3412, w3413);
  FullAdder U126 (w3413, w3316, IN29[3], w3414, w3415);
  FullAdder U127 (w3415, w3318, IN30[3], w3416, w3417);
  FullAdder U128 (w3417, w3320, IN31[3], w3418, w3419);
  FullAdder U129 (w3419, w3322, IN32[3], w3420, w3421);
  FullAdder U130 (w3421, w3324, IN33[3], w3422, w3423);
  FullAdder U131 (w3423, w3326, IN34[3], w3424, w3425);
  FullAdder U132 (w3425, w3328, IN35[3], w3426, w3427);
  FullAdder U133 (w3427, w3330, IN36[3], w3428, w3429);
  FullAdder U134 (w3429, w3332, IN37[3], w3430, w3431);
  FullAdder U135 (w3431, w3334, IN38[3], w3432, w3433);
  FullAdder U136 (w3433, w3336, IN39[3], w3434, w3435);
  FullAdder U137 (w3435, w3338, IN40[3], w3436, w3437);
  FullAdder U138 (w3437, w3340, IN41[3], w3438, w3439);
  FullAdder U139 (w3439, w3342, IN42[3], w3440, w3441);
  FullAdder U140 (w3441, w3344, IN43[3], w3442, w3443);
  FullAdder U141 (w3443, w3346, IN44[3], w3444, w3445);
  FullAdder U142 (w3445, w3348, IN45[3], w3446, w3447);
  FullAdder U143 (w3447, w3350, IN46[3], w3448, w3449);
  FullAdder U144 (w3449, w3352, IN47[3], w3450, w3451);
  FullAdder U145 (w3451, w3354, IN48[3], w3452, w3453);
  FullAdder U146 (w3453, w3356, IN49[3], w3454, w3455);
  FullAdder U147 (w3455, w3358, IN50[3], w3456, w3457);
  FullAdder U148 (w3457, w3360, IN51[1], w3458, w3459);
  FullAdder U149 (w3459, w3361, IN52[0], w3460, w3461);
  HalfAdder U150 (w3364, IN4[4], Out1[4], w3463);
  FullAdder U151 (w3463, w3366, IN5[4], w3464, w3465);
  FullAdder U152 (w3465, w3368, IN6[4], w3466, w3467);
  FullAdder U153 (w3467, w3370, IN7[4], w3468, w3469);
  FullAdder U154 (w3469, w3372, IN8[4], w3470, w3471);
  FullAdder U155 (w3471, w3374, IN9[4], w3472, w3473);
  FullAdder U156 (w3473, w3376, IN10[4], w3474, w3475);
  FullAdder U157 (w3475, w3378, IN11[4], w3476, w3477);
  FullAdder U158 (w3477, w3380, IN12[4], w3478, w3479);
  FullAdder U159 (w3479, w3382, IN13[4], w3480, w3481);
  FullAdder U160 (w3481, w3384, IN14[4], w3482, w3483);
  FullAdder U161 (w3483, w3386, IN15[4], w3484, w3485);
  FullAdder U162 (w3485, w3388, IN16[4], w3486, w3487);
  FullAdder U163 (w3487, w3390, IN17[4], w3488, w3489);
  FullAdder U164 (w3489, w3392, IN18[4], w3490, w3491);
  FullAdder U165 (w3491, w3394, IN19[4], w3492, w3493);
  FullAdder U166 (w3493, w3396, IN20[4], w3494, w3495);
  FullAdder U167 (w3495, w3398, IN21[4], w3496, w3497);
  FullAdder U168 (w3497, w3400, IN22[4], w3498, w3499);
  FullAdder U169 (w3499, w3402, IN23[4], w3500, w3501);
  FullAdder U170 (w3501, w3404, IN24[4], w3502, w3503);
  FullAdder U171 (w3503, w3406, IN25[4], w3504, w3505);
  FullAdder U172 (w3505, w3408, IN26[4], w3506, w3507);
  FullAdder U173 (w3507, w3410, IN27[4], w3508, w3509);
  FullAdder U174 (w3509, w3412, IN28[4], w3510, w3511);
  FullAdder U175 (w3511, w3414, IN29[4], w3512, w3513);
  FullAdder U176 (w3513, w3416, IN30[4], w3514, w3515);
  FullAdder U177 (w3515, w3418, IN31[4], w3516, w3517);
  FullAdder U178 (w3517, w3420, IN32[4], w3518, w3519);
  FullAdder U179 (w3519, w3422, IN33[4], w3520, w3521);
  FullAdder U180 (w3521, w3424, IN34[4], w3522, w3523);
  FullAdder U181 (w3523, w3426, IN35[4], w3524, w3525);
  FullAdder U182 (w3525, w3428, IN36[4], w3526, w3527);
  FullAdder U183 (w3527, w3430, IN37[4], w3528, w3529);
  FullAdder U184 (w3529, w3432, IN38[4], w3530, w3531);
  FullAdder U185 (w3531, w3434, IN39[4], w3532, w3533);
  FullAdder U186 (w3533, w3436, IN40[4], w3534, w3535);
  FullAdder U187 (w3535, w3438, IN41[4], w3536, w3537);
  FullAdder U188 (w3537, w3440, IN42[4], w3538, w3539);
  FullAdder U189 (w3539, w3442, IN43[4], w3540, w3541);
  FullAdder U190 (w3541, w3444, IN44[4], w3542, w3543);
  FullAdder U191 (w3543, w3446, IN45[4], w3544, w3545);
  FullAdder U192 (w3545, w3448, IN46[4], w3546, w3547);
  FullAdder U193 (w3547, w3450, IN47[4], w3548, w3549);
  FullAdder U194 (w3549, w3452, IN48[4], w3550, w3551);
  FullAdder U195 (w3551, w3454, IN49[4], w3552, w3553);
  FullAdder U196 (w3553, w3456, IN50[4], w3554, w3555);
  FullAdder U197 (w3555, w3458, IN51[2], w3556, w3557);
  FullAdder U198 (w3557, w3460, IN52[1], w3558, w3559);
  FullAdder U199 (w3559, w3461, IN53[0], w3560, w3561);
  HalfAdder U200 (w3464, IN5[5], Out1[5], w3563);
  FullAdder U201 (w3563, w3466, IN6[5], w3564, w3565);
  FullAdder U202 (w3565, w3468, IN7[5], w3566, w3567);
  FullAdder U203 (w3567, w3470, IN8[5], w3568, w3569);
  FullAdder U204 (w3569, w3472, IN9[5], w3570, w3571);
  FullAdder U205 (w3571, w3474, IN10[5], w3572, w3573);
  FullAdder U206 (w3573, w3476, IN11[5], w3574, w3575);
  FullAdder U207 (w3575, w3478, IN12[5], w3576, w3577);
  FullAdder U208 (w3577, w3480, IN13[5], w3578, w3579);
  FullAdder U209 (w3579, w3482, IN14[5], w3580, w3581);
  FullAdder U210 (w3581, w3484, IN15[5], w3582, w3583);
  FullAdder U211 (w3583, w3486, IN16[5], w3584, w3585);
  FullAdder U212 (w3585, w3488, IN17[5], w3586, w3587);
  FullAdder U213 (w3587, w3490, IN18[5], w3588, w3589);
  FullAdder U214 (w3589, w3492, IN19[5], w3590, w3591);
  FullAdder U215 (w3591, w3494, IN20[5], w3592, w3593);
  FullAdder U216 (w3593, w3496, IN21[5], w3594, w3595);
  FullAdder U217 (w3595, w3498, IN22[5], w3596, w3597);
  FullAdder U218 (w3597, w3500, IN23[5], w3598, w3599);
  FullAdder U219 (w3599, w3502, IN24[5], w3600, w3601);
  FullAdder U220 (w3601, w3504, IN25[5], w3602, w3603);
  FullAdder U221 (w3603, w3506, IN26[5], w3604, w3605);
  FullAdder U222 (w3605, w3508, IN27[5], w3606, w3607);
  FullAdder U223 (w3607, w3510, IN28[5], w3608, w3609);
  FullAdder U224 (w3609, w3512, IN29[5], w3610, w3611);
  FullAdder U225 (w3611, w3514, IN30[5], w3612, w3613);
  FullAdder U226 (w3613, w3516, IN31[5], w3614, w3615);
  FullAdder U227 (w3615, w3518, IN32[5], w3616, w3617);
  FullAdder U228 (w3617, w3520, IN33[5], w3618, w3619);
  FullAdder U229 (w3619, w3522, IN34[5], w3620, w3621);
  FullAdder U230 (w3621, w3524, IN35[5], w3622, w3623);
  FullAdder U231 (w3623, w3526, IN36[5], w3624, w3625);
  FullAdder U232 (w3625, w3528, IN37[5], w3626, w3627);
  FullAdder U233 (w3627, w3530, IN38[5], w3628, w3629);
  FullAdder U234 (w3629, w3532, IN39[5], w3630, w3631);
  FullAdder U235 (w3631, w3534, IN40[5], w3632, w3633);
  FullAdder U236 (w3633, w3536, IN41[5], w3634, w3635);
  FullAdder U237 (w3635, w3538, IN42[5], w3636, w3637);
  FullAdder U238 (w3637, w3540, IN43[5], w3638, w3639);
  FullAdder U239 (w3639, w3542, IN44[5], w3640, w3641);
  FullAdder U240 (w3641, w3544, IN45[5], w3642, w3643);
  FullAdder U241 (w3643, w3546, IN46[5], w3644, w3645);
  FullAdder U242 (w3645, w3548, IN47[5], w3646, w3647);
  FullAdder U243 (w3647, w3550, IN48[5], w3648, w3649);
  FullAdder U244 (w3649, w3552, IN49[5], w3650, w3651);
  FullAdder U245 (w3651, w3554, IN50[5], w3652, w3653);
  FullAdder U246 (w3653, w3556, IN51[3], w3654, w3655);
  FullAdder U247 (w3655, w3558, IN52[2], w3656, w3657);
  FullAdder U248 (w3657, w3560, IN53[1], w3658, w3659);
  FullAdder U249 (w3659, w3561, IN54[0], w3660, w3661);
  HalfAdder U250 (w3564, IN6[6], Out1[6], w3663);
  FullAdder U251 (w3663, w3566, IN7[6], w3664, w3665);
  FullAdder U252 (w3665, w3568, IN8[6], w3666, w3667);
  FullAdder U253 (w3667, w3570, IN9[6], w3668, w3669);
  FullAdder U254 (w3669, w3572, IN10[6], w3670, w3671);
  FullAdder U255 (w3671, w3574, IN11[6], w3672, w3673);
  FullAdder U256 (w3673, w3576, IN12[6], w3674, w3675);
  FullAdder U257 (w3675, w3578, IN13[6], w3676, w3677);
  FullAdder U258 (w3677, w3580, IN14[6], w3678, w3679);
  FullAdder U259 (w3679, w3582, IN15[6], w3680, w3681);
  FullAdder U260 (w3681, w3584, IN16[6], w3682, w3683);
  FullAdder U261 (w3683, w3586, IN17[6], w3684, w3685);
  FullAdder U262 (w3685, w3588, IN18[6], w3686, w3687);
  FullAdder U263 (w3687, w3590, IN19[6], w3688, w3689);
  FullAdder U264 (w3689, w3592, IN20[6], w3690, w3691);
  FullAdder U265 (w3691, w3594, IN21[6], w3692, w3693);
  FullAdder U266 (w3693, w3596, IN22[6], w3694, w3695);
  FullAdder U267 (w3695, w3598, IN23[6], w3696, w3697);
  FullAdder U268 (w3697, w3600, IN24[6], w3698, w3699);
  FullAdder U269 (w3699, w3602, IN25[6], w3700, w3701);
  FullAdder U270 (w3701, w3604, IN26[6], w3702, w3703);
  FullAdder U271 (w3703, w3606, IN27[6], w3704, w3705);
  FullAdder U272 (w3705, w3608, IN28[6], w3706, w3707);
  FullAdder U273 (w3707, w3610, IN29[6], w3708, w3709);
  FullAdder U274 (w3709, w3612, IN30[6], w3710, w3711);
  FullAdder U275 (w3711, w3614, IN31[6], w3712, w3713);
  FullAdder U276 (w3713, w3616, IN32[6], w3714, w3715);
  FullAdder U277 (w3715, w3618, IN33[6], w3716, w3717);
  FullAdder U278 (w3717, w3620, IN34[6], w3718, w3719);
  FullAdder U279 (w3719, w3622, IN35[6], w3720, w3721);
  FullAdder U280 (w3721, w3624, IN36[6], w3722, w3723);
  FullAdder U281 (w3723, w3626, IN37[6], w3724, w3725);
  FullAdder U282 (w3725, w3628, IN38[6], w3726, w3727);
  FullAdder U283 (w3727, w3630, IN39[6], w3728, w3729);
  FullAdder U284 (w3729, w3632, IN40[6], w3730, w3731);
  FullAdder U285 (w3731, w3634, IN41[6], w3732, w3733);
  FullAdder U286 (w3733, w3636, IN42[6], w3734, w3735);
  FullAdder U287 (w3735, w3638, IN43[6], w3736, w3737);
  FullAdder U288 (w3737, w3640, IN44[6], w3738, w3739);
  FullAdder U289 (w3739, w3642, IN45[6], w3740, w3741);
  FullAdder U290 (w3741, w3644, IN46[6], w3742, w3743);
  FullAdder U291 (w3743, w3646, IN47[6], w3744, w3745);
  FullAdder U292 (w3745, w3648, IN48[6], w3746, w3747);
  FullAdder U293 (w3747, w3650, IN49[6], w3748, w3749);
  FullAdder U294 (w3749, w3652, IN50[6], w3750, w3751);
  FullAdder U295 (w3751, w3654, IN51[4], w3752, w3753);
  FullAdder U296 (w3753, w3656, IN52[3], w3754, w3755);
  FullAdder U297 (w3755, w3658, IN53[2], w3756, w3757);
  FullAdder U298 (w3757, w3660, IN54[1], w3758, w3759);
  FullAdder U299 (w3759, w3661, IN55[0], w3760, w3761);
  HalfAdder U300 (w3664, IN7[7], Out1[7], w3763);
  FullAdder U301 (w3763, w3666, IN8[7], w3764, w3765);
  FullAdder U302 (w3765, w3668, IN9[7], w3766, w3767);
  FullAdder U303 (w3767, w3670, IN10[7], w3768, w3769);
  FullAdder U304 (w3769, w3672, IN11[7], w3770, w3771);
  FullAdder U305 (w3771, w3674, IN12[7], w3772, w3773);
  FullAdder U306 (w3773, w3676, IN13[7], w3774, w3775);
  FullAdder U307 (w3775, w3678, IN14[7], w3776, w3777);
  FullAdder U308 (w3777, w3680, IN15[7], w3778, w3779);
  FullAdder U309 (w3779, w3682, IN16[7], w3780, w3781);
  FullAdder U310 (w3781, w3684, IN17[7], w3782, w3783);
  FullAdder U311 (w3783, w3686, IN18[7], w3784, w3785);
  FullAdder U312 (w3785, w3688, IN19[7], w3786, w3787);
  FullAdder U313 (w3787, w3690, IN20[7], w3788, w3789);
  FullAdder U314 (w3789, w3692, IN21[7], w3790, w3791);
  FullAdder U315 (w3791, w3694, IN22[7], w3792, w3793);
  FullAdder U316 (w3793, w3696, IN23[7], w3794, w3795);
  FullAdder U317 (w3795, w3698, IN24[7], w3796, w3797);
  FullAdder U318 (w3797, w3700, IN25[7], w3798, w3799);
  FullAdder U319 (w3799, w3702, IN26[7], w3800, w3801);
  FullAdder U320 (w3801, w3704, IN27[7], w3802, w3803);
  FullAdder U321 (w3803, w3706, IN28[7], w3804, w3805);
  FullAdder U322 (w3805, w3708, IN29[7], w3806, w3807);
  FullAdder U323 (w3807, w3710, IN30[7], w3808, w3809);
  FullAdder U324 (w3809, w3712, IN31[7], w3810, w3811);
  FullAdder U325 (w3811, w3714, IN32[7], w3812, w3813);
  FullAdder U326 (w3813, w3716, IN33[7], w3814, w3815);
  FullAdder U327 (w3815, w3718, IN34[7], w3816, w3817);
  FullAdder U328 (w3817, w3720, IN35[7], w3818, w3819);
  FullAdder U329 (w3819, w3722, IN36[7], w3820, w3821);
  FullAdder U330 (w3821, w3724, IN37[7], w3822, w3823);
  FullAdder U331 (w3823, w3726, IN38[7], w3824, w3825);
  FullAdder U332 (w3825, w3728, IN39[7], w3826, w3827);
  FullAdder U333 (w3827, w3730, IN40[7], w3828, w3829);
  FullAdder U334 (w3829, w3732, IN41[7], w3830, w3831);
  FullAdder U335 (w3831, w3734, IN42[7], w3832, w3833);
  FullAdder U336 (w3833, w3736, IN43[7], w3834, w3835);
  FullAdder U337 (w3835, w3738, IN44[7], w3836, w3837);
  FullAdder U338 (w3837, w3740, IN45[7], w3838, w3839);
  FullAdder U339 (w3839, w3742, IN46[7], w3840, w3841);
  FullAdder U340 (w3841, w3744, IN47[7], w3842, w3843);
  FullAdder U341 (w3843, w3746, IN48[7], w3844, w3845);
  FullAdder U342 (w3845, w3748, IN49[7], w3846, w3847);
  FullAdder U343 (w3847, w3750, IN50[7], w3848, w3849);
  FullAdder U344 (w3849, w3752, IN51[5], w3850, w3851);
  FullAdder U345 (w3851, w3754, IN52[4], w3852, w3853);
  FullAdder U346 (w3853, w3756, IN53[3], w3854, w3855);
  FullAdder U347 (w3855, w3758, IN54[2], w3856, w3857);
  FullAdder U348 (w3857, w3760, IN55[1], w3858, w3859);
  FullAdder U349 (w3859, w3761, IN56[0], w3860, w3861);
  HalfAdder U350 (w3764, IN8[8], Out1[8], w3863);
  FullAdder U351 (w3863, w3766, IN9[8], w3864, w3865);
  FullAdder U352 (w3865, w3768, IN10[8], w3866, w3867);
  FullAdder U353 (w3867, w3770, IN11[8], w3868, w3869);
  FullAdder U354 (w3869, w3772, IN12[8], w3870, w3871);
  FullAdder U355 (w3871, w3774, IN13[8], w3872, w3873);
  FullAdder U356 (w3873, w3776, IN14[8], w3874, w3875);
  FullAdder U357 (w3875, w3778, IN15[8], w3876, w3877);
  FullAdder U358 (w3877, w3780, IN16[8], w3878, w3879);
  FullAdder U359 (w3879, w3782, IN17[8], w3880, w3881);
  FullAdder U360 (w3881, w3784, IN18[8], w3882, w3883);
  FullAdder U361 (w3883, w3786, IN19[8], w3884, w3885);
  FullAdder U362 (w3885, w3788, IN20[8], w3886, w3887);
  FullAdder U363 (w3887, w3790, IN21[8], w3888, w3889);
  FullAdder U364 (w3889, w3792, IN22[8], w3890, w3891);
  FullAdder U365 (w3891, w3794, IN23[8], w3892, w3893);
  FullAdder U366 (w3893, w3796, IN24[8], w3894, w3895);
  FullAdder U367 (w3895, w3798, IN25[8], w3896, w3897);
  FullAdder U368 (w3897, w3800, IN26[8], w3898, w3899);
  FullAdder U369 (w3899, w3802, IN27[8], w3900, w3901);
  FullAdder U370 (w3901, w3804, IN28[8], w3902, w3903);
  FullAdder U371 (w3903, w3806, IN29[8], w3904, w3905);
  FullAdder U372 (w3905, w3808, IN30[8], w3906, w3907);
  FullAdder U373 (w3907, w3810, IN31[8], w3908, w3909);
  FullAdder U374 (w3909, w3812, IN32[8], w3910, w3911);
  FullAdder U375 (w3911, w3814, IN33[8], w3912, w3913);
  FullAdder U376 (w3913, w3816, IN34[8], w3914, w3915);
  FullAdder U377 (w3915, w3818, IN35[8], w3916, w3917);
  FullAdder U378 (w3917, w3820, IN36[8], w3918, w3919);
  FullAdder U379 (w3919, w3822, IN37[8], w3920, w3921);
  FullAdder U380 (w3921, w3824, IN38[8], w3922, w3923);
  FullAdder U381 (w3923, w3826, IN39[8], w3924, w3925);
  FullAdder U382 (w3925, w3828, IN40[8], w3926, w3927);
  FullAdder U383 (w3927, w3830, IN41[8], w3928, w3929);
  FullAdder U384 (w3929, w3832, IN42[8], w3930, w3931);
  FullAdder U385 (w3931, w3834, IN43[8], w3932, w3933);
  FullAdder U386 (w3933, w3836, IN44[8], w3934, w3935);
  FullAdder U387 (w3935, w3838, IN45[8], w3936, w3937);
  FullAdder U388 (w3937, w3840, IN46[8], w3938, w3939);
  FullAdder U389 (w3939, w3842, IN47[8], w3940, w3941);
  FullAdder U390 (w3941, w3844, IN48[8], w3942, w3943);
  FullAdder U391 (w3943, w3846, IN49[8], w3944, w3945);
  FullAdder U392 (w3945, w3848, IN50[8], w3946, w3947);
  FullAdder U393 (w3947, w3850, IN51[6], w3948, w3949);
  FullAdder U394 (w3949, w3852, IN52[5], w3950, w3951);
  FullAdder U395 (w3951, w3854, IN53[4], w3952, w3953);
  FullAdder U396 (w3953, w3856, IN54[3], w3954, w3955);
  FullAdder U397 (w3955, w3858, IN55[2], w3956, w3957);
  FullAdder U398 (w3957, w3860, IN56[1], w3958, w3959);
  FullAdder U399 (w3959, w3861, IN57[0], w3960, w3961);
  HalfAdder U400 (w3864, IN9[9], Out1[9], w3963);
  FullAdder U401 (w3963, w3866, IN10[9], w3964, w3965);
  FullAdder U402 (w3965, w3868, IN11[9], w3966, w3967);
  FullAdder U403 (w3967, w3870, IN12[9], w3968, w3969);
  FullAdder U404 (w3969, w3872, IN13[9], w3970, w3971);
  FullAdder U405 (w3971, w3874, IN14[9], w3972, w3973);
  FullAdder U406 (w3973, w3876, IN15[9], w3974, w3975);
  FullAdder U407 (w3975, w3878, IN16[9], w3976, w3977);
  FullAdder U408 (w3977, w3880, IN17[9], w3978, w3979);
  FullAdder U409 (w3979, w3882, IN18[9], w3980, w3981);
  FullAdder U410 (w3981, w3884, IN19[9], w3982, w3983);
  FullAdder U411 (w3983, w3886, IN20[9], w3984, w3985);
  FullAdder U412 (w3985, w3888, IN21[9], w3986, w3987);
  FullAdder U413 (w3987, w3890, IN22[9], w3988, w3989);
  FullAdder U414 (w3989, w3892, IN23[9], w3990, w3991);
  FullAdder U415 (w3991, w3894, IN24[9], w3992, w3993);
  FullAdder U416 (w3993, w3896, IN25[9], w3994, w3995);
  FullAdder U417 (w3995, w3898, IN26[9], w3996, w3997);
  FullAdder U418 (w3997, w3900, IN27[9], w3998, w3999);
  FullAdder U419 (w3999, w3902, IN28[9], w4000, w4001);
  FullAdder U420 (w4001, w3904, IN29[9], w4002, w4003);
  FullAdder U421 (w4003, w3906, IN30[9], w4004, w4005);
  FullAdder U422 (w4005, w3908, IN31[9], w4006, w4007);
  FullAdder U423 (w4007, w3910, IN32[9], w4008, w4009);
  FullAdder U424 (w4009, w3912, IN33[9], w4010, w4011);
  FullAdder U425 (w4011, w3914, IN34[9], w4012, w4013);
  FullAdder U426 (w4013, w3916, IN35[9], w4014, w4015);
  FullAdder U427 (w4015, w3918, IN36[9], w4016, w4017);
  FullAdder U428 (w4017, w3920, IN37[9], w4018, w4019);
  FullAdder U429 (w4019, w3922, IN38[9], w4020, w4021);
  FullAdder U430 (w4021, w3924, IN39[9], w4022, w4023);
  FullAdder U431 (w4023, w3926, IN40[9], w4024, w4025);
  FullAdder U432 (w4025, w3928, IN41[9], w4026, w4027);
  FullAdder U433 (w4027, w3930, IN42[9], w4028, w4029);
  FullAdder U434 (w4029, w3932, IN43[9], w4030, w4031);
  FullAdder U435 (w4031, w3934, IN44[9], w4032, w4033);
  FullAdder U436 (w4033, w3936, IN45[9], w4034, w4035);
  FullAdder U437 (w4035, w3938, IN46[9], w4036, w4037);
  FullAdder U438 (w4037, w3940, IN47[9], w4038, w4039);
  FullAdder U439 (w4039, w3942, IN48[9], w4040, w4041);
  FullAdder U440 (w4041, w3944, IN49[9], w4042, w4043);
  FullAdder U441 (w4043, w3946, IN50[9], w4044, w4045);
  FullAdder U442 (w4045, w3948, IN51[7], w4046, w4047);
  FullAdder U443 (w4047, w3950, IN52[6], w4048, w4049);
  FullAdder U444 (w4049, w3952, IN53[5], w4050, w4051);
  FullAdder U445 (w4051, w3954, IN54[4], w4052, w4053);
  FullAdder U446 (w4053, w3956, IN55[3], w4054, w4055);
  FullAdder U447 (w4055, w3958, IN56[2], w4056, w4057);
  FullAdder U448 (w4057, w3960, IN57[1], w4058, w4059);
  FullAdder U449 (w4059, w3961, IN58[0], w4060, w4061);
  HalfAdder U450 (w3964, IN10[10], Out1[10], w4063);
  FullAdder U451 (w4063, w3966, IN11[10], w4064, w4065);
  FullAdder U452 (w4065, w3968, IN12[10], w4066, w4067);
  FullAdder U453 (w4067, w3970, IN13[10], w4068, w4069);
  FullAdder U454 (w4069, w3972, IN14[10], w4070, w4071);
  FullAdder U455 (w4071, w3974, IN15[10], w4072, w4073);
  FullAdder U456 (w4073, w3976, IN16[10], w4074, w4075);
  FullAdder U457 (w4075, w3978, IN17[10], w4076, w4077);
  FullAdder U458 (w4077, w3980, IN18[10], w4078, w4079);
  FullAdder U459 (w4079, w3982, IN19[10], w4080, w4081);
  FullAdder U460 (w4081, w3984, IN20[10], w4082, w4083);
  FullAdder U461 (w4083, w3986, IN21[10], w4084, w4085);
  FullAdder U462 (w4085, w3988, IN22[10], w4086, w4087);
  FullAdder U463 (w4087, w3990, IN23[10], w4088, w4089);
  FullAdder U464 (w4089, w3992, IN24[10], w4090, w4091);
  FullAdder U465 (w4091, w3994, IN25[10], w4092, w4093);
  FullAdder U466 (w4093, w3996, IN26[10], w4094, w4095);
  FullAdder U467 (w4095, w3998, IN27[10], w4096, w4097);
  FullAdder U468 (w4097, w4000, IN28[10], w4098, w4099);
  FullAdder U469 (w4099, w4002, IN29[10], w4100, w4101);
  FullAdder U470 (w4101, w4004, IN30[10], w4102, w4103);
  FullAdder U471 (w4103, w4006, IN31[10], w4104, w4105);
  FullAdder U472 (w4105, w4008, IN32[10], w4106, w4107);
  FullAdder U473 (w4107, w4010, IN33[10], w4108, w4109);
  FullAdder U474 (w4109, w4012, IN34[10], w4110, w4111);
  FullAdder U475 (w4111, w4014, IN35[10], w4112, w4113);
  FullAdder U476 (w4113, w4016, IN36[10], w4114, w4115);
  FullAdder U477 (w4115, w4018, IN37[10], w4116, w4117);
  FullAdder U478 (w4117, w4020, IN38[10], w4118, w4119);
  FullAdder U479 (w4119, w4022, IN39[10], w4120, w4121);
  FullAdder U480 (w4121, w4024, IN40[10], w4122, w4123);
  FullAdder U481 (w4123, w4026, IN41[10], w4124, w4125);
  FullAdder U482 (w4125, w4028, IN42[10], w4126, w4127);
  FullAdder U483 (w4127, w4030, IN43[10], w4128, w4129);
  FullAdder U484 (w4129, w4032, IN44[10], w4130, w4131);
  FullAdder U485 (w4131, w4034, IN45[10], w4132, w4133);
  FullAdder U486 (w4133, w4036, IN46[10], w4134, w4135);
  FullAdder U487 (w4135, w4038, IN47[10], w4136, w4137);
  FullAdder U488 (w4137, w4040, IN48[10], w4138, w4139);
  FullAdder U489 (w4139, w4042, IN49[10], w4140, w4141);
  FullAdder U490 (w4141, w4044, IN50[10], w4142, w4143);
  FullAdder U491 (w4143, w4046, IN51[8], w4144, w4145);
  FullAdder U492 (w4145, w4048, IN52[7], w4146, w4147);
  FullAdder U493 (w4147, w4050, IN53[6], w4148, w4149);
  FullAdder U494 (w4149, w4052, IN54[5], w4150, w4151);
  FullAdder U495 (w4151, w4054, IN55[4], w4152, w4153);
  FullAdder U496 (w4153, w4056, IN56[3], w4154, w4155);
  FullAdder U497 (w4155, w4058, IN57[2], w4156, w4157);
  FullAdder U498 (w4157, w4060, IN58[1], w4158, w4159);
  FullAdder U499 (w4159, w4061, IN59[0], w4160, w4161);
  HalfAdder U500 (w4064, IN11[11], Out1[11], w4163);
  FullAdder U501 (w4163, w4066, IN12[11], w4164, w4165);
  FullAdder U502 (w4165, w4068, IN13[11], w4166, w4167);
  FullAdder U503 (w4167, w4070, IN14[11], w4168, w4169);
  FullAdder U504 (w4169, w4072, IN15[11], w4170, w4171);
  FullAdder U505 (w4171, w4074, IN16[11], w4172, w4173);
  FullAdder U506 (w4173, w4076, IN17[11], w4174, w4175);
  FullAdder U507 (w4175, w4078, IN18[11], w4176, w4177);
  FullAdder U508 (w4177, w4080, IN19[11], w4178, w4179);
  FullAdder U509 (w4179, w4082, IN20[11], w4180, w4181);
  FullAdder U510 (w4181, w4084, IN21[11], w4182, w4183);
  FullAdder U511 (w4183, w4086, IN22[11], w4184, w4185);
  FullAdder U512 (w4185, w4088, IN23[11], w4186, w4187);
  FullAdder U513 (w4187, w4090, IN24[11], w4188, w4189);
  FullAdder U514 (w4189, w4092, IN25[11], w4190, w4191);
  FullAdder U515 (w4191, w4094, IN26[11], w4192, w4193);
  FullAdder U516 (w4193, w4096, IN27[11], w4194, w4195);
  FullAdder U517 (w4195, w4098, IN28[11], w4196, w4197);
  FullAdder U518 (w4197, w4100, IN29[11], w4198, w4199);
  FullAdder U519 (w4199, w4102, IN30[11], w4200, w4201);
  FullAdder U520 (w4201, w4104, IN31[11], w4202, w4203);
  FullAdder U521 (w4203, w4106, IN32[11], w4204, w4205);
  FullAdder U522 (w4205, w4108, IN33[11], w4206, w4207);
  FullAdder U523 (w4207, w4110, IN34[11], w4208, w4209);
  FullAdder U524 (w4209, w4112, IN35[11], w4210, w4211);
  FullAdder U525 (w4211, w4114, IN36[11], w4212, w4213);
  FullAdder U526 (w4213, w4116, IN37[11], w4214, w4215);
  FullAdder U527 (w4215, w4118, IN38[11], w4216, w4217);
  FullAdder U528 (w4217, w4120, IN39[11], w4218, w4219);
  FullAdder U529 (w4219, w4122, IN40[11], w4220, w4221);
  FullAdder U530 (w4221, w4124, IN41[11], w4222, w4223);
  FullAdder U531 (w4223, w4126, IN42[11], w4224, w4225);
  FullAdder U532 (w4225, w4128, IN43[11], w4226, w4227);
  FullAdder U533 (w4227, w4130, IN44[11], w4228, w4229);
  FullAdder U534 (w4229, w4132, IN45[11], w4230, w4231);
  FullAdder U535 (w4231, w4134, IN46[11], w4232, w4233);
  FullAdder U536 (w4233, w4136, IN47[11], w4234, w4235);
  FullAdder U537 (w4235, w4138, IN48[11], w4236, w4237);
  FullAdder U538 (w4237, w4140, IN49[11], w4238, w4239);
  FullAdder U539 (w4239, w4142, IN50[11], w4240, w4241);
  FullAdder U540 (w4241, w4144, IN51[9], w4242, w4243);
  FullAdder U541 (w4243, w4146, IN52[8], w4244, w4245);
  FullAdder U542 (w4245, w4148, IN53[7], w4246, w4247);
  FullAdder U543 (w4247, w4150, IN54[6], w4248, w4249);
  FullAdder U544 (w4249, w4152, IN55[5], w4250, w4251);
  FullAdder U545 (w4251, w4154, IN56[4], w4252, w4253);
  FullAdder U546 (w4253, w4156, IN57[3], w4254, w4255);
  FullAdder U547 (w4255, w4158, IN58[2], w4256, w4257);
  FullAdder U548 (w4257, w4160, IN59[1], w4258, w4259);
  FullAdder U549 (w4259, w4161, IN60[0], w4260, w4261);
  HalfAdder U550 (w4164, IN12[12], Out1[12], w4263);
  FullAdder U551 (w4263, w4166, IN13[12], w4264, w4265);
  FullAdder U552 (w4265, w4168, IN14[12], w4266, w4267);
  FullAdder U553 (w4267, w4170, IN15[12], w4268, w4269);
  FullAdder U554 (w4269, w4172, IN16[12], w4270, w4271);
  FullAdder U555 (w4271, w4174, IN17[12], w4272, w4273);
  FullAdder U556 (w4273, w4176, IN18[12], w4274, w4275);
  FullAdder U557 (w4275, w4178, IN19[12], w4276, w4277);
  FullAdder U558 (w4277, w4180, IN20[12], w4278, w4279);
  FullAdder U559 (w4279, w4182, IN21[12], w4280, w4281);
  FullAdder U560 (w4281, w4184, IN22[12], w4282, w4283);
  FullAdder U561 (w4283, w4186, IN23[12], w4284, w4285);
  FullAdder U562 (w4285, w4188, IN24[12], w4286, w4287);
  FullAdder U563 (w4287, w4190, IN25[12], w4288, w4289);
  FullAdder U564 (w4289, w4192, IN26[12], w4290, w4291);
  FullAdder U565 (w4291, w4194, IN27[12], w4292, w4293);
  FullAdder U566 (w4293, w4196, IN28[12], w4294, w4295);
  FullAdder U567 (w4295, w4198, IN29[12], w4296, w4297);
  FullAdder U568 (w4297, w4200, IN30[12], w4298, w4299);
  FullAdder U569 (w4299, w4202, IN31[12], w4300, w4301);
  FullAdder U570 (w4301, w4204, IN32[12], w4302, w4303);
  FullAdder U571 (w4303, w4206, IN33[12], w4304, w4305);
  FullAdder U572 (w4305, w4208, IN34[12], w4306, w4307);
  FullAdder U573 (w4307, w4210, IN35[12], w4308, w4309);
  FullAdder U574 (w4309, w4212, IN36[12], w4310, w4311);
  FullAdder U575 (w4311, w4214, IN37[12], w4312, w4313);
  FullAdder U576 (w4313, w4216, IN38[12], w4314, w4315);
  FullAdder U577 (w4315, w4218, IN39[12], w4316, w4317);
  FullAdder U578 (w4317, w4220, IN40[12], w4318, w4319);
  FullAdder U579 (w4319, w4222, IN41[12], w4320, w4321);
  FullAdder U580 (w4321, w4224, IN42[12], w4322, w4323);
  FullAdder U581 (w4323, w4226, IN43[12], w4324, w4325);
  FullAdder U582 (w4325, w4228, IN44[12], w4326, w4327);
  FullAdder U583 (w4327, w4230, IN45[12], w4328, w4329);
  FullAdder U584 (w4329, w4232, IN46[12], w4330, w4331);
  FullAdder U585 (w4331, w4234, IN47[12], w4332, w4333);
  FullAdder U586 (w4333, w4236, IN48[12], w4334, w4335);
  FullAdder U587 (w4335, w4238, IN49[12], w4336, w4337);
  FullAdder U588 (w4337, w4240, IN50[12], w4338, w4339);
  FullAdder U589 (w4339, w4242, IN51[10], w4340, w4341);
  FullAdder U590 (w4341, w4244, IN52[9], w4342, w4343);
  FullAdder U591 (w4343, w4246, IN53[8], w4344, w4345);
  FullAdder U592 (w4345, w4248, IN54[7], w4346, w4347);
  FullAdder U593 (w4347, w4250, IN55[6], w4348, w4349);
  FullAdder U594 (w4349, w4252, IN56[5], w4350, w4351);
  FullAdder U595 (w4351, w4254, IN57[4], w4352, w4353);
  FullAdder U596 (w4353, w4256, IN58[3], w4354, w4355);
  FullAdder U597 (w4355, w4258, IN59[2], w4356, w4357);
  FullAdder U598 (w4357, w4260, IN60[1], w4358, w4359);
  FullAdder U599 (w4359, w4261, IN61[0], w4360, w4361);
  HalfAdder U600 (w4264, IN13[13], Out1[13], w4363);
  FullAdder U601 (w4363, w4266, IN14[13], w4364, w4365);
  FullAdder U602 (w4365, w4268, IN15[13], w4366, w4367);
  FullAdder U603 (w4367, w4270, IN16[13], w4368, w4369);
  FullAdder U604 (w4369, w4272, IN17[13], w4370, w4371);
  FullAdder U605 (w4371, w4274, IN18[13], w4372, w4373);
  FullAdder U606 (w4373, w4276, IN19[13], w4374, w4375);
  FullAdder U607 (w4375, w4278, IN20[13], w4376, w4377);
  FullAdder U608 (w4377, w4280, IN21[13], w4378, w4379);
  FullAdder U609 (w4379, w4282, IN22[13], w4380, w4381);
  FullAdder U610 (w4381, w4284, IN23[13], w4382, w4383);
  FullAdder U611 (w4383, w4286, IN24[13], w4384, w4385);
  FullAdder U612 (w4385, w4288, IN25[13], w4386, w4387);
  FullAdder U613 (w4387, w4290, IN26[13], w4388, w4389);
  FullAdder U614 (w4389, w4292, IN27[13], w4390, w4391);
  FullAdder U615 (w4391, w4294, IN28[13], w4392, w4393);
  FullAdder U616 (w4393, w4296, IN29[13], w4394, w4395);
  FullAdder U617 (w4395, w4298, IN30[13], w4396, w4397);
  FullAdder U618 (w4397, w4300, IN31[13], w4398, w4399);
  FullAdder U619 (w4399, w4302, IN32[13], w4400, w4401);
  FullAdder U620 (w4401, w4304, IN33[13], w4402, w4403);
  FullAdder U621 (w4403, w4306, IN34[13], w4404, w4405);
  FullAdder U622 (w4405, w4308, IN35[13], w4406, w4407);
  FullAdder U623 (w4407, w4310, IN36[13], w4408, w4409);
  FullAdder U624 (w4409, w4312, IN37[13], w4410, w4411);
  FullAdder U625 (w4411, w4314, IN38[13], w4412, w4413);
  FullAdder U626 (w4413, w4316, IN39[13], w4414, w4415);
  FullAdder U627 (w4415, w4318, IN40[13], w4416, w4417);
  FullAdder U628 (w4417, w4320, IN41[13], w4418, w4419);
  FullAdder U629 (w4419, w4322, IN42[13], w4420, w4421);
  FullAdder U630 (w4421, w4324, IN43[13], w4422, w4423);
  FullAdder U631 (w4423, w4326, IN44[13], w4424, w4425);
  FullAdder U632 (w4425, w4328, IN45[13], w4426, w4427);
  FullAdder U633 (w4427, w4330, IN46[13], w4428, w4429);
  FullAdder U634 (w4429, w4332, IN47[13], w4430, w4431);
  FullAdder U635 (w4431, w4334, IN48[13], w4432, w4433);
  FullAdder U636 (w4433, w4336, IN49[13], w4434, w4435);
  FullAdder U637 (w4435, w4338, IN50[13], w4436, w4437);
  FullAdder U638 (w4437, w4340, IN51[11], w4438, w4439);
  FullAdder U639 (w4439, w4342, IN52[10], w4440, w4441);
  FullAdder U640 (w4441, w4344, IN53[9], w4442, w4443);
  FullAdder U641 (w4443, w4346, IN54[8], w4444, w4445);
  FullAdder U642 (w4445, w4348, IN55[7], w4446, w4447);
  FullAdder U643 (w4447, w4350, IN56[6], w4448, w4449);
  FullAdder U644 (w4449, w4352, IN57[5], w4450, w4451);
  FullAdder U645 (w4451, w4354, IN58[4], w4452, w4453);
  FullAdder U646 (w4453, w4356, IN59[3], w4454, w4455);
  FullAdder U647 (w4455, w4358, IN60[2], w4456, w4457);
  FullAdder U648 (w4457, w4360, IN61[1], w4458, w4459);
  FullAdder U649 (w4459, w4361, IN62[0], w4460, w4461);
  HalfAdder U650 (w4364, IN14[14], Out1[14], w4463);
  FullAdder U651 (w4463, w4366, IN15[14], w4464, w4465);
  FullAdder U652 (w4465, w4368, IN16[14], w4466, w4467);
  FullAdder U653 (w4467, w4370, IN17[14], w4468, w4469);
  FullAdder U654 (w4469, w4372, IN18[14], w4470, w4471);
  FullAdder U655 (w4471, w4374, IN19[14], w4472, w4473);
  FullAdder U656 (w4473, w4376, IN20[14], w4474, w4475);
  FullAdder U657 (w4475, w4378, IN21[14], w4476, w4477);
  FullAdder U658 (w4477, w4380, IN22[14], w4478, w4479);
  FullAdder U659 (w4479, w4382, IN23[14], w4480, w4481);
  FullAdder U660 (w4481, w4384, IN24[14], w4482, w4483);
  FullAdder U661 (w4483, w4386, IN25[14], w4484, w4485);
  FullAdder U662 (w4485, w4388, IN26[14], w4486, w4487);
  FullAdder U663 (w4487, w4390, IN27[14], w4488, w4489);
  FullAdder U664 (w4489, w4392, IN28[14], w4490, w4491);
  FullAdder U665 (w4491, w4394, IN29[14], w4492, w4493);
  FullAdder U666 (w4493, w4396, IN30[14], w4494, w4495);
  FullAdder U667 (w4495, w4398, IN31[14], w4496, w4497);
  FullAdder U668 (w4497, w4400, IN32[14], w4498, w4499);
  FullAdder U669 (w4499, w4402, IN33[14], w4500, w4501);
  FullAdder U670 (w4501, w4404, IN34[14], w4502, w4503);
  FullAdder U671 (w4503, w4406, IN35[14], w4504, w4505);
  FullAdder U672 (w4505, w4408, IN36[14], w4506, w4507);
  FullAdder U673 (w4507, w4410, IN37[14], w4508, w4509);
  FullAdder U674 (w4509, w4412, IN38[14], w4510, w4511);
  FullAdder U675 (w4511, w4414, IN39[14], w4512, w4513);
  FullAdder U676 (w4513, w4416, IN40[14], w4514, w4515);
  FullAdder U677 (w4515, w4418, IN41[14], w4516, w4517);
  FullAdder U678 (w4517, w4420, IN42[14], w4518, w4519);
  FullAdder U679 (w4519, w4422, IN43[14], w4520, w4521);
  FullAdder U680 (w4521, w4424, IN44[14], w4522, w4523);
  FullAdder U681 (w4523, w4426, IN45[14], w4524, w4525);
  FullAdder U682 (w4525, w4428, IN46[14], w4526, w4527);
  FullAdder U683 (w4527, w4430, IN47[14], w4528, w4529);
  FullAdder U684 (w4529, w4432, IN48[14], w4530, w4531);
  FullAdder U685 (w4531, w4434, IN49[14], w4532, w4533);
  FullAdder U686 (w4533, w4436, IN50[14], w4534, w4535);
  FullAdder U687 (w4535, w4438, IN51[12], w4536, w4537);
  FullAdder U688 (w4537, w4440, IN52[11], w4538, w4539);
  FullAdder U689 (w4539, w4442, IN53[10], w4540, w4541);
  FullAdder U690 (w4541, w4444, IN54[9], w4542, w4543);
  FullAdder U691 (w4543, w4446, IN55[8], w4544, w4545);
  FullAdder U692 (w4545, w4448, IN56[7], w4546, w4547);
  FullAdder U693 (w4547, w4450, IN57[6], w4548, w4549);
  FullAdder U694 (w4549, w4452, IN58[5], w4550, w4551);
  FullAdder U695 (w4551, w4454, IN59[4], w4552, w4553);
  FullAdder U696 (w4553, w4456, IN60[3], w4554, w4555);
  FullAdder U697 (w4555, w4458, IN61[2], w4556, w4557);
  FullAdder U698 (w4557, w4460, IN62[1], w4558, w4559);
  FullAdder U699 (w4559, w4461, IN63[0], w4560, w4561);
  HalfAdder U700 (w4464, IN15[15], Out1[15], w4563);
  FullAdder U701 (w4563, w4466, IN16[15], w4564, w4565);
  FullAdder U702 (w4565, w4468, IN17[15], w4566, w4567);
  FullAdder U703 (w4567, w4470, IN18[15], w4568, w4569);
  FullAdder U704 (w4569, w4472, IN19[15], w4570, w4571);
  FullAdder U705 (w4571, w4474, IN20[15], w4572, w4573);
  FullAdder U706 (w4573, w4476, IN21[15], w4574, w4575);
  FullAdder U707 (w4575, w4478, IN22[15], w4576, w4577);
  FullAdder U708 (w4577, w4480, IN23[15], w4578, w4579);
  FullAdder U709 (w4579, w4482, IN24[15], w4580, w4581);
  FullAdder U710 (w4581, w4484, IN25[15], w4582, w4583);
  FullAdder U711 (w4583, w4486, IN26[15], w4584, w4585);
  FullAdder U712 (w4585, w4488, IN27[15], w4586, w4587);
  FullAdder U713 (w4587, w4490, IN28[15], w4588, w4589);
  FullAdder U714 (w4589, w4492, IN29[15], w4590, w4591);
  FullAdder U715 (w4591, w4494, IN30[15], w4592, w4593);
  FullAdder U716 (w4593, w4496, IN31[15], w4594, w4595);
  FullAdder U717 (w4595, w4498, IN32[15], w4596, w4597);
  FullAdder U718 (w4597, w4500, IN33[15], w4598, w4599);
  FullAdder U719 (w4599, w4502, IN34[15], w4600, w4601);
  FullAdder U720 (w4601, w4504, IN35[15], w4602, w4603);
  FullAdder U721 (w4603, w4506, IN36[15], w4604, w4605);
  FullAdder U722 (w4605, w4508, IN37[15], w4606, w4607);
  FullAdder U723 (w4607, w4510, IN38[15], w4608, w4609);
  FullAdder U724 (w4609, w4512, IN39[15], w4610, w4611);
  FullAdder U725 (w4611, w4514, IN40[15], w4612, w4613);
  FullAdder U726 (w4613, w4516, IN41[15], w4614, w4615);
  FullAdder U727 (w4615, w4518, IN42[15], w4616, w4617);
  FullAdder U728 (w4617, w4520, IN43[15], w4618, w4619);
  FullAdder U729 (w4619, w4522, IN44[15], w4620, w4621);
  FullAdder U730 (w4621, w4524, IN45[15], w4622, w4623);
  FullAdder U731 (w4623, w4526, IN46[15], w4624, w4625);
  FullAdder U732 (w4625, w4528, IN47[15], w4626, w4627);
  FullAdder U733 (w4627, w4530, IN48[15], w4628, w4629);
  FullAdder U734 (w4629, w4532, IN49[15], w4630, w4631);
  FullAdder U735 (w4631, w4534, IN50[15], w4632, w4633);
  FullAdder U736 (w4633, w4536, IN51[13], w4634, w4635);
  FullAdder U737 (w4635, w4538, IN52[12], w4636, w4637);
  FullAdder U738 (w4637, w4540, IN53[11], w4638, w4639);
  FullAdder U739 (w4639, w4542, IN54[10], w4640, w4641);
  FullAdder U740 (w4641, w4544, IN55[9], w4642, w4643);
  FullAdder U741 (w4643, w4546, IN56[8], w4644, w4645);
  FullAdder U742 (w4645, w4548, IN57[7], w4646, w4647);
  FullAdder U743 (w4647, w4550, IN58[6], w4648, w4649);
  FullAdder U744 (w4649, w4552, IN59[5], w4650, w4651);
  FullAdder U745 (w4651, w4554, IN60[4], w4652, w4653);
  FullAdder U746 (w4653, w4556, IN61[3], w4654, w4655);
  FullAdder U747 (w4655, w4558, IN62[2], w4656, w4657);
  FullAdder U748 (w4657, w4560, IN63[1], w4658, w4659);
  FullAdder U749 (w4659, w4561, IN64[0], w4660, w4661);
  HalfAdder U750 (w4564, IN16[16], Out1[16], w4663);
  FullAdder U751 (w4663, w4566, IN17[16], w4664, w4665);
  FullAdder U752 (w4665, w4568, IN18[16], w4666, w4667);
  FullAdder U753 (w4667, w4570, IN19[16], w4668, w4669);
  FullAdder U754 (w4669, w4572, IN20[16], w4670, w4671);
  FullAdder U755 (w4671, w4574, IN21[16], w4672, w4673);
  FullAdder U756 (w4673, w4576, IN22[16], w4674, w4675);
  FullAdder U757 (w4675, w4578, IN23[16], w4676, w4677);
  FullAdder U758 (w4677, w4580, IN24[16], w4678, w4679);
  FullAdder U759 (w4679, w4582, IN25[16], w4680, w4681);
  FullAdder U760 (w4681, w4584, IN26[16], w4682, w4683);
  FullAdder U761 (w4683, w4586, IN27[16], w4684, w4685);
  FullAdder U762 (w4685, w4588, IN28[16], w4686, w4687);
  FullAdder U763 (w4687, w4590, IN29[16], w4688, w4689);
  FullAdder U764 (w4689, w4592, IN30[16], w4690, w4691);
  FullAdder U765 (w4691, w4594, IN31[16], w4692, w4693);
  FullAdder U766 (w4693, w4596, IN32[16], w4694, w4695);
  FullAdder U767 (w4695, w4598, IN33[16], w4696, w4697);
  FullAdder U768 (w4697, w4600, IN34[16], w4698, w4699);
  FullAdder U769 (w4699, w4602, IN35[16], w4700, w4701);
  FullAdder U770 (w4701, w4604, IN36[16], w4702, w4703);
  FullAdder U771 (w4703, w4606, IN37[16], w4704, w4705);
  FullAdder U772 (w4705, w4608, IN38[16], w4706, w4707);
  FullAdder U773 (w4707, w4610, IN39[16], w4708, w4709);
  FullAdder U774 (w4709, w4612, IN40[16], w4710, w4711);
  FullAdder U775 (w4711, w4614, IN41[16], w4712, w4713);
  FullAdder U776 (w4713, w4616, IN42[16], w4714, w4715);
  FullAdder U777 (w4715, w4618, IN43[16], w4716, w4717);
  FullAdder U778 (w4717, w4620, IN44[16], w4718, w4719);
  FullAdder U779 (w4719, w4622, IN45[16], w4720, w4721);
  FullAdder U780 (w4721, w4624, IN46[16], w4722, w4723);
  FullAdder U781 (w4723, w4626, IN47[16], w4724, w4725);
  FullAdder U782 (w4725, w4628, IN48[16], w4726, w4727);
  FullAdder U783 (w4727, w4630, IN49[16], w4728, w4729);
  FullAdder U784 (w4729, w4632, IN50[16], w4730, w4731);
  FullAdder U785 (w4731, w4634, IN51[14], w4732, w4733);
  FullAdder U786 (w4733, w4636, IN52[13], w4734, w4735);
  FullAdder U787 (w4735, w4638, IN53[12], w4736, w4737);
  FullAdder U788 (w4737, w4640, IN54[11], w4738, w4739);
  FullAdder U789 (w4739, w4642, IN55[10], w4740, w4741);
  FullAdder U790 (w4741, w4644, IN56[9], w4742, w4743);
  FullAdder U791 (w4743, w4646, IN57[8], w4744, w4745);
  FullAdder U792 (w4745, w4648, IN58[7], w4746, w4747);
  FullAdder U793 (w4747, w4650, IN59[6], w4748, w4749);
  FullAdder U794 (w4749, w4652, IN60[5], w4750, w4751);
  FullAdder U795 (w4751, w4654, IN61[4], w4752, w4753);
  FullAdder U796 (w4753, w4656, IN62[3], w4754, w4755);
  FullAdder U797 (w4755, w4658, IN63[2], w4756, w4757);
  FullAdder U798 (w4757, w4660, IN64[1], w4758, w4759);
  FullAdder U799 (w4759, w4661, IN65[0], w4760, w4761);
  HalfAdder U800 (w4664, IN17[17], Out1[17], w4763);
  FullAdder U801 (w4763, w4666, IN18[17], w4764, w4765);
  FullAdder U802 (w4765, w4668, IN19[17], w4766, w4767);
  FullAdder U803 (w4767, w4670, IN20[17], w4768, w4769);
  FullAdder U804 (w4769, w4672, IN21[17], w4770, w4771);
  FullAdder U805 (w4771, w4674, IN22[17], w4772, w4773);
  FullAdder U806 (w4773, w4676, IN23[17], w4774, w4775);
  FullAdder U807 (w4775, w4678, IN24[17], w4776, w4777);
  FullAdder U808 (w4777, w4680, IN25[17], w4778, w4779);
  FullAdder U809 (w4779, w4682, IN26[17], w4780, w4781);
  FullAdder U810 (w4781, w4684, IN27[17], w4782, w4783);
  FullAdder U811 (w4783, w4686, IN28[17], w4784, w4785);
  FullAdder U812 (w4785, w4688, IN29[17], w4786, w4787);
  FullAdder U813 (w4787, w4690, IN30[17], w4788, w4789);
  FullAdder U814 (w4789, w4692, IN31[17], w4790, w4791);
  FullAdder U815 (w4791, w4694, IN32[17], w4792, w4793);
  FullAdder U816 (w4793, w4696, IN33[17], w4794, w4795);
  FullAdder U817 (w4795, w4698, IN34[17], w4796, w4797);
  FullAdder U818 (w4797, w4700, IN35[17], w4798, w4799);
  FullAdder U819 (w4799, w4702, IN36[17], w4800, w4801);
  FullAdder U820 (w4801, w4704, IN37[17], w4802, w4803);
  FullAdder U821 (w4803, w4706, IN38[17], w4804, w4805);
  FullAdder U822 (w4805, w4708, IN39[17], w4806, w4807);
  FullAdder U823 (w4807, w4710, IN40[17], w4808, w4809);
  FullAdder U824 (w4809, w4712, IN41[17], w4810, w4811);
  FullAdder U825 (w4811, w4714, IN42[17], w4812, w4813);
  FullAdder U826 (w4813, w4716, IN43[17], w4814, w4815);
  FullAdder U827 (w4815, w4718, IN44[17], w4816, w4817);
  FullAdder U828 (w4817, w4720, IN45[17], w4818, w4819);
  FullAdder U829 (w4819, w4722, IN46[17], w4820, w4821);
  FullAdder U830 (w4821, w4724, IN47[17], w4822, w4823);
  FullAdder U831 (w4823, w4726, IN48[17], w4824, w4825);
  FullAdder U832 (w4825, w4728, IN49[17], w4826, w4827);
  FullAdder U833 (w4827, w4730, IN50[17], w4828, w4829);
  FullAdder U834 (w4829, w4732, IN51[15], w4830, w4831);
  FullAdder U835 (w4831, w4734, IN52[14], w4832, w4833);
  FullAdder U836 (w4833, w4736, IN53[13], w4834, w4835);
  FullAdder U837 (w4835, w4738, IN54[12], w4836, w4837);
  FullAdder U838 (w4837, w4740, IN55[11], w4838, w4839);
  FullAdder U839 (w4839, w4742, IN56[10], w4840, w4841);
  FullAdder U840 (w4841, w4744, IN57[9], w4842, w4843);
  FullAdder U841 (w4843, w4746, IN58[8], w4844, w4845);
  FullAdder U842 (w4845, w4748, IN59[7], w4846, w4847);
  FullAdder U843 (w4847, w4750, IN60[6], w4848, w4849);
  FullAdder U844 (w4849, w4752, IN61[5], w4850, w4851);
  FullAdder U845 (w4851, w4754, IN62[4], w4852, w4853);
  FullAdder U846 (w4853, w4756, IN63[3], w4854, w4855);
  FullAdder U847 (w4855, w4758, IN64[2], w4856, w4857);
  FullAdder U848 (w4857, w4760, IN65[1], w4858, w4859);
  FullAdder U849 (w4859, w4761, IN66[0], w4860, w4861);
  HalfAdder U850 (w4764, IN18[18], Out1[18], w4863);
  FullAdder U851 (w4863, w4766, IN19[18], w4864, w4865);
  FullAdder U852 (w4865, w4768, IN20[18], w4866, w4867);
  FullAdder U853 (w4867, w4770, IN21[18], w4868, w4869);
  FullAdder U854 (w4869, w4772, IN22[18], w4870, w4871);
  FullAdder U855 (w4871, w4774, IN23[18], w4872, w4873);
  FullAdder U856 (w4873, w4776, IN24[18], w4874, w4875);
  FullAdder U857 (w4875, w4778, IN25[18], w4876, w4877);
  FullAdder U858 (w4877, w4780, IN26[18], w4878, w4879);
  FullAdder U859 (w4879, w4782, IN27[18], w4880, w4881);
  FullAdder U860 (w4881, w4784, IN28[18], w4882, w4883);
  FullAdder U861 (w4883, w4786, IN29[18], w4884, w4885);
  FullAdder U862 (w4885, w4788, IN30[18], w4886, w4887);
  FullAdder U863 (w4887, w4790, IN31[18], w4888, w4889);
  FullAdder U864 (w4889, w4792, IN32[18], w4890, w4891);
  FullAdder U865 (w4891, w4794, IN33[18], w4892, w4893);
  FullAdder U866 (w4893, w4796, IN34[18], w4894, w4895);
  FullAdder U867 (w4895, w4798, IN35[18], w4896, w4897);
  FullAdder U868 (w4897, w4800, IN36[18], w4898, w4899);
  FullAdder U869 (w4899, w4802, IN37[18], w4900, w4901);
  FullAdder U870 (w4901, w4804, IN38[18], w4902, w4903);
  FullAdder U871 (w4903, w4806, IN39[18], w4904, w4905);
  FullAdder U872 (w4905, w4808, IN40[18], w4906, w4907);
  FullAdder U873 (w4907, w4810, IN41[18], w4908, w4909);
  FullAdder U874 (w4909, w4812, IN42[18], w4910, w4911);
  FullAdder U875 (w4911, w4814, IN43[18], w4912, w4913);
  FullAdder U876 (w4913, w4816, IN44[18], w4914, w4915);
  FullAdder U877 (w4915, w4818, IN45[18], w4916, w4917);
  FullAdder U878 (w4917, w4820, IN46[18], w4918, w4919);
  FullAdder U879 (w4919, w4822, IN47[18], w4920, w4921);
  FullAdder U880 (w4921, w4824, IN48[18], w4922, w4923);
  FullAdder U881 (w4923, w4826, IN49[18], w4924, w4925);
  FullAdder U882 (w4925, w4828, IN50[18], w4926, w4927);
  FullAdder U883 (w4927, w4830, IN51[16], w4928, w4929);
  FullAdder U884 (w4929, w4832, IN52[15], w4930, w4931);
  FullAdder U885 (w4931, w4834, IN53[14], w4932, w4933);
  FullAdder U886 (w4933, w4836, IN54[13], w4934, w4935);
  FullAdder U887 (w4935, w4838, IN55[12], w4936, w4937);
  FullAdder U888 (w4937, w4840, IN56[11], w4938, w4939);
  FullAdder U889 (w4939, w4842, IN57[10], w4940, w4941);
  FullAdder U890 (w4941, w4844, IN58[9], w4942, w4943);
  FullAdder U891 (w4943, w4846, IN59[8], w4944, w4945);
  FullAdder U892 (w4945, w4848, IN60[7], w4946, w4947);
  FullAdder U893 (w4947, w4850, IN61[6], w4948, w4949);
  FullAdder U894 (w4949, w4852, IN62[5], w4950, w4951);
  FullAdder U895 (w4951, w4854, IN63[4], w4952, w4953);
  FullAdder U896 (w4953, w4856, IN64[3], w4954, w4955);
  FullAdder U897 (w4955, w4858, IN65[2], w4956, w4957);
  FullAdder U898 (w4957, w4860, IN66[1], w4958, w4959);
  FullAdder U899 (w4959, w4861, IN67[0], w4960, w4961);
  HalfAdder U900 (w4864, IN19[19], Out1[19], w4963);
  FullAdder U901 (w4963, w4866, IN20[19], w4964, w4965);
  FullAdder U902 (w4965, w4868, IN21[19], w4966, w4967);
  FullAdder U903 (w4967, w4870, IN22[19], w4968, w4969);
  FullAdder U904 (w4969, w4872, IN23[19], w4970, w4971);
  FullAdder U905 (w4971, w4874, IN24[19], w4972, w4973);
  FullAdder U906 (w4973, w4876, IN25[19], w4974, w4975);
  FullAdder U907 (w4975, w4878, IN26[19], w4976, w4977);
  FullAdder U908 (w4977, w4880, IN27[19], w4978, w4979);
  FullAdder U909 (w4979, w4882, IN28[19], w4980, w4981);
  FullAdder U910 (w4981, w4884, IN29[19], w4982, w4983);
  FullAdder U911 (w4983, w4886, IN30[19], w4984, w4985);
  FullAdder U912 (w4985, w4888, IN31[19], w4986, w4987);
  FullAdder U913 (w4987, w4890, IN32[19], w4988, w4989);
  FullAdder U914 (w4989, w4892, IN33[19], w4990, w4991);
  FullAdder U915 (w4991, w4894, IN34[19], w4992, w4993);
  FullAdder U916 (w4993, w4896, IN35[19], w4994, w4995);
  FullAdder U917 (w4995, w4898, IN36[19], w4996, w4997);
  FullAdder U918 (w4997, w4900, IN37[19], w4998, w4999);
  FullAdder U919 (w4999, w4902, IN38[19], w5000, w5001);
  FullAdder U920 (w5001, w4904, IN39[19], w5002, w5003);
  FullAdder U921 (w5003, w4906, IN40[19], w5004, w5005);
  FullAdder U922 (w5005, w4908, IN41[19], w5006, w5007);
  FullAdder U923 (w5007, w4910, IN42[19], w5008, w5009);
  FullAdder U924 (w5009, w4912, IN43[19], w5010, w5011);
  FullAdder U925 (w5011, w4914, IN44[19], w5012, w5013);
  FullAdder U926 (w5013, w4916, IN45[19], w5014, w5015);
  FullAdder U927 (w5015, w4918, IN46[19], w5016, w5017);
  FullAdder U928 (w5017, w4920, IN47[19], w5018, w5019);
  FullAdder U929 (w5019, w4922, IN48[19], w5020, w5021);
  FullAdder U930 (w5021, w4924, IN49[19], w5022, w5023);
  FullAdder U931 (w5023, w4926, IN50[19], w5024, w5025);
  FullAdder U932 (w5025, w4928, IN51[17], w5026, w5027);
  FullAdder U933 (w5027, w4930, IN52[16], w5028, w5029);
  FullAdder U934 (w5029, w4932, IN53[15], w5030, w5031);
  FullAdder U935 (w5031, w4934, IN54[14], w5032, w5033);
  FullAdder U936 (w5033, w4936, IN55[13], w5034, w5035);
  FullAdder U937 (w5035, w4938, IN56[12], w5036, w5037);
  FullAdder U938 (w5037, w4940, IN57[11], w5038, w5039);
  FullAdder U939 (w5039, w4942, IN58[10], w5040, w5041);
  FullAdder U940 (w5041, w4944, IN59[9], w5042, w5043);
  FullAdder U941 (w5043, w4946, IN60[8], w5044, w5045);
  FullAdder U942 (w5045, w4948, IN61[7], w5046, w5047);
  FullAdder U943 (w5047, w4950, IN62[6], w5048, w5049);
  FullAdder U944 (w5049, w4952, IN63[5], w5050, w5051);
  FullAdder U945 (w5051, w4954, IN64[4], w5052, w5053);
  FullAdder U946 (w5053, w4956, IN65[3], w5054, w5055);
  FullAdder U947 (w5055, w4958, IN66[2], w5056, w5057);
  FullAdder U948 (w5057, w4960, IN67[1], w5058, w5059);
  FullAdder U949 (w5059, w4961, IN68[0], w5060, w5061);
  HalfAdder U950 (w4964, IN20[20], Out1[20], w5063);
  FullAdder U951 (w5063, w4966, IN21[20], w5064, w5065);
  FullAdder U952 (w5065, w4968, IN22[20], w5066, w5067);
  FullAdder U953 (w5067, w4970, IN23[20], w5068, w5069);
  FullAdder U954 (w5069, w4972, IN24[20], w5070, w5071);
  FullAdder U955 (w5071, w4974, IN25[20], w5072, w5073);
  FullAdder U956 (w5073, w4976, IN26[20], w5074, w5075);
  FullAdder U957 (w5075, w4978, IN27[20], w5076, w5077);
  FullAdder U958 (w5077, w4980, IN28[20], w5078, w5079);
  FullAdder U959 (w5079, w4982, IN29[20], w5080, w5081);
  FullAdder U960 (w5081, w4984, IN30[20], w5082, w5083);
  FullAdder U961 (w5083, w4986, IN31[20], w5084, w5085);
  FullAdder U962 (w5085, w4988, IN32[20], w5086, w5087);
  FullAdder U963 (w5087, w4990, IN33[20], w5088, w5089);
  FullAdder U964 (w5089, w4992, IN34[20], w5090, w5091);
  FullAdder U965 (w5091, w4994, IN35[20], w5092, w5093);
  FullAdder U966 (w5093, w4996, IN36[20], w5094, w5095);
  FullAdder U967 (w5095, w4998, IN37[20], w5096, w5097);
  FullAdder U968 (w5097, w5000, IN38[20], w5098, w5099);
  FullAdder U969 (w5099, w5002, IN39[20], w5100, w5101);
  FullAdder U970 (w5101, w5004, IN40[20], w5102, w5103);
  FullAdder U971 (w5103, w5006, IN41[20], w5104, w5105);
  FullAdder U972 (w5105, w5008, IN42[20], w5106, w5107);
  FullAdder U973 (w5107, w5010, IN43[20], w5108, w5109);
  FullAdder U974 (w5109, w5012, IN44[20], w5110, w5111);
  FullAdder U975 (w5111, w5014, IN45[20], w5112, w5113);
  FullAdder U976 (w5113, w5016, IN46[20], w5114, w5115);
  FullAdder U977 (w5115, w5018, IN47[20], w5116, w5117);
  FullAdder U978 (w5117, w5020, IN48[20], w5118, w5119);
  FullAdder U979 (w5119, w5022, IN49[20], w5120, w5121);
  FullAdder U980 (w5121, w5024, IN50[20], w5122, w5123);
  FullAdder U981 (w5123, w5026, IN51[18], w5124, w5125);
  FullAdder U982 (w5125, w5028, IN52[17], w5126, w5127);
  FullAdder U983 (w5127, w5030, IN53[16], w5128, w5129);
  FullAdder U984 (w5129, w5032, IN54[15], w5130, w5131);
  FullAdder U985 (w5131, w5034, IN55[14], w5132, w5133);
  FullAdder U986 (w5133, w5036, IN56[13], w5134, w5135);
  FullAdder U987 (w5135, w5038, IN57[12], w5136, w5137);
  FullAdder U988 (w5137, w5040, IN58[11], w5138, w5139);
  FullAdder U989 (w5139, w5042, IN59[10], w5140, w5141);
  FullAdder U990 (w5141, w5044, IN60[9], w5142, w5143);
  FullAdder U991 (w5143, w5046, IN61[8], w5144, w5145);
  FullAdder U992 (w5145, w5048, IN62[7], w5146, w5147);
  FullAdder U993 (w5147, w5050, IN63[6], w5148, w5149);
  FullAdder U994 (w5149, w5052, IN64[5], w5150, w5151);
  FullAdder U995 (w5151, w5054, IN65[4], w5152, w5153);
  FullAdder U996 (w5153, w5056, IN66[3], w5154, w5155);
  FullAdder U997 (w5155, w5058, IN67[2], w5156, w5157);
  FullAdder U998 (w5157, w5060, IN68[1], w5158, w5159);
  FullAdder U999 (w5159, w5061, IN69[0], w5160, w5161);
  HalfAdder U1000 (w5064, IN21[21], Out1[21], w5163);
  FullAdder U1001 (w5163, w5066, IN22[21], w5164, w5165);
  FullAdder U1002 (w5165, w5068, IN23[21], w5166, w5167);
  FullAdder U1003 (w5167, w5070, IN24[21], w5168, w5169);
  FullAdder U1004 (w5169, w5072, IN25[21], w5170, w5171);
  FullAdder U1005 (w5171, w5074, IN26[21], w5172, w5173);
  FullAdder U1006 (w5173, w5076, IN27[21], w5174, w5175);
  FullAdder U1007 (w5175, w5078, IN28[21], w5176, w5177);
  FullAdder U1008 (w5177, w5080, IN29[21], w5178, w5179);
  FullAdder U1009 (w5179, w5082, IN30[21], w5180, w5181);
  FullAdder U1010 (w5181, w5084, IN31[21], w5182, w5183);
  FullAdder U1011 (w5183, w5086, IN32[21], w5184, w5185);
  FullAdder U1012 (w5185, w5088, IN33[21], w5186, w5187);
  FullAdder U1013 (w5187, w5090, IN34[21], w5188, w5189);
  FullAdder U1014 (w5189, w5092, IN35[21], w5190, w5191);
  FullAdder U1015 (w5191, w5094, IN36[21], w5192, w5193);
  FullAdder U1016 (w5193, w5096, IN37[21], w5194, w5195);
  FullAdder U1017 (w5195, w5098, IN38[21], w5196, w5197);
  FullAdder U1018 (w5197, w5100, IN39[21], w5198, w5199);
  FullAdder U1019 (w5199, w5102, IN40[21], w5200, w5201);
  FullAdder U1020 (w5201, w5104, IN41[21], w5202, w5203);
  FullAdder U1021 (w5203, w5106, IN42[21], w5204, w5205);
  FullAdder U1022 (w5205, w5108, IN43[21], w5206, w5207);
  FullAdder U1023 (w5207, w5110, IN44[21], w5208, w5209);
  FullAdder U1024 (w5209, w5112, IN45[21], w5210, w5211);
  FullAdder U1025 (w5211, w5114, IN46[21], w5212, w5213);
  FullAdder U1026 (w5213, w5116, IN47[21], w5214, w5215);
  FullAdder U1027 (w5215, w5118, IN48[21], w5216, w5217);
  FullAdder U1028 (w5217, w5120, IN49[21], w5218, w5219);
  FullAdder U1029 (w5219, w5122, IN50[21], w5220, w5221);
  FullAdder U1030 (w5221, w5124, IN51[19], w5222, w5223);
  FullAdder U1031 (w5223, w5126, IN52[18], w5224, w5225);
  FullAdder U1032 (w5225, w5128, IN53[17], w5226, w5227);
  FullAdder U1033 (w5227, w5130, IN54[16], w5228, w5229);
  FullAdder U1034 (w5229, w5132, IN55[15], w5230, w5231);
  FullAdder U1035 (w5231, w5134, IN56[14], w5232, w5233);
  FullAdder U1036 (w5233, w5136, IN57[13], w5234, w5235);
  FullAdder U1037 (w5235, w5138, IN58[12], w5236, w5237);
  FullAdder U1038 (w5237, w5140, IN59[11], w5238, w5239);
  FullAdder U1039 (w5239, w5142, IN60[10], w5240, w5241);
  FullAdder U1040 (w5241, w5144, IN61[9], w5242, w5243);
  FullAdder U1041 (w5243, w5146, IN62[8], w5244, w5245);
  FullAdder U1042 (w5245, w5148, IN63[7], w5246, w5247);
  FullAdder U1043 (w5247, w5150, IN64[6], w5248, w5249);
  FullAdder U1044 (w5249, w5152, IN65[5], w5250, w5251);
  FullAdder U1045 (w5251, w5154, IN66[4], w5252, w5253);
  FullAdder U1046 (w5253, w5156, IN67[3], w5254, w5255);
  FullAdder U1047 (w5255, w5158, IN68[2], w5256, w5257);
  FullAdder U1048 (w5257, w5160, IN69[1], w5258, w5259);
  FullAdder U1049 (w5259, w5161, IN70[0], w5260, w5261);
  HalfAdder U1050 (w5164, IN22[22], Out1[22], w5263);
  FullAdder U1051 (w5263, w5166, IN23[22], w5264, w5265);
  FullAdder U1052 (w5265, w5168, IN24[22], w5266, w5267);
  FullAdder U1053 (w5267, w5170, IN25[22], w5268, w5269);
  FullAdder U1054 (w5269, w5172, IN26[22], w5270, w5271);
  FullAdder U1055 (w5271, w5174, IN27[22], w5272, w5273);
  FullAdder U1056 (w5273, w5176, IN28[22], w5274, w5275);
  FullAdder U1057 (w5275, w5178, IN29[22], w5276, w5277);
  FullAdder U1058 (w5277, w5180, IN30[22], w5278, w5279);
  FullAdder U1059 (w5279, w5182, IN31[22], w5280, w5281);
  FullAdder U1060 (w5281, w5184, IN32[22], w5282, w5283);
  FullAdder U1061 (w5283, w5186, IN33[22], w5284, w5285);
  FullAdder U1062 (w5285, w5188, IN34[22], w5286, w5287);
  FullAdder U1063 (w5287, w5190, IN35[22], w5288, w5289);
  FullAdder U1064 (w5289, w5192, IN36[22], w5290, w5291);
  FullAdder U1065 (w5291, w5194, IN37[22], w5292, w5293);
  FullAdder U1066 (w5293, w5196, IN38[22], w5294, w5295);
  FullAdder U1067 (w5295, w5198, IN39[22], w5296, w5297);
  FullAdder U1068 (w5297, w5200, IN40[22], w5298, w5299);
  FullAdder U1069 (w5299, w5202, IN41[22], w5300, w5301);
  FullAdder U1070 (w5301, w5204, IN42[22], w5302, w5303);
  FullAdder U1071 (w5303, w5206, IN43[22], w5304, w5305);
  FullAdder U1072 (w5305, w5208, IN44[22], w5306, w5307);
  FullAdder U1073 (w5307, w5210, IN45[22], w5308, w5309);
  FullAdder U1074 (w5309, w5212, IN46[22], w5310, w5311);
  FullAdder U1075 (w5311, w5214, IN47[22], w5312, w5313);
  FullAdder U1076 (w5313, w5216, IN48[22], w5314, w5315);
  FullAdder U1077 (w5315, w5218, IN49[22], w5316, w5317);
  FullAdder U1078 (w5317, w5220, IN50[22], w5318, w5319);
  FullAdder U1079 (w5319, w5222, IN51[20], w5320, w5321);
  FullAdder U1080 (w5321, w5224, IN52[19], w5322, w5323);
  FullAdder U1081 (w5323, w5226, IN53[18], w5324, w5325);
  FullAdder U1082 (w5325, w5228, IN54[17], w5326, w5327);
  FullAdder U1083 (w5327, w5230, IN55[16], w5328, w5329);
  FullAdder U1084 (w5329, w5232, IN56[15], w5330, w5331);
  FullAdder U1085 (w5331, w5234, IN57[14], w5332, w5333);
  FullAdder U1086 (w5333, w5236, IN58[13], w5334, w5335);
  FullAdder U1087 (w5335, w5238, IN59[12], w5336, w5337);
  FullAdder U1088 (w5337, w5240, IN60[11], w5338, w5339);
  FullAdder U1089 (w5339, w5242, IN61[10], w5340, w5341);
  FullAdder U1090 (w5341, w5244, IN62[9], w5342, w5343);
  FullAdder U1091 (w5343, w5246, IN63[8], w5344, w5345);
  FullAdder U1092 (w5345, w5248, IN64[7], w5346, w5347);
  FullAdder U1093 (w5347, w5250, IN65[6], w5348, w5349);
  FullAdder U1094 (w5349, w5252, IN66[5], w5350, w5351);
  FullAdder U1095 (w5351, w5254, IN67[4], w5352, w5353);
  FullAdder U1096 (w5353, w5256, IN68[3], w5354, w5355);
  FullAdder U1097 (w5355, w5258, IN69[2], w5356, w5357);
  FullAdder U1098 (w5357, w5260, IN70[1], w5358, w5359);
  FullAdder U1099 (w5359, w5261, IN71[0], w5360, w5361);
  HalfAdder U1100 (w5264, IN23[23], Out1[23], w5363);
  FullAdder U1101 (w5363, w5266, IN24[23], w5364, w5365);
  FullAdder U1102 (w5365, w5268, IN25[23], w5366, w5367);
  FullAdder U1103 (w5367, w5270, IN26[23], w5368, w5369);
  FullAdder U1104 (w5369, w5272, IN27[23], w5370, w5371);
  FullAdder U1105 (w5371, w5274, IN28[23], w5372, w5373);
  FullAdder U1106 (w5373, w5276, IN29[23], w5374, w5375);
  FullAdder U1107 (w5375, w5278, IN30[23], w5376, w5377);
  FullAdder U1108 (w5377, w5280, IN31[23], w5378, w5379);
  FullAdder U1109 (w5379, w5282, IN32[23], w5380, w5381);
  FullAdder U1110 (w5381, w5284, IN33[23], w5382, w5383);
  FullAdder U1111 (w5383, w5286, IN34[23], w5384, w5385);
  FullAdder U1112 (w5385, w5288, IN35[23], w5386, w5387);
  FullAdder U1113 (w5387, w5290, IN36[23], w5388, w5389);
  FullAdder U1114 (w5389, w5292, IN37[23], w5390, w5391);
  FullAdder U1115 (w5391, w5294, IN38[23], w5392, w5393);
  FullAdder U1116 (w5393, w5296, IN39[23], w5394, w5395);
  FullAdder U1117 (w5395, w5298, IN40[23], w5396, w5397);
  FullAdder U1118 (w5397, w5300, IN41[23], w5398, w5399);
  FullAdder U1119 (w5399, w5302, IN42[23], w5400, w5401);
  FullAdder U1120 (w5401, w5304, IN43[23], w5402, w5403);
  FullAdder U1121 (w5403, w5306, IN44[23], w5404, w5405);
  FullAdder U1122 (w5405, w5308, IN45[23], w5406, w5407);
  FullAdder U1123 (w5407, w5310, IN46[23], w5408, w5409);
  FullAdder U1124 (w5409, w5312, IN47[23], w5410, w5411);
  FullAdder U1125 (w5411, w5314, IN48[23], w5412, w5413);
  FullAdder U1126 (w5413, w5316, IN49[23], w5414, w5415);
  FullAdder U1127 (w5415, w5318, IN50[23], w5416, w5417);
  FullAdder U1128 (w5417, w5320, IN51[21], w5418, w5419);
  FullAdder U1129 (w5419, w5322, IN52[20], w5420, w5421);
  FullAdder U1130 (w5421, w5324, IN53[19], w5422, w5423);
  FullAdder U1131 (w5423, w5326, IN54[18], w5424, w5425);
  FullAdder U1132 (w5425, w5328, IN55[17], w5426, w5427);
  FullAdder U1133 (w5427, w5330, IN56[16], w5428, w5429);
  FullAdder U1134 (w5429, w5332, IN57[15], w5430, w5431);
  FullAdder U1135 (w5431, w5334, IN58[14], w5432, w5433);
  FullAdder U1136 (w5433, w5336, IN59[13], w5434, w5435);
  FullAdder U1137 (w5435, w5338, IN60[12], w5436, w5437);
  FullAdder U1138 (w5437, w5340, IN61[11], w5438, w5439);
  FullAdder U1139 (w5439, w5342, IN62[10], w5440, w5441);
  FullAdder U1140 (w5441, w5344, IN63[9], w5442, w5443);
  FullAdder U1141 (w5443, w5346, IN64[8], w5444, w5445);
  FullAdder U1142 (w5445, w5348, IN65[7], w5446, w5447);
  FullAdder U1143 (w5447, w5350, IN66[6], w5448, w5449);
  FullAdder U1144 (w5449, w5352, IN67[5], w5450, w5451);
  FullAdder U1145 (w5451, w5354, IN68[4], w5452, w5453);
  FullAdder U1146 (w5453, w5356, IN69[3], w5454, w5455);
  FullAdder U1147 (w5455, w5358, IN70[2], w5456, w5457);
  FullAdder U1148 (w5457, w5360, IN71[1], w5458, w5459);
  FullAdder U1149 (w5459, w5361, IN72[0], w5460, w5461);
  HalfAdder U1150 (w5364, IN24[24], Out1[24], w5463);
  FullAdder U1151 (w5463, w5366, IN25[24], w5464, w5465);
  FullAdder U1152 (w5465, w5368, IN26[24], w5466, w5467);
  FullAdder U1153 (w5467, w5370, IN27[24], w5468, w5469);
  FullAdder U1154 (w5469, w5372, IN28[24], w5470, w5471);
  FullAdder U1155 (w5471, w5374, IN29[24], w5472, w5473);
  FullAdder U1156 (w5473, w5376, IN30[24], w5474, w5475);
  FullAdder U1157 (w5475, w5378, IN31[24], w5476, w5477);
  FullAdder U1158 (w5477, w5380, IN32[24], w5478, w5479);
  FullAdder U1159 (w5479, w5382, IN33[24], w5480, w5481);
  FullAdder U1160 (w5481, w5384, IN34[24], w5482, w5483);
  FullAdder U1161 (w5483, w5386, IN35[24], w5484, w5485);
  FullAdder U1162 (w5485, w5388, IN36[24], w5486, w5487);
  FullAdder U1163 (w5487, w5390, IN37[24], w5488, w5489);
  FullAdder U1164 (w5489, w5392, IN38[24], w5490, w5491);
  FullAdder U1165 (w5491, w5394, IN39[24], w5492, w5493);
  FullAdder U1166 (w5493, w5396, IN40[24], w5494, w5495);
  FullAdder U1167 (w5495, w5398, IN41[24], w5496, w5497);
  FullAdder U1168 (w5497, w5400, IN42[24], w5498, w5499);
  FullAdder U1169 (w5499, w5402, IN43[24], w5500, w5501);
  FullAdder U1170 (w5501, w5404, IN44[24], w5502, w5503);
  FullAdder U1171 (w5503, w5406, IN45[24], w5504, w5505);
  FullAdder U1172 (w5505, w5408, IN46[24], w5506, w5507);
  FullAdder U1173 (w5507, w5410, IN47[24], w5508, w5509);
  FullAdder U1174 (w5509, w5412, IN48[24], w5510, w5511);
  FullAdder U1175 (w5511, w5414, IN49[24], w5512, w5513);
  FullAdder U1176 (w5513, w5416, IN50[24], w5514, w5515);
  FullAdder U1177 (w5515, w5418, IN51[22], w5516, w5517);
  FullAdder U1178 (w5517, w5420, IN52[21], w5518, w5519);
  FullAdder U1179 (w5519, w5422, IN53[20], w5520, w5521);
  FullAdder U1180 (w5521, w5424, IN54[19], w5522, w5523);
  FullAdder U1181 (w5523, w5426, IN55[18], w5524, w5525);
  FullAdder U1182 (w5525, w5428, IN56[17], w5526, w5527);
  FullAdder U1183 (w5527, w5430, IN57[16], w5528, w5529);
  FullAdder U1184 (w5529, w5432, IN58[15], w5530, w5531);
  FullAdder U1185 (w5531, w5434, IN59[14], w5532, w5533);
  FullAdder U1186 (w5533, w5436, IN60[13], w5534, w5535);
  FullAdder U1187 (w5535, w5438, IN61[12], w5536, w5537);
  FullAdder U1188 (w5537, w5440, IN62[11], w5538, w5539);
  FullAdder U1189 (w5539, w5442, IN63[10], w5540, w5541);
  FullAdder U1190 (w5541, w5444, IN64[9], w5542, w5543);
  FullAdder U1191 (w5543, w5446, IN65[8], w5544, w5545);
  FullAdder U1192 (w5545, w5448, IN66[7], w5546, w5547);
  FullAdder U1193 (w5547, w5450, IN67[6], w5548, w5549);
  FullAdder U1194 (w5549, w5452, IN68[5], w5550, w5551);
  FullAdder U1195 (w5551, w5454, IN69[4], w5552, w5553);
  FullAdder U1196 (w5553, w5456, IN70[3], w5554, w5555);
  FullAdder U1197 (w5555, w5458, IN71[2], w5556, w5557);
  FullAdder U1198 (w5557, w5460, IN72[1], w5558, w5559);
  FullAdder U1199 (w5559, w5461, IN73[0], w5560, w5561);
  HalfAdder U1200 (w5464, IN25[25], Out1[25], w5563);
  FullAdder U1201 (w5563, w5466, IN26[25], w5564, w5565);
  FullAdder U1202 (w5565, w5468, IN27[25], w5566, w5567);
  FullAdder U1203 (w5567, w5470, IN28[25], w5568, w5569);
  FullAdder U1204 (w5569, w5472, IN29[25], w5570, w5571);
  FullAdder U1205 (w5571, w5474, IN30[25], w5572, w5573);
  FullAdder U1206 (w5573, w5476, IN31[25], w5574, w5575);
  FullAdder U1207 (w5575, w5478, IN32[25], w5576, w5577);
  FullAdder U1208 (w5577, w5480, IN33[25], w5578, w5579);
  FullAdder U1209 (w5579, w5482, IN34[25], w5580, w5581);
  FullAdder U1210 (w5581, w5484, IN35[25], w5582, w5583);
  FullAdder U1211 (w5583, w5486, IN36[25], w5584, w5585);
  FullAdder U1212 (w5585, w5488, IN37[25], w5586, w5587);
  FullAdder U1213 (w5587, w5490, IN38[25], w5588, w5589);
  FullAdder U1214 (w5589, w5492, IN39[25], w5590, w5591);
  FullAdder U1215 (w5591, w5494, IN40[25], w5592, w5593);
  FullAdder U1216 (w5593, w5496, IN41[25], w5594, w5595);
  FullAdder U1217 (w5595, w5498, IN42[25], w5596, w5597);
  FullAdder U1218 (w5597, w5500, IN43[25], w5598, w5599);
  FullAdder U1219 (w5599, w5502, IN44[25], w5600, w5601);
  FullAdder U1220 (w5601, w5504, IN45[25], w5602, w5603);
  FullAdder U1221 (w5603, w5506, IN46[25], w5604, w5605);
  FullAdder U1222 (w5605, w5508, IN47[25], w5606, w5607);
  FullAdder U1223 (w5607, w5510, IN48[25], w5608, w5609);
  FullAdder U1224 (w5609, w5512, IN49[25], w5610, w5611);
  FullAdder U1225 (w5611, w5514, IN50[25], w5612, w5613);
  FullAdder U1226 (w5613, w5516, IN51[23], w5614, w5615);
  FullAdder U1227 (w5615, w5518, IN52[22], w5616, w5617);
  FullAdder U1228 (w5617, w5520, IN53[21], w5618, w5619);
  FullAdder U1229 (w5619, w5522, IN54[20], w5620, w5621);
  FullAdder U1230 (w5621, w5524, IN55[19], w5622, w5623);
  FullAdder U1231 (w5623, w5526, IN56[18], w5624, w5625);
  FullAdder U1232 (w5625, w5528, IN57[17], w5626, w5627);
  FullAdder U1233 (w5627, w5530, IN58[16], w5628, w5629);
  FullAdder U1234 (w5629, w5532, IN59[15], w5630, w5631);
  FullAdder U1235 (w5631, w5534, IN60[14], w5632, w5633);
  FullAdder U1236 (w5633, w5536, IN61[13], w5634, w5635);
  FullAdder U1237 (w5635, w5538, IN62[12], w5636, w5637);
  FullAdder U1238 (w5637, w5540, IN63[11], w5638, w5639);
  FullAdder U1239 (w5639, w5542, IN64[10], w5640, w5641);
  FullAdder U1240 (w5641, w5544, IN65[9], w5642, w5643);
  FullAdder U1241 (w5643, w5546, IN66[8], w5644, w5645);
  FullAdder U1242 (w5645, w5548, IN67[7], w5646, w5647);
  FullAdder U1243 (w5647, w5550, IN68[6], w5648, w5649);
  FullAdder U1244 (w5649, w5552, IN69[5], w5650, w5651);
  FullAdder U1245 (w5651, w5554, IN70[4], w5652, w5653);
  FullAdder U1246 (w5653, w5556, IN71[3], w5654, w5655);
  FullAdder U1247 (w5655, w5558, IN72[2], w5656, w5657);
  FullAdder U1248 (w5657, w5560, IN73[1], w5658, w5659);
  FullAdder U1249 (w5659, w5561, IN74[0], w5660, w5661);
  HalfAdder U1250 (w5564, IN26[26], Out1[26], w5663);
  FullAdder U1251 (w5663, w5566, IN27[26], w5664, w5665);
  FullAdder U1252 (w5665, w5568, IN28[26], w5666, w5667);
  FullAdder U1253 (w5667, w5570, IN29[26], w5668, w5669);
  FullAdder U1254 (w5669, w5572, IN30[26], w5670, w5671);
  FullAdder U1255 (w5671, w5574, IN31[26], w5672, w5673);
  FullAdder U1256 (w5673, w5576, IN32[26], w5674, w5675);
  FullAdder U1257 (w5675, w5578, IN33[26], w5676, w5677);
  FullAdder U1258 (w5677, w5580, IN34[26], w5678, w5679);
  FullAdder U1259 (w5679, w5582, IN35[26], w5680, w5681);
  FullAdder U1260 (w5681, w5584, IN36[26], w5682, w5683);
  FullAdder U1261 (w5683, w5586, IN37[26], w5684, w5685);
  FullAdder U1262 (w5685, w5588, IN38[26], w5686, w5687);
  FullAdder U1263 (w5687, w5590, IN39[26], w5688, w5689);
  FullAdder U1264 (w5689, w5592, IN40[26], w5690, w5691);
  FullAdder U1265 (w5691, w5594, IN41[26], w5692, w5693);
  FullAdder U1266 (w5693, w5596, IN42[26], w5694, w5695);
  FullAdder U1267 (w5695, w5598, IN43[26], w5696, w5697);
  FullAdder U1268 (w5697, w5600, IN44[26], w5698, w5699);
  FullAdder U1269 (w5699, w5602, IN45[26], w5700, w5701);
  FullAdder U1270 (w5701, w5604, IN46[26], w5702, w5703);
  FullAdder U1271 (w5703, w5606, IN47[26], w5704, w5705);
  FullAdder U1272 (w5705, w5608, IN48[26], w5706, w5707);
  FullAdder U1273 (w5707, w5610, IN49[26], w5708, w5709);
  FullAdder U1274 (w5709, w5612, IN50[26], w5710, w5711);
  FullAdder U1275 (w5711, w5614, IN51[24], w5712, w5713);
  FullAdder U1276 (w5713, w5616, IN52[23], w5714, w5715);
  FullAdder U1277 (w5715, w5618, IN53[22], w5716, w5717);
  FullAdder U1278 (w5717, w5620, IN54[21], w5718, w5719);
  FullAdder U1279 (w5719, w5622, IN55[20], w5720, w5721);
  FullAdder U1280 (w5721, w5624, IN56[19], w5722, w5723);
  FullAdder U1281 (w5723, w5626, IN57[18], w5724, w5725);
  FullAdder U1282 (w5725, w5628, IN58[17], w5726, w5727);
  FullAdder U1283 (w5727, w5630, IN59[16], w5728, w5729);
  FullAdder U1284 (w5729, w5632, IN60[15], w5730, w5731);
  FullAdder U1285 (w5731, w5634, IN61[14], w5732, w5733);
  FullAdder U1286 (w5733, w5636, IN62[13], w5734, w5735);
  FullAdder U1287 (w5735, w5638, IN63[12], w5736, w5737);
  FullAdder U1288 (w5737, w5640, IN64[11], w5738, w5739);
  FullAdder U1289 (w5739, w5642, IN65[10], w5740, w5741);
  FullAdder U1290 (w5741, w5644, IN66[9], w5742, w5743);
  FullAdder U1291 (w5743, w5646, IN67[8], w5744, w5745);
  FullAdder U1292 (w5745, w5648, IN68[7], w5746, w5747);
  FullAdder U1293 (w5747, w5650, IN69[6], w5748, w5749);
  FullAdder U1294 (w5749, w5652, IN70[5], w5750, w5751);
  FullAdder U1295 (w5751, w5654, IN71[4], w5752, w5753);
  FullAdder U1296 (w5753, w5656, IN72[3], w5754, w5755);
  FullAdder U1297 (w5755, w5658, IN73[2], w5756, w5757);
  FullAdder U1298 (w5757, w5660, IN74[1], w5758, w5759);
  FullAdder U1299 (w5759, w5661, IN75[0], w5760, w5761);
  HalfAdder U1300 (w5664, IN27[27], Out1[27], w5763);
  FullAdder U1301 (w5763, w5666, IN28[27], w5764, w5765);
  FullAdder U1302 (w5765, w5668, IN29[27], w5766, w5767);
  FullAdder U1303 (w5767, w5670, IN30[27], w5768, w5769);
  FullAdder U1304 (w5769, w5672, IN31[27], w5770, w5771);
  FullAdder U1305 (w5771, w5674, IN32[27], w5772, w5773);
  FullAdder U1306 (w5773, w5676, IN33[27], w5774, w5775);
  FullAdder U1307 (w5775, w5678, IN34[27], w5776, w5777);
  FullAdder U1308 (w5777, w5680, IN35[27], w5778, w5779);
  FullAdder U1309 (w5779, w5682, IN36[27], w5780, w5781);
  FullAdder U1310 (w5781, w5684, IN37[27], w5782, w5783);
  FullAdder U1311 (w5783, w5686, IN38[27], w5784, w5785);
  FullAdder U1312 (w5785, w5688, IN39[27], w5786, w5787);
  FullAdder U1313 (w5787, w5690, IN40[27], w5788, w5789);
  FullAdder U1314 (w5789, w5692, IN41[27], w5790, w5791);
  FullAdder U1315 (w5791, w5694, IN42[27], w5792, w5793);
  FullAdder U1316 (w5793, w5696, IN43[27], w5794, w5795);
  FullAdder U1317 (w5795, w5698, IN44[27], w5796, w5797);
  FullAdder U1318 (w5797, w5700, IN45[27], w5798, w5799);
  FullAdder U1319 (w5799, w5702, IN46[27], w5800, w5801);
  FullAdder U1320 (w5801, w5704, IN47[27], w5802, w5803);
  FullAdder U1321 (w5803, w5706, IN48[27], w5804, w5805);
  FullAdder U1322 (w5805, w5708, IN49[27], w5806, w5807);
  FullAdder U1323 (w5807, w5710, IN50[27], w5808, w5809);
  FullAdder U1324 (w5809, w5712, IN51[25], w5810, w5811);
  FullAdder U1325 (w5811, w5714, IN52[24], w5812, w5813);
  FullAdder U1326 (w5813, w5716, IN53[23], w5814, w5815);
  FullAdder U1327 (w5815, w5718, IN54[22], w5816, w5817);
  FullAdder U1328 (w5817, w5720, IN55[21], w5818, w5819);
  FullAdder U1329 (w5819, w5722, IN56[20], w5820, w5821);
  FullAdder U1330 (w5821, w5724, IN57[19], w5822, w5823);
  FullAdder U1331 (w5823, w5726, IN58[18], w5824, w5825);
  FullAdder U1332 (w5825, w5728, IN59[17], w5826, w5827);
  FullAdder U1333 (w5827, w5730, IN60[16], w5828, w5829);
  FullAdder U1334 (w5829, w5732, IN61[15], w5830, w5831);
  FullAdder U1335 (w5831, w5734, IN62[14], w5832, w5833);
  FullAdder U1336 (w5833, w5736, IN63[13], w5834, w5835);
  FullAdder U1337 (w5835, w5738, IN64[12], w5836, w5837);
  FullAdder U1338 (w5837, w5740, IN65[11], w5838, w5839);
  FullAdder U1339 (w5839, w5742, IN66[10], w5840, w5841);
  FullAdder U1340 (w5841, w5744, IN67[9], w5842, w5843);
  FullAdder U1341 (w5843, w5746, IN68[8], w5844, w5845);
  FullAdder U1342 (w5845, w5748, IN69[7], w5846, w5847);
  FullAdder U1343 (w5847, w5750, IN70[6], w5848, w5849);
  FullAdder U1344 (w5849, w5752, IN71[5], w5850, w5851);
  FullAdder U1345 (w5851, w5754, IN72[4], w5852, w5853);
  FullAdder U1346 (w5853, w5756, IN73[3], w5854, w5855);
  FullAdder U1347 (w5855, w5758, IN74[2], w5856, w5857);
  FullAdder U1348 (w5857, w5760, IN75[1], w5858, w5859);
  FullAdder U1349 (w5859, w5761, IN76[0], w5860, w5861);
  HalfAdder U1350 (w5764, IN28[28], Out1[28], w5863);
  FullAdder U1351 (w5863, w5766, IN29[28], w5864, w5865);
  FullAdder U1352 (w5865, w5768, IN30[28], w5866, w5867);
  FullAdder U1353 (w5867, w5770, IN31[28], w5868, w5869);
  FullAdder U1354 (w5869, w5772, IN32[28], w5870, w5871);
  FullAdder U1355 (w5871, w5774, IN33[28], w5872, w5873);
  FullAdder U1356 (w5873, w5776, IN34[28], w5874, w5875);
  FullAdder U1357 (w5875, w5778, IN35[28], w5876, w5877);
  FullAdder U1358 (w5877, w5780, IN36[28], w5878, w5879);
  FullAdder U1359 (w5879, w5782, IN37[28], w5880, w5881);
  FullAdder U1360 (w5881, w5784, IN38[28], w5882, w5883);
  FullAdder U1361 (w5883, w5786, IN39[28], w5884, w5885);
  FullAdder U1362 (w5885, w5788, IN40[28], w5886, w5887);
  FullAdder U1363 (w5887, w5790, IN41[28], w5888, w5889);
  FullAdder U1364 (w5889, w5792, IN42[28], w5890, w5891);
  FullAdder U1365 (w5891, w5794, IN43[28], w5892, w5893);
  FullAdder U1366 (w5893, w5796, IN44[28], w5894, w5895);
  FullAdder U1367 (w5895, w5798, IN45[28], w5896, w5897);
  FullAdder U1368 (w5897, w5800, IN46[28], w5898, w5899);
  FullAdder U1369 (w5899, w5802, IN47[28], w5900, w5901);
  FullAdder U1370 (w5901, w5804, IN48[28], w5902, w5903);
  FullAdder U1371 (w5903, w5806, IN49[28], w5904, w5905);
  FullAdder U1372 (w5905, w5808, IN50[28], w5906, w5907);
  FullAdder U1373 (w5907, w5810, IN51[26], w5908, w5909);
  FullAdder U1374 (w5909, w5812, IN52[25], w5910, w5911);
  FullAdder U1375 (w5911, w5814, IN53[24], w5912, w5913);
  FullAdder U1376 (w5913, w5816, IN54[23], w5914, w5915);
  FullAdder U1377 (w5915, w5818, IN55[22], w5916, w5917);
  FullAdder U1378 (w5917, w5820, IN56[21], w5918, w5919);
  FullAdder U1379 (w5919, w5822, IN57[20], w5920, w5921);
  FullAdder U1380 (w5921, w5824, IN58[19], w5922, w5923);
  FullAdder U1381 (w5923, w5826, IN59[18], w5924, w5925);
  FullAdder U1382 (w5925, w5828, IN60[17], w5926, w5927);
  FullAdder U1383 (w5927, w5830, IN61[16], w5928, w5929);
  FullAdder U1384 (w5929, w5832, IN62[15], w5930, w5931);
  FullAdder U1385 (w5931, w5834, IN63[14], w5932, w5933);
  FullAdder U1386 (w5933, w5836, IN64[13], w5934, w5935);
  FullAdder U1387 (w5935, w5838, IN65[12], w5936, w5937);
  FullAdder U1388 (w5937, w5840, IN66[11], w5938, w5939);
  FullAdder U1389 (w5939, w5842, IN67[10], w5940, w5941);
  FullAdder U1390 (w5941, w5844, IN68[9], w5942, w5943);
  FullAdder U1391 (w5943, w5846, IN69[8], w5944, w5945);
  FullAdder U1392 (w5945, w5848, IN70[7], w5946, w5947);
  FullAdder U1393 (w5947, w5850, IN71[6], w5948, w5949);
  FullAdder U1394 (w5949, w5852, IN72[5], w5950, w5951);
  FullAdder U1395 (w5951, w5854, IN73[4], w5952, w5953);
  FullAdder U1396 (w5953, w5856, IN74[3], w5954, w5955);
  FullAdder U1397 (w5955, w5858, IN75[2], w5956, w5957);
  FullAdder U1398 (w5957, w5860, IN76[1], w5958, w5959);
  FullAdder U1399 (w5959, w5861, IN77[0], w5960, w5961);
  HalfAdder U1400 (w5864, IN29[29], Out1[29], w5963);
  FullAdder U1401 (w5963, w5866, IN30[29], w5964, w5965);
  FullAdder U1402 (w5965, w5868, IN31[29], w5966, w5967);
  FullAdder U1403 (w5967, w5870, IN32[29], w5968, w5969);
  FullAdder U1404 (w5969, w5872, IN33[29], w5970, w5971);
  FullAdder U1405 (w5971, w5874, IN34[29], w5972, w5973);
  FullAdder U1406 (w5973, w5876, IN35[29], w5974, w5975);
  FullAdder U1407 (w5975, w5878, IN36[29], w5976, w5977);
  FullAdder U1408 (w5977, w5880, IN37[29], w5978, w5979);
  FullAdder U1409 (w5979, w5882, IN38[29], w5980, w5981);
  FullAdder U1410 (w5981, w5884, IN39[29], w5982, w5983);
  FullAdder U1411 (w5983, w5886, IN40[29], w5984, w5985);
  FullAdder U1412 (w5985, w5888, IN41[29], w5986, w5987);
  FullAdder U1413 (w5987, w5890, IN42[29], w5988, w5989);
  FullAdder U1414 (w5989, w5892, IN43[29], w5990, w5991);
  FullAdder U1415 (w5991, w5894, IN44[29], w5992, w5993);
  FullAdder U1416 (w5993, w5896, IN45[29], w5994, w5995);
  FullAdder U1417 (w5995, w5898, IN46[29], w5996, w5997);
  FullAdder U1418 (w5997, w5900, IN47[29], w5998, w5999);
  FullAdder U1419 (w5999, w5902, IN48[29], w6000, w6001);
  FullAdder U1420 (w6001, w5904, IN49[29], w6002, w6003);
  FullAdder U1421 (w6003, w5906, IN50[29], w6004, w6005);
  FullAdder U1422 (w6005, w5908, IN51[27], w6006, w6007);
  FullAdder U1423 (w6007, w5910, IN52[26], w6008, w6009);
  FullAdder U1424 (w6009, w5912, IN53[25], w6010, w6011);
  FullAdder U1425 (w6011, w5914, IN54[24], w6012, w6013);
  FullAdder U1426 (w6013, w5916, IN55[23], w6014, w6015);
  FullAdder U1427 (w6015, w5918, IN56[22], w6016, w6017);
  FullAdder U1428 (w6017, w5920, IN57[21], w6018, w6019);
  FullAdder U1429 (w6019, w5922, IN58[20], w6020, w6021);
  FullAdder U1430 (w6021, w5924, IN59[19], w6022, w6023);
  FullAdder U1431 (w6023, w5926, IN60[18], w6024, w6025);
  FullAdder U1432 (w6025, w5928, IN61[17], w6026, w6027);
  FullAdder U1433 (w6027, w5930, IN62[16], w6028, w6029);
  FullAdder U1434 (w6029, w5932, IN63[15], w6030, w6031);
  FullAdder U1435 (w6031, w5934, IN64[14], w6032, w6033);
  FullAdder U1436 (w6033, w5936, IN65[13], w6034, w6035);
  FullAdder U1437 (w6035, w5938, IN66[12], w6036, w6037);
  FullAdder U1438 (w6037, w5940, IN67[11], w6038, w6039);
  FullAdder U1439 (w6039, w5942, IN68[10], w6040, w6041);
  FullAdder U1440 (w6041, w5944, IN69[9], w6042, w6043);
  FullAdder U1441 (w6043, w5946, IN70[8], w6044, w6045);
  FullAdder U1442 (w6045, w5948, IN71[7], w6046, w6047);
  FullAdder U1443 (w6047, w5950, IN72[6], w6048, w6049);
  FullAdder U1444 (w6049, w5952, IN73[5], w6050, w6051);
  FullAdder U1445 (w6051, w5954, IN74[4], w6052, w6053);
  FullAdder U1446 (w6053, w5956, IN75[3], w6054, w6055);
  FullAdder U1447 (w6055, w5958, IN76[2], w6056, w6057);
  FullAdder U1448 (w6057, w5960, IN77[1], w6058, w6059);
  FullAdder U1449 (w6059, w5961, IN78[0], w6060, w6061);
  HalfAdder U1450 (w5964, IN30[30], Out1[30], w6063);
  FullAdder U1451 (w6063, w5966, IN31[30], w6064, w6065);
  FullAdder U1452 (w6065, w5968, IN32[30], w6066, w6067);
  FullAdder U1453 (w6067, w5970, IN33[30], w6068, w6069);
  FullAdder U1454 (w6069, w5972, IN34[30], w6070, w6071);
  FullAdder U1455 (w6071, w5974, IN35[30], w6072, w6073);
  FullAdder U1456 (w6073, w5976, IN36[30], w6074, w6075);
  FullAdder U1457 (w6075, w5978, IN37[30], w6076, w6077);
  FullAdder U1458 (w6077, w5980, IN38[30], w6078, w6079);
  FullAdder U1459 (w6079, w5982, IN39[30], w6080, w6081);
  FullAdder U1460 (w6081, w5984, IN40[30], w6082, w6083);
  FullAdder U1461 (w6083, w5986, IN41[30], w6084, w6085);
  FullAdder U1462 (w6085, w5988, IN42[30], w6086, w6087);
  FullAdder U1463 (w6087, w5990, IN43[30], w6088, w6089);
  FullAdder U1464 (w6089, w5992, IN44[30], w6090, w6091);
  FullAdder U1465 (w6091, w5994, IN45[30], w6092, w6093);
  FullAdder U1466 (w6093, w5996, IN46[30], w6094, w6095);
  FullAdder U1467 (w6095, w5998, IN47[30], w6096, w6097);
  FullAdder U1468 (w6097, w6000, IN48[30], w6098, w6099);
  FullAdder U1469 (w6099, w6002, IN49[30], w6100, w6101);
  FullAdder U1470 (w6101, w6004, IN50[30], w6102, w6103);
  FullAdder U1471 (w6103, w6006, IN51[28], w6104, w6105);
  FullAdder U1472 (w6105, w6008, IN52[27], w6106, w6107);
  FullAdder U1473 (w6107, w6010, IN53[26], w6108, w6109);
  FullAdder U1474 (w6109, w6012, IN54[25], w6110, w6111);
  FullAdder U1475 (w6111, w6014, IN55[24], w6112, w6113);
  FullAdder U1476 (w6113, w6016, IN56[23], w6114, w6115);
  FullAdder U1477 (w6115, w6018, IN57[22], w6116, w6117);
  FullAdder U1478 (w6117, w6020, IN58[21], w6118, w6119);
  FullAdder U1479 (w6119, w6022, IN59[20], w6120, w6121);
  FullAdder U1480 (w6121, w6024, IN60[19], w6122, w6123);
  FullAdder U1481 (w6123, w6026, IN61[18], w6124, w6125);
  FullAdder U1482 (w6125, w6028, IN62[17], w6126, w6127);
  FullAdder U1483 (w6127, w6030, IN63[16], w6128, w6129);
  FullAdder U1484 (w6129, w6032, IN64[15], w6130, w6131);
  FullAdder U1485 (w6131, w6034, IN65[14], w6132, w6133);
  FullAdder U1486 (w6133, w6036, IN66[13], w6134, w6135);
  FullAdder U1487 (w6135, w6038, IN67[12], w6136, w6137);
  FullAdder U1488 (w6137, w6040, IN68[11], w6138, w6139);
  FullAdder U1489 (w6139, w6042, IN69[10], w6140, w6141);
  FullAdder U1490 (w6141, w6044, IN70[9], w6142, w6143);
  FullAdder U1491 (w6143, w6046, IN71[8], w6144, w6145);
  FullAdder U1492 (w6145, w6048, IN72[7], w6146, w6147);
  FullAdder U1493 (w6147, w6050, IN73[6], w6148, w6149);
  FullAdder U1494 (w6149, w6052, IN74[5], w6150, w6151);
  FullAdder U1495 (w6151, w6054, IN75[4], w6152, w6153);
  FullAdder U1496 (w6153, w6056, IN76[3], w6154, w6155);
  FullAdder U1497 (w6155, w6058, IN77[2], w6156, w6157);
  FullAdder U1498 (w6157, w6060, IN78[1], w6158, w6159);
  FullAdder U1499 (w6159, w6061, IN79[0], w6160, w6161);
  HalfAdder U1500 (w6064, IN31[31], Out1[31], w6163);
  FullAdder U1501 (w6163, w6066, IN32[31], w6164, w6165);
  FullAdder U1502 (w6165, w6068, IN33[31], w6166, w6167);
  FullAdder U1503 (w6167, w6070, IN34[31], w6168, w6169);
  FullAdder U1504 (w6169, w6072, IN35[31], w6170, w6171);
  FullAdder U1505 (w6171, w6074, IN36[31], w6172, w6173);
  FullAdder U1506 (w6173, w6076, IN37[31], w6174, w6175);
  FullAdder U1507 (w6175, w6078, IN38[31], w6176, w6177);
  FullAdder U1508 (w6177, w6080, IN39[31], w6178, w6179);
  FullAdder U1509 (w6179, w6082, IN40[31], w6180, w6181);
  FullAdder U1510 (w6181, w6084, IN41[31], w6182, w6183);
  FullAdder U1511 (w6183, w6086, IN42[31], w6184, w6185);
  FullAdder U1512 (w6185, w6088, IN43[31], w6186, w6187);
  FullAdder U1513 (w6187, w6090, IN44[31], w6188, w6189);
  FullAdder U1514 (w6189, w6092, IN45[31], w6190, w6191);
  FullAdder U1515 (w6191, w6094, IN46[31], w6192, w6193);
  FullAdder U1516 (w6193, w6096, IN47[31], w6194, w6195);
  FullAdder U1517 (w6195, w6098, IN48[31], w6196, w6197);
  FullAdder U1518 (w6197, w6100, IN49[31], w6198, w6199);
  FullAdder U1519 (w6199, w6102, IN50[31], w6200, w6201);
  FullAdder U1520 (w6201, w6104, IN51[29], w6202, w6203);
  FullAdder U1521 (w6203, w6106, IN52[28], w6204, w6205);
  FullAdder U1522 (w6205, w6108, IN53[27], w6206, w6207);
  FullAdder U1523 (w6207, w6110, IN54[26], w6208, w6209);
  FullAdder U1524 (w6209, w6112, IN55[25], w6210, w6211);
  FullAdder U1525 (w6211, w6114, IN56[24], w6212, w6213);
  FullAdder U1526 (w6213, w6116, IN57[23], w6214, w6215);
  FullAdder U1527 (w6215, w6118, IN58[22], w6216, w6217);
  FullAdder U1528 (w6217, w6120, IN59[21], w6218, w6219);
  FullAdder U1529 (w6219, w6122, IN60[20], w6220, w6221);
  FullAdder U1530 (w6221, w6124, IN61[19], w6222, w6223);
  FullAdder U1531 (w6223, w6126, IN62[18], w6224, w6225);
  FullAdder U1532 (w6225, w6128, IN63[17], w6226, w6227);
  FullAdder U1533 (w6227, w6130, IN64[16], w6228, w6229);
  FullAdder U1534 (w6229, w6132, IN65[15], w6230, w6231);
  FullAdder U1535 (w6231, w6134, IN66[14], w6232, w6233);
  FullAdder U1536 (w6233, w6136, IN67[13], w6234, w6235);
  FullAdder U1537 (w6235, w6138, IN68[12], w6236, w6237);
  FullAdder U1538 (w6237, w6140, IN69[11], w6238, w6239);
  FullAdder U1539 (w6239, w6142, IN70[10], w6240, w6241);
  FullAdder U1540 (w6241, w6144, IN71[9], w6242, w6243);
  FullAdder U1541 (w6243, w6146, IN72[8], w6244, w6245);
  FullAdder U1542 (w6245, w6148, IN73[7], w6246, w6247);
  FullAdder U1543 (w6247, w6150, IN74[6], w6248, w6249);
  FullAdder U1544 (w6249, w6152, IN75[5], w6250, w6251);
  FullAdder U1545 (w6251, w6154, IN76[4], w6252, w6253);
  FullAdder U1546 (w6253, w6156, IN77[3], w6254, w6255);
  FullAdder U1547 (w6255, w6158, IN78[2], w6256, w6257);
  FullAdder U1548 (w6257, w6160, IN79[1], w6258, w6259);
  FullAdder U1549 (w6259, w6161, IN80[0], w6260, w6261);
  HalfAdder U1550 (w6164, IN32[32], Out1[32], w6263);
  FullAdder U1551 (w6263, w6166, IN33[32], w6264, w6265);
  FullAdder U1552 (w6265, w6168, IN34[32], w6266, w6267);
  FullAdder U1553 (w6267, w6170, IN35[32], w6268, w6269);
  FullAdder U1554 (w6269, w6172, IN36[32], w6270, w6271);
  FullAdder U1555 (w6271, w6174, IN37[32], w6272, w6273);
  FullAdder U1556 (w6273, w6176, IN38[32], w6274, w6275);
  FullAdder U1557 (w6275, w6178, IN39[32], w6276, w6277);
  FullAdder U1558 (w6277, w6180, IN40[32], w6278, w6279);
  FullAdder U1559 (w6279, w6182, IN41[32], w6280, w6281);
  FullAdder U1560 (w6281, w6184, IN42[32], w6282, w6283);
  FullAdder U1561 (w6283, w6186, IN43[32], w6284, w6285);
  FullAdder U1562 (w6285, w6188, IN44[32], w6286, w6287);
  FullAdder U1563 (w6287, w6190, IN45[32], w6288, w6289);
  FullAdder U1564 (w6289, w6192, IN46[32], w6290, w6291);
  FullAdder U1565 (w6291, w6194, IN47[32], w6292, w6293);
  FullAdder U1566 (w6293, w6196, IN48[32], w6294, w6295);
  FullAdder U1567 (w6295, w6198, IN49[32], w6296, w6297);
  FullAdder U1568 (w6297, w6200, IN50[32], w6298, w6299);
  FullAdder U1569 (w6299, w6202, IN51[30], w6300, w6301);
  FullAdder U1570 (w6301, w6204, IN52[29], w6302, w6303);
  FullAdder U1571 (w6303, w6206, IN53[28], w6304, w6305);
  FullAdder U1572 (w6305, w6208, IN54[27], w6306, w6307);
  FullAdder U1573 (w6307, w6210, IN55[26], w6308, w6309);
  FullAdder U1574 (w6309, w6212, IN56[25], w6310, w6311);
  FullAdder U1575 (w6311, w6214, IN57[24], w6312, w6313);
  FullAdder U1576 (w6313, w6216, IN58[23], w6314, w6315);
  FullAdder U1577 (w6315, w6218, IN59[22], w6316, w6317);
  FullAdder U1578 (w6317, w6220, IN60[21], w6318, w6319);
  FullAdder U1579 (w6319, w6222, IN61[20], w6320, w6321);
  FullAdder U1580 (w6321, w6224, IN62[19], w6322, w6323);
  FullAdder U1581 (w6323, w6226, IN63[18], w6324, w6325);
  FullAdder U1582 (w6325, w6228, IN64[17], w6326, w6327);
  FullAdder U1583 (w6327, w6230, IN65[16], w6328, w6329);
  FullAdder U1584 (w6329, w6232, IN66[15], w6330, w6331);
  FullAdder U1585 (w6331, w6234, IN67[14], w6332, w6333);
  FullAdder U1586 (w6333, w6236, IN68[13], w6334, w6335);
  FullAdder U1587 (w6335, w6238, IN69[12], w6336, w6337);
  FullAdder U1588 (w6337, w6240, IN70[11], w6338, w6339);
  FullAdder U1589 (w6339, w6242, IN71[10], w6340, w6341);
  FullAdder U1590 (w6341, w6244, IN72[9], w6342, w6343);
  FullAdder U1591 (w6343, w6246, IN73[8], w6344, w6345);
  FullAdder U1592 (w6345, w6248, IN74[7], w6346, w6347);
  FullAdder U1593 (w6347, w6250, IN75[6], w6348, w6349);
  FullAdder U1594 (w6349, w6252, IN76[5], w6350, w6351);
  FullAdder U1595 (w6351, w6254, IN77[4], w6352, w6353);
  FullAdder U1596 (w6353, w6256, IN78[3], w6354, w6355);
  FullAdder U1597 (w6355, w6258, IN79[2], w6356, w6357);
  FullAdder U1598 (w6357, w6260, IN80[1], w6358, w6359);
  FullAdder U1599 (w6359, w6261, IN81[0], w6360, w6361);
  HalfAdder U1600 (w6264, IN33[33], Out1[33], w6363);
  FullAdder U1601 (w6363, w6266, IN34[33], w6364, w6365);
  FullAdder U1602 (w6365, w6268, IN35[33], w6366, w6367);
  FullAdder U1603 (w6367, w6270, IN36[33], w6368, w6369);
  FullAdder U1604 (w6369, w6272, IN37[33], w6370, w6371);
  FullAdder U1605 (w6371, w6274, IN38[33], w6372, w6373);
  FullAdder U1606 (w6373, w6276, IN39[33], w6374, w6375);
  FullAdder U1607 (w6375, w6278, IN40[33], w6376, w6377);
  FullAdder U1608 (w6377, w6280, IN41[33], w6378, w6379);
  FullAdder U1609 (w6379, w6282, IN42[33], w6380, w6381);
  FullAdder U1610 (w6381, w6284, IN43[33], w6382, w6383);
  FullAdder U1611 (w6383, w6286, IN44[33], w6384, w6385);
  FullAdder U1612 (w6385, w6288, IN45[33], w6386, w6387);
  FullAdder U1613 (w6387, w6290, IN46[33], w6388, w6389);
  FullAdder U1614 (w6389, w6292, IN47[33], w6390, w6391);
  FullAdder U1615 (w6391, w6294, IN48[33], w6392, w6393);
  FullAdder U1616 (w6393, w6296, IN49[33], w6394, w6395);
  FullAdder U1617 (w6395, w6298, IN50[33], w6396, w6397);
  FullAdder U1618 (w6397, w6300, IN51[31], w6398, w6399);
  FullAdder U1619 (w6399, w6302, IN52[30], w6400, w6401);
  FullAdder U1620 (w6401, w6304, IN53[29], w6402, w6403);
  FullAdder U1621 (w6403, w6306, IN54[28], w6404, w6405);
  FullAdder U1622 (w6405, w6308, IN55[27], w6406, w6407);
  FullAdder U1623 (w6407, w6310, IN56[26], w6408, w6409);
  FullAdder U1624 (w6409, w6312, IN57[25], w6410, w6411);
  FullAdder U1625 (w6411, w6314, IN58[24], w6412, w6413);
  FullAdder U1626 (w6413, w6316, IN59[23], w6414, w6415);
  FullAdder U1627 (w6415, w6318, IN60[22], w6416, w6417);
  FullAdder U1628 (w6417, w6320, IN61[21], w6418, w6419);
  FullAdder U1629 (w6419, w6322, IN62[20], w6420, w6421);
  FullAdder U1630 (w6421, w6324, IN63[19], w6422, w6423);
  FullAdder U1631 (w6423, w6326, IN64[18], w6424, w6425);
  FullAdder U1632 (w6425, w6328, IN65[17], w6426, w6427);
  FullAdder U1633 (w6427, w6330, IN66[16], w6428, w6429);
  FullAdder U1634 (w6429, w6332, IN67[15], w6430, w6431);
  FullAdder U1635 (w6431, w6334, IN68[14], w6432, w6433);
  FullAdder U1636 (w6433, w6336, IN69[13], w6434, w6435);
  FullAdder U1637 (w6435, w6338, IN70[12], w6436, w6437);
  FullAdder U1638 (w6437, w6340, IN71[11], w6438, w6439);
  FullAdder U1639 (w6439, w6342, IN72[10], w6440, w6441);
  FullAdder U1640 (w6441, w6344, IN73[9], w6442, w6443);
  FullAdder U1641 (w6443, w6346, IN74[8], w6444, w6445);
  FullAdder U1642 (w6445, w6348, IN75[7], w6446, w6447);
  FullAdder U1643 (w6447, w6350, IN76[6], w6448, w6449);
  FullAdder U1644 (w6449, w6352, IN77[5], w6450, w6451);
  FullAdder U1645 (w6451, w6354, IN78[4], w6452, w6453);
  FullAdder U1646 (w6453, w6356, IN79[3], w6454, w6455);
  FullAdder U1647 (w6455, w6358, IN80[2], w6456, w6457);
  FullAdder U1648 (w6457, w6360, IN81[1], w6458, w6459);
  FullAdder U1649 (w6459, w6361, IN82[0], w6460, w6461);
  HalfAdder U1650 (w6364, IN34[34], Out1[34], w6463);
  FullAdder U1651 (w6463, w6366, IN35[34], w6464, w6465);
  FullAdder U1652 (w6465, w6368, IN36[34], w6466, w6467);
  FullAdder U1653 (w6467, w6370, IN37[34], w6468, w6469);
  FullAdder U1654 (w6469, w6372, IN38[34], w6470, w6471);
  FullAdder U1655 (w6471, w6374, IN39[34], w6472, w6473);
  FullAdder U1656 (w6473, w6376, IN40[34], w6474, w6475);
  FullAdder U1657 (w6475, w6378, IN41[34], w6476, w6477);
  FullAdder U1658 (w6477, w6380, IN42[34], w6478, w6479);
  FullAdder U1659 (w6479, w6382, IN43[34], w6480, w6481);
  FullAdder U1660 (w6481, w6384, IN44[34], w6482, w6483);
  FullAdder U1661 (w6483, w6386, IN45[34], w6484, w6485);
  FullAdder U1662 (w6485, w6388, IN46[34], w6486, w6487);
  FullAdder U1663 (w6487, w6390, IN47[34], w6488, w6489);
  FullAdder U1664 (w6489, w6392, IN48[34], w6490, w6491);
  FullAdder U1665 (w6491, w6394, IN49[34], w6492, w6493);
  FullAdder U1666 (w6493, w6396, IN50[34], w6494, w6495);
  FullAdder U1667 (w6495, w6398, IN51[32], w6496, w6497);
  FullAdder U1668 (w6497, w6400, IN52[31], w6498, w6499);
  FullAdder U1669 (w6499, w6402, IN53[30], w6500, w6501);
  FullAdder U1670 (w6501, w6404, IN54[29], w6502, w6503);
  FullAdder U1671 (w6503, w6406, IN55[28], w6504, w6505);
  FullAdder U1672 (w6505, w6408, IN56[27], w6506, w6507);
  FullAdder U1673 (w6507, w6410, IN57[26], w6508, w6509);
  FullAdder U1674 (w6509, w6412, IN58[25], w6510, w6511);
  FullAdder U1675 (w6511, w6414, IN59[24], w6512, w6513);
  FullAdder U1676 (w6513, w6416, IN60[23], w6514, w6515);
  FullAdder U1677 (w6515, w6418, IN61[22], w6516, w6517);
  FullAdder U1678 (w6517, w6420, IN62[21], w6518, w6519);
  FullAdder U1679 (w6519, w6422, IN63[20], w6520, w6521);
  FullAdder U1680 (w6521, w6424, IN64[19], w6522, w6523);
  FullAdder U1681 (w6523, w6426, IN65[18], w6524, w6525);
  FullAdder U1682 (w6525, w6428, IN66[17], w6526, w6527);
  FullAdder U1683 (w6527, w6430, IN67[16], w6528, w6529);
  FullAdder U1684 (w6529, w6432, IN68[15], w6530, w6531);
  FullAdder U1685 (w6531, w6434, IN69[14], w6532, w6533);
  FullAdder U1686 (w6533, w6436, IN70[13], w6534, w6535);
  FullAdder U1687 (w6535, w6438, IN71[12], w6536, w6537);
  FullAdder U1688 (w6537, w6440, IN72[11], w6538, w6539);
  FullAdder U1689 (w6539, w6442, IN73[10], w6540, w6541);
  FullAdder U1690 (w6541, w6444, IN74[9], w6542, w6543);
  FullAdder U1691 (w6543, w6446, IN75[8], w6544, w6545);
  FullAdder U1692 (w6545, w6448, IN76[7], w6546, w6547);
  FullAdder U1693 (w6547, w6450, IN77[6], w6548, w6549);
  FullAdder U1694 (w6549, w6452, IN78[5], w6550, w6551);
  FullAdder U1695 (w6551, w6454, IN79[4], w6552, w6553);
  FullAdder U1696 (w6553, w6456, IN80[3], w6554, w6555);
  FullAdder U1697 (w6555, w6458, IN81[2], w6556, w6557);
  FullAdder U1698 (w6557, w6460, IN82[1], w6558, w6559);
  FullAdder U1699 (w6559, w6461, IN83[0], w6560, w6561);
  HalfAdder U1700 (w6464, IN35[35], Out1[35], w6563);
  FullAdder U1701 (w6563, w6466, IN36[35], w6564, w6565);
  FullAdder U1702 (w6565, w6468, IN37[35], w6566, w6567);
  FullAdder U1703 (w6567, w6470, IN38[35], w6568, w6569);
  FullAdder U1704 (w6569, w6472, IN39[35], w6570, w6571);
  FullAdder U1705 (w6571, w6474, IN40[35], w6572, w6573);
  FullAdder U1706 (w6573, w6476, IN41[35], w6574, w6575);
  FullAdder U1707 (w6575, w6478, IN42[35], w6576, w6577);
  FullAdder U1708 (w6577, w6480, IN43[35], w6578, w6579);
  FullAdder U1709 (w6579, w6482, IN44[35], w6580, w6581);
  FullAdder U1710 (w6581, w6484, IN45[35], w6582, w6583);
  FullAdder U1711 (w6583, w6486, IN46[35], w6584, w6585);
  FullAdder U1712 (w6585, w6488, IN47[35], w6586, w6587);
  FullAdder U1713 (w6587, w6490, IN48[35], w6588, w6589);
  FullAdder U1714 (w6589, w6492, IN49[35], w6590, w6591);
  FullAdder U1715 (w6591, w6494, IN50[35], w6592, w6593);
  FullAdder U1716 (w6593, w6496, IN51[33], w6594, w6595);
  FullAdder U1717 (w6595, w6498, IN52[32], w6596, w6597);
  FullAdder U1718 (w6597, w6500, IN53[31], w6598, w6599);
  FullAdder U1719 (w6599, w6502, IN54[30], w6600, w6601);
  FullAdder U1720 (w6601, w6504, IN55[29], w6602, w6603);
  FullAdder U1721 (w6603, w6506, IN56[28], w6604, w6605);
  FullAdder U1722 (w6605, w6508, IN57[27], w6606, w6607);
  FullAdder U1723 (w6607, w6510, IN58[26], w6608, w6609);
  FullAdder U1724 (w6609, w6512, IN59[25], w6610, w6611);
  FullAdder U1725 (w6611, w6514, IN60[24], w6612, w6613);
  FullAdder U1726 (w6613, w6516, IN61[23], w6614, w6615);
  FullAdder U1727 (w6615, w6518, IN62[22], w6616, w6617);
  FullAdder U1728 (w6617, w6520, IN63[21], w6618, w6619);
  FullAdder U1729 (w6619, w6522, IN64[20], w6620, w6621);
  FullAdder U1730 (w6621, w6524, IN65[19], w6622, w6623);
  FullAdder U1731 (w6623, w6526, IN66[18], w6624, w6625);
  FullAdder U1732 (w6625, w6528, IN67[17], w6626, w6627);
  FullAdder U1733 (w6627, w6530, IN68[16], w6628, w6629);
  FullAdder U1734 (w6629, w6532, IN69[15], w6630, w6631);
  FullAdder U1735 (w6631, w6534, IN70[14], w6632, w6633);
  FullAdder U1736 (w6633, w6536, IN71[13], w6634, w6635);
  FullAdder U1737 (w6635, w6538, IN72[12], w6636, w6637);
  FullAdder U1738 (w6637, w6540, IN73[11], w6638, w6639);
  FullAdder U1739 (w6639, w6542, IN74[10], w6640, w6641);
  FullAdder U1740 (w6641, w6544, IN75[9], w6642, w6643);
  FullAdder U1741 (w6643, w6546, IN76[8], w6644, w6645);
  FullAdder U1742 (w6645, w6548, IN77[7], w6646, w6647);
  FullAdder U1743 (w6647, w6550, IN78[6], w6648, w6649);
  FullAdder U1744 (w6649, w6552, IN79[5], w6650, w6651);
  FullAdder U1745 (w6651, w6554, IN80[4], w6652, w6653);
  FullAdder U1746 (w6653, w6556, IN81[3], w6654, w6655);
  FullAdder U1747 (w6655, w6558, IN82[2], w6656, w6657);
  FullAdder U1748 (w6657, w6560, IN83[1], w6658, w6659);
  FullAdder U1749 (w6659, w6561, IN84[0], w6660, w6661);
  HalfAdder U1750 (w6564, IN36[36], Out1[36], w6663);
  FullAdder U1751 (w6663, w6566, IN37[36], w6664, w6665);
  FullAdder U1752 (w6665, w6568, IN38[36], w6666, w6667);
  FullAdder U1753 (w6667, w6570, IN39[36], w6668, w6669);
  FullAdder U1754 (w6669, w6572, IN40[36], w6670, w6671);
  FullAdder U1755 (w6671, w6574, IN41[36], w6672, w6673);
  FullAdder U1756 (w6673, w6576, IN42[36], w6674, w6675);
  FullAdder U1757 (w6675, w6578, IN43[36], w6676, w6677);
  FullAdder U1758 (w6677, w6580, IN44[36], w6678, w6679);
  FullAdder U1759 (w6679, w6582, IN45[36], w6680, w6681);
  FullAdder U1760 (w6681, w6584, IN46[36], w6682, w6683);
  FullAdder U1761 (w6683, w6586, IN47[36], w6684, w6685);
  FullAdder U1762 (w6685, w6588, IN48[36], w6686, w6687);
  FullAdder U1763 (w6687, w6590, IN49[36], w6688, w6689);
  FullAdder U1764 (w6689, w6592, IN50[36], w6690, w6691);
  FullAdder U1765 (w6691, w6594, IN51[34], w6692, w6693);
  FullAdder U1766 (w6693, w6596, IN52[33], w6694, w6695);
  FullAdder U1767 (w6695, w6598, IN53[32], w6696, w6697);
  FullAdder U1768 (w6697, w6600, IN54[31], w6698, w6699);
  FullAdder U1769 (w6699, w6602, IN55[30], w6700, w6701);
  FullAdder U1770 (w6701, w6604, IN56[29], w6702, w6703);
  FullAdder U1771 (w6703, w6606, IN57[28], w6704, w6705);
  FullAdder U1772 (w6705, w6608, IN58[27], w6706, w6707);
  FullAdder U1773 (w6707, w6610, IN59[26], w6708, w6709);
  FullAdder U1774 (w6709, w6612, IN60[25], w6710, w6711);
  FullAdder U1775 (w6711, w6614, IN61[24], w6712, w6713);
  FullAdder U1776 (w6713, w6616, IN62[23], w6714, w6715);
  FullAdder U1777 (w6715, w6618, IN63[22], w6716, w6717);
  FullAdder U1778 (w6717, w6620, IN64[21], w6718, w6719);
  FullAdder U1779 (w6719, w6622, IN65[20], w6720, w6721);
  FullAdder U1780 (w6721, w6624, IN66[19], w6722, w6723);
  FullAdder U1781 (w6723, w6626, IN67[18], w6724, w6725);
  FullAdder U1782 (w6725, w6628, IN68[17], w6726, w6727);
  FullAdder U1783 (w6727, w6630, IN69[16], w6728, w6729);
  FullAdder U1784 (w6729, w6632, IN70[15], w6730, w6731);
  FullAdder U1785 (w6731, w6634, IN71[14], w6732, w6733);
  FullAdder U1786 (w6733, w6636, IN72[13], w6734, w6735);
  FullAdder U1787 (w6735, w6638, IN73[12], w6736, w6737);
  FullAdder U1788 (w6737, w6640, IN74[11], w6738, w6739);
  FullAdder U1789 (w6739, w6642, IN75[10], w6740, w6741);
  FullAdder U1790 (w6741, w6644, IN76[9], w6742, w6743);
  FullAdder U1791 (w6743, w6646, IN77[8], w6744, w6745);
  FullAdder U1792 (w6745, w6648, IN78[7], w6746, w6747);
  FullAdder U1793 (w6747, w6650, IN79[6], w6748, w6749);
  FullAdder U1794 (w6749, w6652, IN80[5], w6750, w6751);
  FullAdder U1795 (w6751, w6654, IN81[4], w6752, w6753);
  FullAdder U1796 (w6753, w6656, IN82[3], w6754, w6755);
  FullAdder U1797 (w6755, w6658, IN83[2], w6756, w6757);
  FullAdder U1798 (w6757, w6660, IN84[1], w6758, w6759);
  FullAdder U1799 (w6759, w6661, IN85[0], w6760, w6761);
  HalfAdder U1800 (w6664, IN37[37], Out1[37], w6763);
  FullAdder U1801 (w6763, w6666, IN38[37], w6764, w6765);
  FullAdder U1802 (w6765, w6668, IN39[37], w6766, w6767);
  FullAdder U1803 (w6767, w6670, IN40[37], w6768, w6769);
  FullAdder U1804 (w6769, w6672, IN41[37], w6770, w6771);
  FullAdder U1805 (w6771, w6674, IN42[37], w6772, w6773);
  FullAdder U1806 (w6773, w6676, IN43[37], w6774, w6775);
  FullAdder U1807 (w6775, w6678, IN44[37], w6776, w6777);
  FullAdder U1808 (w6777, w6680, IN45[37], w6778, w6779);
  FullAdder U1809 (w6779, w6682, IN46[37], w6780, w6781);
  FullAdder U1810 (w6781, w6684, IN47[37], w6782, w6783);
  FullAdder U1811 (w6783, w6686, IN48[37], w6784, w6785);
  FullAdder U1812 (w6785, w6688, IN49[37], w6786, w6787);
  FullAdder U1813 (w6787, w6690, IN50[37], w6788, w6789);
  FullAdder U1814 (w6789, w6692, IN51[35], w6790, w6791);
  FullAdder U1815 (w6791, w6694, IN52[34], w6792, w6793);
  FullAdder U1816 (w6793, w6696, IN53[33], w6794, w6795);
  FullAdder U1817 (w6795, w6698, IN54[32], w6796, w6797);
  FullAdder U1818 (w6797, w6700, IN55[31], w6798, w6799);
  FullAdder U1819 (w6799, w6702, IN56[30], w6800, w6801);
  FullAdder U1820 (w6801, w6704, IN57[29], w6802, w6803);
  FullAdder U1821 (w6803, w6706, IN58[28], w6804, w6805);
  FullAdder U1822 (w6805, w6708, IN59[27], w6806, w6807);
  FullAdder U1823 (w6807, w6710, IN60[26], w6808, w6809);
  FullAdder U1824 (w6809, w6712, IN61[25], w6810, w6811);
  FullAdder U1825 (w6811, w6714, IN62[24], w6812, w6813);
  FullAdder U1826 (w6813, w6716, IN63[23], w6814, w6815);
  FullAdder U1827 (w6815, w6718, IN64[22], w6816, w6817);
  FullAdder U1828 (w6817, w6720, IN65[21], w6818, w6819);
  FullAdder U1829 (w6819, w6722, IN66[20], w6820, w6821);
  FullAdder U1830 (w6821, w6724, IN67[19], w6822, w6823);
  FullAdder U1831 (w6823, w6726, IN68[18], w6824, w6825);
  FullAdder U1832 (w6825, w6728, IN69[17], w6826, w6827);
  FullAdder U1833 (w6827, w6730, IN70[16], w6828, w6829);
  FullAdder U1834 (w6829, w6732, IN71[15], w6830, w6831);
  FullAdder U1835 (w6831, w6734, IN72[14], w6832, w6833);
  FullAdder U1836 (w6833, w6736, IN73[13], w6834, w6835);
  FullAdder U1837 (w6835, w6738, IN74[12], w6836, w6837);
  FullAdder U1838 (w6837, w6740, IN75[11], w6838, w6839);
  FullAdder U1839 (w6839, w6742, IN76[10], w6840, w6841);
  FullAdder U1840 (w6841, w6744, IN77[9], w6842, w6843);
  FullAdder U1841 (w6843, w6746, IN78[8], w6844, w6845);
  FullAdder U1842 (w6845, w6748, IN79[7], w6846, w6847);
  FullAdder U1843 (w6847, w6750, IN80[6], w6848, w6849);
  FullAdder U1844 (w6849, w6752, IN81[5], w6850, w6851);
  FullAdder U1845 (w6851, w6754, IN82[4], w6852, w6853);
  FullAdder U1846 (w6853, w6756, IN83[3], w6854, w6855);
  FullAdder U1847 (w6855, w6758, IN84[2], w6856, w6857);
  FullAdder U1848 (w6857, w6760, IN85[1], w6858, w6859);
  FullAdder U1849 (w6859, w6761, IN86[0], w6860, w6861);
  HalfAdder U1850 (w6764, IN38[38], Out1[38], w6863);
  FullAdder U1851 (w6863, w6766, IN39[38], w6864, w6865);
  FullAdder U1852 (w6865, w6768, IN40[38], w6866, w6867);
  FullAdder U1853 (w6867, w6770, IN41[38], w6868, w6869);
  FullAdder U1854 (w6869, w6772, IN42[38], w6870, w6871);
  FullAdder U1855 (w6871, w6774, IN43[38], w6872, w6873);
  FullAdder U1856 (w6873, w6776, IN44[38], w6874, w6875);
  FullAdder U1857 (w6875, w6778, IN45[38], w6876, w6877);
  FullAdder U1858 (w6877, w6780, IN46[38], w6878, w6879);
  FullAdder U1859 (w6879, w6782, IN47[38], w6880, w6881);
  FullAdder U1860 (w6881, w6784, IN48[38], w6882, w6883);
  FullAdder U1861 (w6883, w6786, IN49[38], w6884, w6885);
  FullAdder U1862 (w6885, w6788, IN50[38], w6886, w6887);
  FullAdder U1863 (w6887, w6790, IN51[36], w6888, w6889);
  FullAdder U1864 (w6889, w6792, IN52[35], w6890, w6891);
  FullAdder U1865 (w6891, w6794, IN53[34], w6892, w6893);
  FullAdder U1866 (w6893, w6796, IN54[33], w6894, w6895);
  FullAdder U1867 (w6895, w6798, IN55[32], w6896, w6897);
  FullAdder U1868 (w6897, w6800, IN56[31], w6898, w6899);
  FullAdder U1869 (w6899, w6802, IN57[30], w6900, w6901);
  FullAdder U1870 (w6901, w6804, IN58[29], w6902, w6903);
  FullAdder U1871 (w6903, w6806, IN59[28], w6904, w6905);
  FullAdder U1872 (w6905, w6808, IN60[27], w6906, w6907);
  FullAdder U1873 (w6907, w6810, IN61[26], w6908, w6909);
  FullAdder U1874 (w6909, w6812, IN62[25], w6910, w6911);
  FullAdder U1875 (w6911, w6814, IN63[24], w6912, w6913);
  FullAdder U1876 (w6913, w6816, IN64[23], w6914, w6915);
  FullAdder U1877 (w6915, w6818, IN65[22], w6916, w6917);
  FullAdder U1878 (w6917, w6820, IN66[21], w6918, w6919);
  FullAdder U1879 (w6919, w6822, IN67[20], w6920, w6921);
  FullAdder U1880 (w6921, w6824, IN68[19], w6922, w6923);
  FullAdder U1881 (w6923, w6826, IN69[18], w6924, w6925);
  FullAdder U1882 (w6925, w6828, IN70[17], w6926, w6927);
  FullAdder U1883 (w6927, w6830, IN71[16], w6928, w6929);
  FullAdder U1884 (w6929, w6832, IN72[15], w6930, w6931);
  FullAdder U1885 (w6931, w6834, IN73[14], w6932, w6933);
  FullAdder U1886 (w6933, w6836, IN74[13], w6934, w6935);
  FullAdder U1887 (w6935, w6838, IN75[12], w6936, w6937);
  FullAdder U1888 (w6937, w6840, IN76[11], w6938, w6939);
  FullAdder U1889 (w6939, w6842, IN77[10], w6940, w6941);
  FullAdder U1890 (w6941, w6844, IN78[9], w6942, w6943);
  FullAdder U1891 (w6943, w6846, IN79[8], w6944, w6945);
  FullAdder U1892 (w6945, w6848, IN80[7], w6946, w6947);
  FullAdder U1893 (w6947, w6850, IN81[6], w6948, w6949);
  FullAdder U1894 (w6949, w6852, IN82[5], w6950, w6951);
  FullAdder U1895 (w6951, w6854, IN83[4], w6952, w6953);
  FullAdder U1896 (w6953, w6856, IN84[3], w6954, w6955);
  FullAdder U1897 (w6955, w6858, IN85[2], w6956, w6957);
  FullAdder U1898 (w6957, w6860, IN86[1], w6958, w6959);
  FullAdder U1899 (w6959, w6861, IN87[0], w6960, w6961);
  HalfAdder U1900 (w6864, IN39[39], Out1[39], w6963);
  FullAdder U1901 (w6963, w6866, IN40[39], w6964, w6965);
  FullAdder U1902 (w6965, w6868, IN41[39], w6966, w6967);
  FullAdder U1903 (w6967, w6870, IN42[39], w6968, w6969);
  FullAdder U1904 (w6969, w6872, IN43[39], w6970, w6971);
  FullAdder U1905 (w6971, w6874, IN44[39], w6972, w6973);
  FullAdder U1906 (w6973, w6876, IN45[39], w6974, w6975);
  FullAdder U1907 (w6975, w6878, IN46[39], w6976, w6977);
  FullAdder U1908 (w6977, w6880, IN47[39], w6978, w6979);
  FullAdder U1909 (w6979, w6882, IN48[39], w6980, w6981);
  FullAdder U1910 (w6981, w6884, IN49[39], w6982, w6983);
  FullAdder U1911 (w6983, w6886, IN50[39], w6984, w6985);
  FullAdder U1912 (w6985, w6888, IN51[37], w6986, w6987);
  FullAdder U1913 (w6987, w6890, IN52[36], w6988, w6989);
  FullAdder U1914 (w6989, w6892, IN53[35], w6990, w6991);
  FullAdder U1915 (w6991, w6894, IN54[34], w6992, w6993);
  FullAdder U1916 (w6993, w6896, IN55[33], w6994, w6995);
  FullAdder U1917 (w6995, w6898, IN56[32], w6996, w6997);
  FullAdder U1918 (w6997, w6900, IN57[31], w6998, w6999);
  FullAdder U1919 (w6999, w6902, IN58[30], w7000, w7001);
  FullAdder U1920 (w7001, w6904, IN59[29], w7002, w7003);
  FullAdder U1921 (w7003, w6906, IN60[28], w7004, w7005);
  FullAdder U1922 (w7005, w6908, IN61[27], w7006, w7007);
  FullAdder U1923 (w7007, w6910, IN62[26], w7008, w7009);
  FullAdder U1924 (w7009, w6912, IN63[25], w7010, w7011);
  FullAdder U1925 (w7011, w6914, IN64[24], w7012, w7013);
  FullAdder U1926 (w7013, w6916, IN65[23], w7014, w7015);
  FullAdder U1927 (w7015, w6918, IN66[22], w7016, w7017);
  FullAdder U1928 (w7017, w6920, IN67[21], w7018, w7019);
  FullAdder U1929 (w7019, w6922, IN68[20], w7020, w7021);
  FullAdder U1930 (w7021, w6924, IN69[19], w7022, w7023);
  FullAdder U1931 (w7023, w6926, IN70[18], w7024, w7025);
  FullAdder U1932 (w7025, w6928, IN71[17], w7026, w7027);
  FullAdder U1933 (w7027, w6930, IN72[16], w7028, w7029);
  FullAdder U1934 (w7029, w6932, IN73[15], w7030, w7031);
  FullAdder U1935 (w7031, w6934, IN74[14], w7032, w7033);
  FullAdder U1936 (w7033, w6936, IN75[13], w7034, w7035);
  FullAdder U1937 (w7035, w6938, IN76[12], w7036, w7037);
  FullAdder U1938 (w7037, w6940, IN77[11], w7038, w7039);
  FullAdder U1939 (w7039, w6942, IN78[10], w7040, w7041);
  FullAdder U1940 (w7041, w6944, IN79[9], w7042, w7043);
  FullAdder U1941 (w7043, w6946, IN80[8], w7044, w7045);
  FullAdder U1942 (w7045, w6948, IN81[7], w7046, w7047);
  FullAdder U1943 (w7047, w6950, IN82[6], w7048, w7049);
  FullAdder U1944 (w7049, w6952, IN83[5], w7050, w7051);
  FullAdder U1945 (w7051, w6954, IN84[4], w7052, w7053);
  FullAdder U1946 (w7053, w6956, IN85[3], w7054, w7055);
  FullAdder U1947 (w7055, w6958, IN86[2], w7056, w7057);
  FullAdder U1948 (w7057, w6960, IN87[1], w7058, w7059);
  FullAdder U1949 (w7059, w6961, IN88[0], w7060, w7061);
  HalfAdder U1950 (w6964, IN40[40], Out1[40], w7063);
  FullAdder U1951 (w7063, w6966, IN41[40], w7064, w7065);
  FullAdder U1952 (w7065, w6968, IN42[40], w7066, w7067);
  FullAdder U1953 (w7067, w6970, IN43[40], w7068, w7069);
  FullAdder U1954 (w7069, w6972, IN44[40], w7070, w7071);
  FullAdder U1955 (w7071, w6974, IN45[40], w7072, w7073);
  FullAdder U1956 (w7073, w6976, IN46[40], w7074, w7075);
  FullAdder U1957 (w7075, w6978, IN47[40], w7076, w7077);
  FullAdder U1958 (w7077, w6980, IN48[40], w7078, w7079);
  FullAdder U1959 (w7079, w6982, IN49[40], w7080, w7081);
  FullAdder U1960 (w7081, w6984, IN50[40], w7082, w7083);
  FullAdder U1961 (w7083, w6986, IN51[38], w7084, w7085);
  FullAdder U1962 (w7085, w6988, IN52[37], w7086, w7087);
  FullAdder U1963 (w7087, w6990, IN53[36], w7088, w7089);
  FullAdder U1964 (w7089, w6992, IN54[35], w7090, w7091);
  FullAdder U1965 (w7091, w6994, IN55[34], w7092, w7093);
  FullAdder U1966 (w7093, w6996, IN56[33], w7094, w7095);
  FullAdder U1967 (w7095, w6998, IN57[32], w7096, w7097);
  FullAdder U1968 (w7097, w7000, IN58[31], w7098, w7099);
  FullAdder U1969 (w7099, w7002, IN59[30], w7100, w7101);
  FullAdder U1970 (w7101, w7004, IN60[29], w7102, w7103);
  FullAdder U1971 (w7103, w7006, IN61[28], w7104, w7105);
  FullAdder U1972 (w7105, w7008, IN62[27], w7106, w7107);
  FullAdder U1973 (w7107, w7010, IN63[26], w7108, w7109);
  FullAdder U1974 (w7109, w7012, IN64[25], w7110, w7111);
  FullAdder U1975 (w7111, w7014, IN65[24], w7112, w7113);
  FullAdder U1976 (w7113, w7016, IN66[23], w7114, w7115);
  FullAdder U1977 (w7115, w7018, IN67[22], w7116, w7117);
  FullAdder U1978 (w7117, w7020, IN68[21], w7118, w7119);
  FullAdder U1979 (w7119, w7022, IN69[20], w7120, w7121);
  FullAdder U1980 (w7121, w7024, IN70[19], w7122, w7123);
  FullAdder U1981 (w7123, w7026, IN71[18], w7124, w7125);
  FullAdder U1982 (w7125, w7028, IN72[17], w7126, w7127);
  FullAdder U1983 (w7127, w7030, IN73[16], w7128, w7129);
  FullAdder U1984 (w7129, w7032, IN74[15], w7130, w7131);
  FullAdder U1985 (w7131, w7034, IN75[14], w7132, w7133);
  FullAdder U1986 (w7133, w7036, IN76[13], w7134, w7135);
  FullAdder U1987 (w7135, w7038, IN77[12], w7136, w7137);
  FullAdder U1988 (w7137, w7040, IN78[11], w7138, w7139);
  FullAdder U1989 (w7139, w7042, IN79[10], w7140, w7141);
  FullAdder U1990 (w7141, w7044, IN80[9], w7142, w7143);
  FullAdder U1991 (w7143, w7046, IN81[8], w7144, w7145);
  FullAdder U1992 (w7145, w7048, IN82[7], w7146, w7147);
  FullAdder U1993 (w7147, w7050, IN83[6], w7148, w7149);
  FullAdder U1994 (w7149, w7052, IN84[5], w7150, w7151);
  FullAdder U1995 (w7151, w7054, IN85[4], w7152, w7153);
  FullAdder U1996 (w7153, w7056, IN86[3], w7154, w7155);
  FullAdder U1997 (w7155, w7058, IN87[2], w7156, w7157);
  FullAdder U1998 (w7157, w7060, IN88[1], w7158, w7159);
  FullAdder U1999 (w7159, w7061, IN89[0], w7160, w7161);
  HalfAdder U2000 (w7064, IN41[41], Out1[41], w7163);
  FullAdder U2001 (w7163, w7066, IN42[41], w7164, w7165);
  FullAdder U2002 (w7165, w7068, IN43[41], w7166, w7167);
  FullAdder U2003 (w7167, w7070, IN44[41], w7168, w7169);
  FullAdder U2004 (w7169, w7072, IN45[41], w7170, w7171);
  FullAdder U2005 (w7171, w7074, IN46[41], w7172, w7173);
  FullAdder U2006 (w7173, w7076, IN47[41], w7174, w7175);
  FullAdder U2007 (w7175, w7078, IN48[41], w7176, w7177);
  FullAdder U2008 (w7177, w7080, IN49[41], w7178, w7179);
  FullAdder U2009 (w7179, w7082, IN50[41], w7180, w7181);
  FullAdder U2010 (w7181, w7084, IN51[39], w7182, w7183);
  FullAdder U2011 (w7183, w7086, IN52[38], w7184, w7185);
  FullAdder U2012 (w7185, w7088, IN53[37], w7186, w7187);
  FullAdder U2013 (w7187, w7090, IN54[36], w7188, w7189);
  FullAdder U2014 (w7189, w7092, IN55[35], w7190, w7191);
  FullAdder U2015 (w7191, w7094, IN56[34], w7192, w7193);
  FullAdder U2016 (w7193, w7096, IN57[33], w7194, w7195);
  FullAdder U2017 (w7195, w7098, IN58[32], w7196, w7197);
  FullAdder U2018 (w7197, w7100, IN59[31], w7198, w7199);
  FullAdder U2019 (w7199, w7102, IN60[30], w7200, w7201);
  FullAdder U2020 (w7201, w7104, IN61[29], w7202, w7203);
  FullAdder U2021 (w7203, w7106, IN62[28], w7204, w7205);
  FullAdder U2022 (w7205, w7108, IN63[27], w7206, w7207);
  FullAdder U2023 (w7207, w7110, IN64[26], w7208, w7209);
  FullAdder U2024 (w7209, w7112, IN65[25], w7210, w7211);
  FullAdder U2025 (w7211, w7114, IN66[24], w7212, w7213);
  FullAdder U2026 (w7213, w7116, IN67[23], w7214, w7215);
  FullAdder U2027 (w7215, w7118, IN68[22], w7216, w7217);
  FullAdder U2028 (w7217, w7120, IN69[21], w7218, w7219);
  FullAdder U2029 (w7219, w7122, IN70[20], w7220, w7221);
  FullAdder U2030 (w7221, w7124, IN71[19], w7222, w7223);
  FullAdder U2031 (w7223, w7126, IN72[18], w7224, w7225);
  FullAdder U2032 (w7225, w7128, IN73[17], w7226, w7227);
  FullAdder U2033 (w7227, w7130, IN74[16], w7228, w7229);
  FullAdder U2034 (w7229, w7132, IN75[15], w7230, w7231);
  FullAdder U2035 (w7231, w7134, IN76[14], w7232, w7233);
  FullAdder U2036 (w7233, w7136, IN77[13], w7234, w7235);
  FullAdder U2037 (w7235, w7138, IN78[12], w7236, w7237);
  FullAdder U2038 (w7237, w7140, IN79[11], w7238, w7239);
  FullAdder U2039 (w7239, w7142, IN80[10], w7240, w7241);
  FullAdder U2040 (w7241, w7144, IN81[9], w7242, w7243);
  FullAdder U2041 (w7243, w7146, IN82[8], w7244, w7245);
  FullAdder U2042 (w7245, w7148, IN83[7], w7246, w7247);
  FullAdder U2043 (w7247, w7150, IN84[6], w7248, w7249);
  FullAdder U2044 (w7249, w7152, IN85[5], w7250, w7251);
  FullAdder U2045 (w7251, w7154, IN86[4], w7252, w7253);
  FullAdder U2046 (w7253, w7156, IN87[3], w7254, w7255);
  FullAdder U2047 (w7255, w7158, IN88[2], w7256, w7257);
  FullAdder U2048 (w7257, w7160, IN89[1], w7258, w7259);
  FullAdder U2049 (w7259, w7161, IN90[0], w7260, w7261);
  HalfAdder U2050 (w7164, IN42[42], Out1[42], w7263);
  FullAdder U2051 (w7263, w7166, IN43[42], w7264, w7265);
  FullAdder U2052 (w7265, w7168, IN44[42], w7266, w7267);
  FullAdder U2053 (w7267, w7170, IN45[42], w7268, w7269);
  FullAdder U2054 (w7269, w7172, IN46[42], w7270, w7271);
  FullAdder U2055 (w7271, w7174, IN47[42], w7272, w7273);
  FullAdder U2056 (w7273, w7176, IN48[42], w7274, w7275);
  FullAdder U2057 (w7275, w7178, IN49[42], w7276, w7277);
  FullAdder U2058 (w7277, w7180, IN50[42], w7278, w7279);
  FullAdder U2059 (w7279, w7182, IN51[40], w7280, w7281);
  FullAdder U2060 (w7281, w7184, IN52[39], w7282, w7283);
  FullAdder U2061 (w7283, w7186, IN53[38], w7284, w7285);
  FullAdder U2062 (w7285, w7188, IN54[37], w7286, w7287);
  FullAdder U2063 (w7287, w7190, IN55[36], w7288, w7289);
  FullAdder U2064 (w7289, w7192, IN56[35], w7290, w7291);
  FullAdder U2065 (w7291, w7194, IN57[34], w7292, w7293);
  FullAdder U2066 (w7293, w7196, IN58[33], w7294, w7295);
  FullAdder U2067 (w7295, w7198, IN59[32], w7296, w7297);
  FullAdder U2068 (w7297, w7200, IN60[31], w7298, w7299);
  FullAdder U2069 (w7299, w7202, IN61[30], w7300, w7301);
  FullAdder U2070 (w7301, w7204, IN62[29], w7302, w7303);
  FullAdder U2071 (w7303, w7206, IN63[28], w7304, w7305);
  FullAdder U2072 (w7305, w7208, IN64[27], w7306, w7307);
  FullAdder U2073 (w7307, w7210, IN65[26], w7308, w7309);
  FullAdder U2074 (w7309, w7212, IN66[25], w7310, w7311);
  FullAdder U2075 (w7311, w7214, IN67[24], w7312, w7313);
  FullAdder U2076 (w7313, w7216, IN68[23], w7314, w7315);
  FullAdder U2077 (w7315, w7218, IN69[22], w7316, w7317);
  FullAdder U2078 (w7317, w7220, IN70[21], w7318, w7319);
  FullAdder U2079 (w7319, w7222, IN71[20], w7320, w7321);
  FullAdder U2080 (w7321, w7224, IN72[19], w7322, w7323);
  FullAdder U2081 (w7323, w7226, IN73[18], w7324, w7325);
  FullAdder U2082 (w7325, w7228, IN74[17], w7326, w7327);
  FullAdder U2083 (w7327, w7230, IN75[16], w7328, w7329);
  FullAdder U2084 (w7329, w7232, IN76[15], w7330, w7331);
  FullAdder U2085 (w7331, w7234, IN77[14], w7332, w7333);
  FullAdder U2086 (w7333, w7236, IN78[13], w7334, w7335);
  FullAdder U2087 (w7335, w7238, IN79[12], w7336, w7337);
  FullAdder U2088 (w7337, w7240, IN80[11], w7338, w7339);
  FullAdder U2089 (w7339, w7242, IN81[10], w7340, w7341);
  FullAdder U2090 (w7341, w7244, IN82[9], w7342, w7343);
  FullAdder U2091 (w7343, w7246, IN83[8], w7344, w7345);
  FullAdder U2092 (w7345, w7248, IN84[7], w7346, w7347);
  FullAdder U2093 (w7347, w7250, IN85[6], w7348, w7349);
  FullAdder U2094 (w7349, w7252, IN86[5], w7350, w7351);
  FullAdder U2095 (w7351, w7254, IN87[4], w7352, w7353);
  FullAdder U2096 (w7353, w7256, IN88[3], w7354, w7355);
  FullAdder U2097 (w7355, w7258, IN89[2], w7356, w7357);
  FullAdder U2098 (w7357, w7260, IN90[1], w7358, w7359);
  FullAdder U2099 (w7359, w7261, IN91[0], w7360, w7361);
  HalfAdder U2100 (w7264, IN43[43], Out1[43], w7363);
  FullAdder U2101 (w7363, w7266, IN44[43], w7364, w7365);
  FullAdder U2102 (w7365, w7268, IN45[43], w7366, w7367);
  FullAdder U2103 (w7367, w7270, IN46[43], w7368, w7369);
  FullAdder U2104 (w7369, w7272, IN47[43], w7370, w7371);
  FullAdder U2105 (w7371, w7274, IN48[43], w7372, w7373);
  FullAdder U2106 (w7373, w7276, IN49[43], w7374, w7375);
  FullAdder U2107 (w7375, w7278, IN50[43], w7376, w7377);
  FullAdder U2108 (w7377, w7280, IN51[41], w7378, w7379);
  FullAdder U2109 (w7379, w7282, IN52[40], w7380, w7381);
  FullAdder U2110 (w7381, w7284, IN53[39], w7382, w7383);
  FullAdder U2111 (w7383, w7286, IN54[38], w7384, w7385);
  FullAdder U2112 (w7385, w7288, IN55[37], w7386, w7387);
  FullAdder U2113 (w7387, w7290, IN56[36], w7388, w7389);
  FullAdder U2114 (w7389, w7292, IN57[35], w7390, w7391);
  FullAdder U2115 (w7391, w7294, IN58[34], w7392, w7393);
  FullAdder U2116 (w7393, w7296, IN59[33], w7394, w7395);
  FullAdder U2117 (w7395, w7298, IN60[32], w7396, w7397);
  FullAdder U2118 (w7397, w7300, IN61[31], w7398, w7399);
  FullAdder U2119 (w7399, w7302, IN62[30], w7400, w7401);
  FullAdder U2120 (w7401, w7304, IN63[29], w7402, w7403);
  FullAdder U2121 (w7403, w7306, IN64[28], w7404, w7405);
  FullAdder U2122 (w7405, w7308, IN65[27], w7406, w7407);
  FullAdder U2123 (w7407, w7310, IN66[26], w7408, w7409);
  FullAdder U2124 (w7409, w7312, IN67[25], w7410, w7411);
  FullAdder U2125 (w7411, w7314, IN68[24], w7412, w7413);
  FullAdder U2126 (w7413, w7316, IN69[23], w7414, w7415);
  FullAdder U2127 (w7415, w7318, IN70[22], w7416, w7417);
  FullAdder U2128 (w7417, w7320, IN71[21], w7418, w7419);
  FullAdder U2129 (w7419, w7322, IN72[20], w7420, w7421);
  FullAdder U2130 (w7421, w7324, IN73[19], w7422, w7423);
  FullAdder U2131 (w7423, w7326, IN74[18], w7424, w7425);
  FullAdder U2132 (w7425, w7328, IN75[17], w7426, w7427);
  FullAdder U2133 (w7427, w7330, IN76[16], w7428, w7429);
  FullAdder U2134 (w7429, w7332, IN77[15], w7430, w7431);
  FullAdder U2135 (w7431, w7334, IN78[14], w7432, w7433);
  FullAdder U2136 (w7433, w7336, IN79[13], w7434, w7435);
  FullAdder U2137 (w7435, w7338, IN80[12], w7436, w7437);
  FullAdder U2138 (w7437, w7340, IN81[11], w7438, w7439);
  FullAdder U2139 (w7439, w7342, IN82[10], w7440, w7441);
  FullAdder U2140 (w7441, w7344, IN83[9], w7442, w7443);
  FullAdder U2141 (w7443, w7346, IN84[8], w7444, w7445);
  FullAdder U2142 (w7445, w7348, IN85[7], w7446, w7447);
  FullAdder U2143 (w7447, w7350, IN86[6], w7448, w7449);
  FullAdder U2144 (w7449, w7352, IN87[5], w7450, w7451);
  FullAdder U2145 (w7451, w7354, IN88[4], w7452, w7453);
  FullAdder U2146 (w7453, w7356, IN89[3], w7454, w7455);
  FullAdder U2147 (w7455, w7358, IN90[2], w7456, w7457);
  FullAdder U2148 (w7457, w7360, IN91[1], w7458, w7459);
  FullAdder U2149 (w7459, w7361, IN92[0], w7460, w7461);
  HalfAdder U2150 (w7364, IN44[44], Out1[44], w7463);
  FullAdder U2151 (w7463, w7366, IN45[44], w7464, w7465);
  FullAdder U2152 (w7465, w7368, IN46[44], w7466, w7467);
  FullAdder U2153 (w7467, w7370, IN47[44], w7468, w7469);
  FullAdder U2154 (w7469, w7372, IN48[44], w7470, w7471);
  FullAdder U2155 (w7471, w7374, IN49[44], w7472, w7473);
  FullAdder U2156 (w7473, w7376, IN50[44], w7474, w7475);
  FullAdder U2157 (w7475, w7378, IN51[42], w7476, w7477);
  FullAdder U2158 (w7477, w7380, IN52[41], w7478, w7479);
  FullAdder U2159 (w7479, w7382, IN53[40], w7480, w7481);
  FullAdder U2160 (w7481, w7384, IN54[39], w7482, w7483);
  FullAdder U2161 (w7483, w7386, IN55[38], w7484, w7485);
  FullAdder U2162 (w7485, w7388, IN56[37], w7486, w7487);
  FullAdder U2163 (w7487, w7390, IN57[36], w7488, w7489);
  FullAdder U2164 (w7489, w7392, IN58[35], w7490, w7491);
  FullAdder U2165 (w7491, w7394, IN59[34], w7492, w7493);
  FullAdder U2166 (w7493, w7396, IN60[33], w7494, w7495);
  FullAdder U2167 (w7495, w7398, IN61[32], w7496, w7497);
  FullAdder U2168 (w7497, w7400, IN62[31], w7498, w7499);
  FullAdder U2169 (w7499, w7402, IN63[30], w7500, w7501);
  FullAdder U2170 (w7501, w7404, IN64[29], w7502, w7503);
  FullAdder U2171 (w7503, w7406, IN65[28], w7504, w7505);
  FullAdder U2172 (w7505, w7408, IN66[27], w7506, w7507);
  FullAdder U2173 (w7507, w7410, IN67[26], w7508, w7509);
  FullAdder U2174 (w7509, w7412, IN68[25], w7510, w7511);
  FullAdder U2175 (w7511, w7414, IN69[24], w7512, w7513);
  FullAdder U2176 (w7513, w7416, IN70[23], w7514, w7515);
  FullAdder U2177 (w7515, w7418, IN71[22], w7516, w7517);
  FullAdder U2178 (w7517, w7420, IN72[21], w7518, w7519);
  FullAdder U2179 (w7519, w7422, IN73[20], w7520, w7521);
  FullAdder U2180 (w7521, w7424, IN74[19], w7522, w7523);
  FullAdder U2181 (w7523, w7426, IN75[18], w7524, w7525);
  FullAdder U2182 (w7525, w7428, IN76[17], w7526, w7527);
  FullAdder U2183 (w7527, w7430, IN77[16], w7528, w7529);
  FullAdder U2184 (w7529, w7432, IN78[15], w7530, w7531);
  FullAdder U2185 (w7531, w7434, IN79[14], w7532, w7533);
  FullAdder U2186 (w7533, w7436, IN80[13], w7534, w7535);
  FullAdder U2187 (w7535, w7438, IN81[12], w7536, w7537);
  FullAdder U2188 (w7537, w7440, IN82[11], w7538, w7539);
  FullAdder U2189 (w7539, w7442, IN83[10], w7540, w7541);
  FullAdder U2190 (w7541, w7444, IN84[9], w7542, w7543);
  FullAdder U2191 (w7543, w7446, IN85[8], w7544, w7545);
  FullAdder U2192 (w7545, w7448, IN86[7], w7546, w7547);
  FullAdder U2193 (w7547, w7450, IN87[6], w7548, w7549);
  FullAdder U2194 (w7549, w7452, IN88[5], w7550, w7551);
  FullAdder U2195 (w7551, w7454, IN89[4], w7552, w7553);
  FullAdder U2196 (w7553, w7456, IN90[3], w7554, w7555);
  FullAdder U2197 (w7555, w7458, IN91[2], w7556, w7557);
  FullAdder U2198 (w7557, w7460, IN92[1], w7558, w7559);
  FullAdder U2199 (w7559, w7461, IN93[0], w7560, w7561);
  HalfAdder U2200 (w7464, IN45[45], Out1[45], w7563);
  FullAdder U2201 (w7563, w7466, IN46[45], w7564, w7565);
  FullAdder U2202 (w7565, w7468, IN47[45], w7566, w7567);
  FullAdder U2203 (w7567, w7470, IN48[45], w7568, w7569);
  FullAdder U2204 (w7569, w7472, IN49[45], w7570, w7571);
  FullAdder U2205 (w7571, w7474, IN50[45], w7572, w7573);
  FullAdder U2206 (w7573, w7476, IN51[43], w7574, w7575);
  FullAdder U2207 (w7575, w7478, IN52[42], w7576, w7577);
  FullAdder U2208 (w7577, w7480, IN53[41], w7578, w7579);
  FullAdder U2209 (w7579, w7482, IN54[40], w7580, w7581);
  FullAdder U2210 (w7581, w7484, IN55[39], w7582, w7583);
  FullAdder U2211 (w7583, w7486, IN56[38], w7584, w7585);
  FullAdder U2212 (w7585, w7488, IN57[37], w7586, w7587);
  FullAdder U2213 (w7587, w7490, IN58[36], w7588, w7589);
  FullAdder U2214 (w7589, w7492, IN59[35], w7590, w7591);
  FullAdder U2215 (w7591, w7494, IN60[34], w7592, w7593);
  FullAdder U2216 (w7593, w7496, IN61[33], w7594, w7595);
  FullAdder U2217 (w7595, w7498, IN62[32], w7596, w7597);
  FullAdder U2218 (w7597, w7500, IN63[31], w7598, w7599);
  FullAdder U2219 (w7599, w7502, IN64[30], w7600, w7601);
  FullAdder U2220 (w7601, w7504, IN65[29], w7602, w7603);
  FullAdder U2221 (w7603, w7506, IN66[28], w7604, w7605);
  FullAdder U2222 (w7605, w7508, IN67[27], w7606, w7607);
  FullAdder U2223 (w7607, w7510, IN68[26], w7608, w7609);
  FullAdder U2224 (w7609, w7512, IN69[25], w7610, w7611);
  FullAdder U2225 (w7611, w7514, IN70[24], w7612, w7613);
  FullAdder U2226 (w7613, w7516, IN71[23], w7614, w7615);
  FullAdder U2227 (w7615, w7518, IN72[22], w7616, w7617);
  FullAdder U2228 (w7617, w7520, IN73[21], w7618, w7619);
  FullAdder U2229 (w7619, w7522, IN74[20], w7620, w7621);
  FullAdder U2230 (w7621, w7524, IN75[19], w7622, w7623);
  FullAdder U2231 (w7623, w7526, IN76[18], w7624, w7625);
  FullAdder U2232 (w7625, w7528, IN77[17], w7626, w7627);
  FullAdder U2233 (w7627, w7530, IN78[16], w7628, w7629);
  FullAdder U2234 (w7629, w7532, IN79[15], w7630, w7631);
  FullAdder U2235 (w7631, w7534, IN80[14], w7632, w7633);
  FullAdder U2236 (w7633, w7536, IN81[13], w7634, w7635);
  FullAdder U2237 (w7635, w7538, IN82[12], w7636, w7637);
  FullAdder U2238 (w7637, w7540, IN83[11], w7638, w7639);
  FullAdder U2239 (w7639, w7542, IN84[10], w7640, w7641);
  FullAdder U2240 (w7641, w7544, IN85[9], w7642, w7643);
  FullAdder U2241 (w7643, w7546, IN86[8], w7644, w7645);
  FullAdder U2242 (w7645, w7548, IN87[7], w7646, w7647);
  FullAdder U2243 (w7647, w7550, IN88[6], w7648, w7649);
  FullAdder U2244 (w7649, w7552, IN89[5], w7650, w7651);
  FullAdder U2245 (w7651, w7554, IN90[4], w7652, w7653);
  FullAdder U2246 (w7653, w7556, IN91[3], w7654, w7655);
  FullAdder U2247 (w7655, w7558, IN92[2], w7656, w7657);
  FullAdder U2248 (w7657, w7560, IN93[1], w7658, w7659);
  FullAdder U2249 (w7659, w7561, IN94[0], w7660, w7661);
  HalfAdder U2250 (w7564, IN46[46], Out1[46], w7663);
  FullAdder U2251 (w7663, w7566, IN47[46], w7664, w7665);
  FullAdder U2252 (w7665, w7568, IN48[46], w7666, w7667);
  FullAdder U2253 (w7667, w7570, IN49[46], w7668, w7669);
  FullAdder U2254 (w7669, w7572, IN50[46], w7670, w7671);
  FullAdder U2255 (w7671, w7574, IN51[44], w7672, w7673);
  FullAdder U2256 (w7673, w7576, IN52[43], w7674, w7675);
  FullAdder U2257 (w7675, w7578, IN53[42], w7676, w7677);
  FullAdder U2258 (w7677, w7580, IN54[41], w7678, w7679);
  FullAdder U2259 (w7679, w7582, IN55[40], w7680, w7681);
  FullAdder U2260 (w7681, w7584, IN56[39], w7682, w7683);
  FullAdder U2261 (w7683, w7586, IN57[38], w7684, w7685);
  FullAdder U2262 (w7685, w7588, IN58[37], w7686, w7687);
  FullAdder U2263 (w7687, w7590, IN59[36], w7688, w7689);
  FullAdder U2264 (w7689, w7592, IN60[35], w7690, w7691);
  FullAdder U2265 (w7691, w7594, IN61[34], w7692, w7693);
  FullAdder U2266 (w7693, w7596, IN62[33], w7694, w7695);
  FullAdder U2267 (w7695, w7598, IN63[32], w7696, w7697);
  FullAdder U2268 (w7697, w7600, IN64[31], w7698, w7699);
  FullAdder U2269 (w7699, w7602, IN65[30], w7700, w7701);
  FullAdder U2270 (w7701, w7604, IN66[29], w7702, w7703);
  FullAdder U2271 (w7703, w7606, IN67[28], w7704, w7705);
  FullAdder U2272 (w7705, w7608, IN68[27], w7706, w7707);
  FullAdder U2273 (w7707, w7610, IN69[26], w7708, w7709);
  FullAdder U2274 (w7709, w7612, IN70[25], w7710, w7711);
  FullAdder U2275 (w7711, w7614, IN71[24], w7712, w7713);
  FullAdder U2276 (w7713, w7616, IN72[23], w7714, w7715);
  FullAdder U2277 (w7715, w7618, IN73[22], w7716, w7717);
  FullAdder U2278 (w7717, w7620, IN74[21], w7718, w7719);
  FullAdder U2279 (w7719, w7622, IN75[20], w7720, w7721);
  FullAdder U2280 (w7721, w7624, IN76[19], w7722, w7723);
  FullAdder U2281 (w7723, w7626, IN77[18], w7724, w7725);
  FullAdder U2282 (w7725, w7628, IN78[17], w7726, w7727);
  FullAdder U2283 (w7727, w7630, IN79[16], w7728, w7729);
  FullAdder U2284 (w7729, w7632, IN80[15], w7730, w7731);
  FullAdder U2285 (w7731, w7634, IN81[14], w7732, w7733);
  FullAdder U2286 (w7733, w7636, IN82[13], w7734, w7735);
  FullAdder U2287 (w7735, w7638, IN83[12], w7736, w7737);
  FullAdder U2288 (w7737, w7640, IN84[11], w7738, w7739);
  FullAdder U2289 (w7739, w7642, IN85[10], w7740, w7741);
  FullAdder U2290 (w7741, w7644, IN86[9], w7742, w7743);
  FullAdder U2291 (w7743, w7646, IN87[8], w7744, w7745);
  FullAdder U2292 (w7745, w7648, IN88[7], w7746, w7747);
  FullAdder U2293 (w7747, w7650, IN89[6], w7748, w7749);
  FullAdder U2294 (w7749, w7652, IN90[5], w7750, w7751);
  FullAdder U2295 (w7751, w7654, IN91[4], w7752, w7753);
  FullAdder U2296 (w7753, w7656, IN92[3], w7754, w7755);
  FullAdder U2297 (w7755, w7658, IN93[2], w7756, w7757);
  FullAdder U2298 (w7757, w7660, IN94[1], w7758, w7759);
  FullAdder U2299 (w7759, w7661, IN95[0], w7760, w7761);
  HalfAdder U2300 (w7664, IN47[47], Out1[47], w7763);
  FullAdder U2301 (w7763, w7666, IN48[47], w7764, w7765);
  FullAdder U2302 (w7765, w7668, IN49[47], w7766, w7767);
  FullAdder U2303 (w7767, w7670, IN50[47], w7768, w7769);
  FullAdder U2304 (w7769, w7672, IN51[45], w7770, w7771);
  FullAdder U2305 (w7771, w7674, IN52[44], w7772, w7773);
  FullAdder U2306 (w7773, w7676, IN53[43], w7774, w7775);
  FullAdder U2307 (w7775, w7678, IN54[42], w7776, w7777);
  FullAdder U2308 (w7777, w7680, IN55[41], w7778, w7779);
  FullAdder U2309 (w7779, w7682, IN56[40], w7780, w7781);
  FullAdder U2310 (w7781, w7684, IN57[39], w7782, w7783);
  FullAdder U2311 (w7783, w7686, IN58[38], w7784, w7785);
  FullAdder U2312 (w7785, w7688, IN59[37], w7786, w7787);
  FullAdder U2313 (w7787, w7690, IN60[36], w7788, w7789);
  FullAdder U2314 (w7789, w7692, IN61[35], w7790, w7791);
  FullAdder U2315 (w7791, w7694, IN62[34], w7792, w7793);
  FullAdder U2316 (w7793, w7696, IN63[33], w7794, w7795);
  FullAdder U2317 (w7795, w7698, IN64[32], w7796, w7797);
  FullAdder U2318 (w7797, w7700, IN65[31], w7798, w7799);
  FullAdder U2319 (w7799, w7702, IN66[30], w7800, w7801);
  FullAdder U2320 (w7801, w7704, IN67[29], w7802, w7803);
  FullAdder U2321 (w7803, w7706, IN68[28], w7804, w7805);
  FullAdder U2322 (w7805, w7708, IN69[27], w7806, w7807);
  FullAdder U2323 (w7807, w7710, IN70[26], w7808, w7809);
  FullAdder U2324 (w7809, w7712, IN71[25], w7810, w7811);
  FullAdder U2325 (w7811, w7714, IN72[24], w7812, w7813);
  FullAdder U2326 (w7813, w7716, IN73[23], w7814, w7815);
  FullAdder U2327 (w7815, w7718, IN74[22], w7816, w7817);
  FullAdder U2328 (w7817, w7720, IN75[21], w7818, w7819);
  FullAdder U2329 (w7819, w7722, IN76[20], w7820, w7821);
  FullAdder U2330 (w7821, w7724, IN77[19], w7822, w7823);
  FullAdder U2331 (w7823, w7726, IN78[18], w7824, w7825);
  FullAdder U2332 (w7825, w7728, IN79[17], w7826, w7827);
  FullAdder U2333 (w7827, w7730, IN80[16], w7828, w7829);
  FullAdder U2334 (w7829, w7732, IN81[15], w7830, w7831);
  FullAdder U2335 (w7831, w7734, IN82[14], w7832, w7833);
  FullAdder U2336 (w7833, w7736, IN83[13], w7834, w7835);
  FullAdder U2337 (w7835, w7738, IN84[12], w7836, w7837);
  FullAdder U2338 (w7837, w7740, IN85[11], w7838, w7839);
  FullAdder U2339 (w7839, w7742, IN86[10], w7840, w7841);
  FullAdder U2340 (w7841, w7744, IN87[9], w7842, w7843);
  FullAdder U2341 (w7843, w7746, IN88[8], w7844, w7845);
  FullAdder U2342 (w7845, w7748, IN89[7], w7846, w7847);
  FullAdder U2343 (w7847, w7750, IN90[6], w7848, w7849);
  FullAdder U2344 (w7849, w7752, IN91[5], w7850, w7851);
  FullAdder U2345 (w7851, w7754, IN92[4], w7852, w7853);
  FullAdder U2346 (w7853, w7756, IN93[3], w7854, w7855);
  FullAdder U2347 (w7855, w7758, IN94[2], w7856, w7857);
  FullAdder U2348 (w7857, w7760, IN95[1], w7858, w7859);
  FullAdder U2349 (w7859, w7761, IN96[0], w7860, w7861);
  HalfAdder U2350 (w7764, IN48[48], Out1[48], w7863);
  FullAdder U2351 (w7863, w7766, IN49[48], w7864, w7865);
  FullAdder U2352 (w7865, w7768, IN50[48], w7866, w7867);
  FullAdder U2353 (w7867, w7770, IN51[46], w7868, w7869);
  FullAdder U2354 (w7869, w7772, IN52[45], w7870, w7871);
  FullAdder U2355 (w7871, w7774, IN53[44], w7872, w7873);
  FullAdder U2356 (w7873, w7776, IN54[43], w7874, w7875);
  FullAdder U2357 (w7875, w7778, IN55[42], w7876, w7877);
  FullAdder U2358 (w7877, w7780, IN56[41], w7878, w7879);
  FullAdder U2359 (w7879, w7782, IN57[40], w7880, w7881);
  FullAdder U2360 (w7881, w7784, IN58[39], w7882, w7883);
  FullAdder U2361 (w7883, w7786, IN59[38], w7884, w7885);
  FullAdder U2362 (w7885, w7788, IN60[37], w7886, w7887);
  FullAdder U2363 (w7887, w7790, IN61[36], w7888, w7889);
  FullAdder U2364 (w7889, w7792, IN62[35], w7890, w7891);
  FullAdder U2365 (w7891, w7794, IN63[34], w7892, w7893);
  FullAdder U2366 (w7893, w7796, IN64[33], w7894, w7895);
  FullAdder U2367 (w7895, w7798, IN65[32], w7896, w7897);
  FullAdder U2368 (w7897, w7800, IN66[31], w7898, w7899);
  FullAdder U2369 (w7899, w7802, IN67[30], w7900, w7901);
  FullAdder U2370 (w7901, w7804, IN68[29], w7902, w7903);
  FullAdder U2371 (w7903, w7806, IN69[28], w7904, w7905);
  FullAdder U2372 (w7905, w7808, IN70[27], w7906, w7907);
  FullAdder U2373 (w7907, w7810, IN71[26], w7908, w7909);
  FullAdder U2374 (w7909, w7812, IN72[25], w7910, w7911);
  FullAdder U2375 (w7911, w7814, IN73[24], w7912, w7913);
  FullAdder U2376 (w7913, w7816, IN74[23], w7914, w7915);
  FullAdder U2377 (w7915, w7818, IN75[22], w7916, w7917);
  FullAdder U2378 (w7917, w7820, IN76[21], w7918, w7919);
  FullAdder U2379 (w7919, w7822, IN77[20], w7920, w7921);
  FullAdder U2380 (w7921, w7824, IN78[19], w7922, w7923);
  FullAdder U2381 (w7923, w7826, IN79[18], w7924, w7925);
  FullAdder U2382 (w7925, w7828, IN80[17], w7926, w7927);
  FullAdder U2383 (w7927, w7830, IN81[16], w7928, w7929);
  FullAdder U2384 (w7929, w7832, IN82[15], w7930, w7931);
  FullAdder U2385 (w7931, w7834, IN83[14], w7932, w7933);
  FullAdder U2386 (w7933, w7836, IN84[13], w7934, w7935);
  FullAdder U2387 (w7935, w7838, IN85[12], w7936, w7937);
  FullAdder U2388 (w7937, w7840, IN86[11], w7938, w7939);
  FullAdder U2389 (w7939, w7842, IN87[10], w7940, w7941);
  FullAdder U2390 (w7941, w7844, IN88[9], w7942, w7943);
  FullAdder U2391 (w7943, w7846, IN89[8], w7944, w7945);
  FullAdder U2392 (w7945, w7848, IN90[7], w7946, w7947);
  FullAdder U2393 (w7947, w7850, IN91[6], w7948, w7949);
  FullAdder U2394 (w7949, w7852, IN92[5], w7950, w7951);
  FullAdder U2395 (w7951, w7854, IN93[4], w7952, w7953);
  FullAdder U2396 (w7953, w7856, IN94[3], w7954, w7955);
  FullAdder U2397 (w7955, w7858, IN95[2], w7956, w7957);
  FullAdder U2398 (w7957, w7860, IN96[1], w7958, w7959);
  FullAdder U2399 (w7959, w7861, IN97[0], w7960, w7961);
  HalfAdder U2400 (w7864, IN49[49], Out1[49], w7963);
  FullAdder U2401 (w7963, w7866, IN50[49], w7964, w7965);
  FullAdder U2402 (w7965, w7868, IN51[47], w7966, w7967);
  FullAdder U2403 (w7967, w7870, IN52[46], w7968, w7969);
  FullAdder U2404 (w7969, w7872, IN53[45], w7970, w7971);
  FullAdder U2405 (w7971, w7874, IN54[44], w7972, w7973);
  FullAdder U2406 (w7973, w7876, IN55[43], w7974, w7975);
  FullAdder U2407 (w7975, w7878, IN56[42], w7976, w7977);
  FullAdder U2408 (w7977, w7880, IN57[41], w7978, w7979);
  FullAdder U2409 (w7979, w7882, IN58[40], w7980, w7981);
  FullAdder U2410 (w7981, w7884, IN59[39], w7982, w7983);
  FullAdder U2411 (w7983, w7886, IN60[38], w7984, w7985);
  FullAdder U2412 (w7985, w7888, IN61[37], w7986, w7987);
  FullAdder U2413 (w7987, w7890, IN62[36], w7988, w7989);
  FullAdder U2414 (w7989, w7892, IN63[35], w7990, w7991);
  FullAdder U2415 (w7991, w7894, IN64[34], w7992, w7993);
  FullAdder U2416 (w7993, w7896, IN65[33], w7994, w7995);
  FullAdder U2417 (w7995, w7898, IN66[32], w7996, w7997);
  FullAdder U2418 (w7997, w7900, IN67[31], w7998, w7999);
  FullAdder U2419 (w7999, w7902, IN68[30], w8000, w8001);
  FullAdder U2420 (w8001, w7904, IN69[29], w8002, w8003);
  FullAdder U2421 (w8003, w7906, IN70[28], w8004, w8005);
  FullAdder U2422 (w8005, w7908, IN71[27], w8006, w8007);
  FullAdder U2423 (w8007, w7910, IN72[26], w8008, w8009);
  FullAdder U2424 (w8009, w7912, IN73[25], w8010, w8011);
  FullAdder U2425 (w8011, w7914, IN74[24], w8012, w8013);
  FullAdder U2426 (w8013, w7916, IN75[23], w8014, w8015);
  FullAdder U2427 (w8015, w7918, IN76[22], w8016, w8017);
  FullAdder U2428 (w8017, w7920, IN77[21], w8018, w8019);
  FullAdder U2429 (w8019, w7922, IN78[20], w8020, w8021);
  FullAdder U2430 (w8021, w7924, IN79[19], w8022, w8023);
  FullAdder U2431 (w8023, w7926, IN80[18], w8024, w8025);
  FullAdder U2432 (w8025, w7928, IN81[17], w8026, w8027);
  FullAdder U2433 (w8027, w7930, IN82[16], w8028, w8029);
  FullAdder U2434 (w8029, w7932, IN83[15], w8030, w8031);
  FullAdder U2435 (w8031, w7934, IN84[14], w8032, w8033);
  FullAdder U2436 (w8033, w7936, IN85[13], w8034, w8035);
  FullAdder U2437 (w8035, w7938, IN86[12], w8036, w8037);
  FullAdder U2438 (w8037, w7940, IN87[11], w8038, w8039);
  FullAdder U2439 (w8039, w7942, IN88[10], w8040, w8041);
  FullAdder U2440 (w8041, w7944, IN89[9], w8042, w8043);
  FullAdder U2441 (w8043, w7946, IN90[8], w8044, w8045);
  FullAdder U2442 (w8045, w7948, IN91[7], w8046, w8047);
  FullAdder U2443 (w8047, w7950, IN92[6], w8048, w8049);
  FullAdder U2444 (w8049, w7952, IN93[5], w8050, w8051);
  FullAdder U2445 (w8051, w7954, IN94[4], w8052, w8053);
  FullAdder U2446 (w8053, w7956, IN95[3], w8054, w8055);
  FullAdder U2447 (w8055, w7958, IN96[2], w8056, w8057);
  FullAdder U2448 (w8057, w7960, IN97[1], w8058, w8059);
  FullAdder U2449 (w8059, w7961, IN98[0], w8060, w8061);
  HalfAdder U2450 (w7964, IN50[50], Out1[50], w8063);
  FullAdder U2451 (w8063, w7966, IN51[48], w8064, w8065);
  FullAdder U2452 (w8065, w7968, IN52[47], w8066, w8067);
  FullAdder U2453 (w8067, w7970, IN53[46], w8068, w8069);
  FullAdder U2454 (w8069, w7972, IN54[45], w8070, w8071);
  FullAdder U2455 (w8071, w7974, IN55[44], w8072, w8073);
  FullAdder U2456 (w8073, w7976, IN56[43], w8074, w8075);
  FullAdder U2457 (w8075, w7978, IN57[42], w8076, w8077);
  FullAdder U2458 (w8077, w7980, IN58[41], w8078, w8079);
  FullAdder U2459 (w8079, w7982, IN59[40], w8080, w8081);
  FullAdder U2460 (w8081, w7984, IN60[39], w8082, w8083);
  FullAdder U2461 (w8083, w7986, IN61[38], w8084, w8085);
  FullAdder U2462 (w8085, w7988, IN62[37], w8086, w8087);
  FullAdder U2463 (w8087, w7990, IN63[36], w8088, w8089);
  FullAdder U2464 (w8089, w7992, IN64[35], w8090, w8091);
  FullAdder U2465 (w8091, w7994, IN65[34], w8092, w8093);
  FullAdder U2466 (w8093, w7996, IN66[33], w8094, w8095);
  FullAdder U2467 (w8095, w7998, IN67[32], w8096, w8097);
  FullAdder U2468 (w8097, w8000, IN68[31], w8098, w8099);
  FullAdder U2469 (w8099, w8002, IN69[30], w8100, w8101);
  FullAdder U2470 (w8101, w8004, IN70[29], w8102, w8103);
  FullAdder U2471 (w8103, w8006, IN71[28], w8104, w8105);
  FullAdder U2472 (w8105, w8008, IN72[27], w8106, w8107);
  FullAdder U2473 (w8107, w8010, IN73[26], w8108, w8109);
  FullAdder U2474 (w8109, w8012, IN74[25], w8110, w8111);
  FullAdder U2475 (w8111, w8014, IN75[24], w8112, w8113);
  FullAdder U2476 (w8113, w8016, IN76[23], w8114, w8115);
  FullAdder U2477 (w8115, w8018, IN77[22], w8116, w8117);
  FullAdder U2478 (w8117, w8020, IN78[21], w8118, w8119);
  FullAdder U2479 (w8119, w8022, IN79[20], w8120, w8121);
  FullAdder U2480 (w8121, w8024, IN80[19], w8122, w8123);
  FullAdder U2481 (w8123, w8026, IN81[18], w8124, w8125);
  FullAdder U2482 (w8125, w8028, IN82[17], w8126, w8127);
  FullAdder U2483 (w8127, w8030, IN83[16], w8128, w8129);
  FullAdder U2484 (w8129, w8032, IN84[15], w8130, w8131);
  FullAdder U2485 (w8131, w8034, IN85[14], w8132, w8133);
  FullAdder U2486 (w8133, w8036, IN86[13], w8134, w8135);
  FullAdder U2487 (w8135, w8038, IN87[12], w8136, w8137);
  FullAdder U2488 (w8137, w8040, IN88[11], w8138, w8139);
  FullAdder U2489 (w8139, w8042, IN89[10], w8140, w8141);
  FullAdder U2490 (w8141, w8044, IN90[9], w8142, w8143);
  FullAdder U2491 (w8143, w8046, IN91[8], w8144, w8145);
  FullAdder U2492 (w8145, w8048, IN92[7], w8146, w8147);
  FullAdder U2493 (w8147, w8050, IN93[6], w8148, w8149);
  FullAdder U2494 (w8149, w8052, IN94[5], w8150, w8151);
  FullAdder U2495 (w8151, w8054, IN95[4], w8152, w8153);
  FullAdder U2496 (w8153, w8056, IN96[3], w8154, w8155);
  FullAdder U2497 (w8155, w8058, IN97[2], w8156, w8157);
  FullAdder U2498 (w8157, w8060, IN98[1], w8158, w8159);
  FullAdder U2499 (w8159, w8061, IN99[0], w8160, w8161);
  HalfAdder U2500 (w8064, IN51[49], Out1[51], w8163);
  FullAdder U2501 (w8163, w8066, IN52[48], w8164, w8165);
  FullAdder U2502 (w8165, w8068, IN53[47], w8166, w8167);
  FullAdder U2503 (w8167, w8070, IN54[46], w8168, w8169);
  FullAdder U2504 (w8169, w8072, IN55[45], w8170, w8171);
  FullAdder U2505 (w8171, w8074, IN56[44], w8172, w8173);
  FullAdder U2506 (w8173, w8076, IN57[43], w8174, w8175);
  FullAdder U2507 (w8175, w8078, IN58[42], w8176, w8177);
  FullAdder U2508 (w8177, w8080, IN59[41], w8178, w8179);
  FullAdder U2509 (w8179, w8082, IN60[40], w8180, w8181);
  FullAdder U2510 (w8181, w8084, IN61[39], w8182, w8183);
  FullAdder U2511 (w8183, w8086, IN62[38], w8184, w8185);
  FullAdder U2512 (w8185, w8088, IN63[37], w8186, w8187);
  FullAdder U2513 (w8187, w8090, IN64[36], w8188, w8189);
  FullAdder U2514 (w8189, w8092, IN65[35], w8190, w8191);
  FullAdder U2515 (w8191, w8094, IN66[34], w8192, w8193);
  FullAdder U2516 (w8193, w8096, IN67[33], w8194, w8195);
  FullAdder U2517 (w8195, w8098, IN68[32], w8196, w8197);
  FullAdder U2518 (w8197, w8100, IN69[31], w8198, w8199);
  FullAdder U2519 (w8199, w8102, IN70[30], w8200, w8201);
  FullAdder U2520 (w8201, w8104, IN71[29], w8202, w8203);
  FullAdder U2521 (w8203, w8106, IN72[28], w8204, w8205);
  FullAdder U2522 (w8205, w8108, IN73[27], w8206, w8207);
  FullAdder U2523 (w8207, w8110, IN74[26], w8208, w8209);
  FullAdder U2524 (w8209, w8112, IN75[25], w8210, w8211);
  FullAdder U2525 (w8211, w8114, IN76[24], w8212, w8213);
  FullAdder U2526 (w8213, w8116, IN77[23], w8214, w8215);
  FullAdder U2527 (w8215, w8118, IN78[22], w8216, w8217);
  FullAdder U2528 (w8217, w8120, IN79[21], w8218, w8219);
  FullAdder U2529 (w8219, w8122, IN80[20], w8220, w8221);
  FullAdder U2530 (w8221, w8124, IN81[19], w8222, w8223);
  FullAdder U2531 (w8223, w8126, IN82[18], w8224, w8225);
  FullAdder U2532 (w8225, w8128, IN83[17], w8226, w8227);
  FullAdder U2533 (w8227, w8130, IN84[16], w8228, w8229);
  FullAdder U2534 (w8229, w8132, IN85[15], w8230, w8231);
  FullAdder U2535 (w8231, w8134, IN86[14], w8232, w8233);
  FullAdder U2536 (w8233, w8136, IN87[13], w8234, w8235);
  FullAdder U2537 (w8235, w8138, IN88[12], w8236, w8237);
  FullAdder U2538 (w8237, w8140, IN89[11], w8238, w8239);
  FullAdder U2539 (w8239, w8142, IN90[10], w8240, w8241);
  FullAdder U2540 (w8241, w8144, IN91[9], w8242, w8243);
  FullAdder U2541 (w8243, w8146, IN92[8], w8244, w8245);
  FullAdder U2542 (w8245, w8148, IN93[7], w8246, w8247);
  FullAdder U2543 (w8247, w8150, IN94[6], w8248, w8249);
  FullAdder U2544 (w8249, w8152, IN95[5], w8250, w8251);
  FullAdder U2545 (w8251, w8154, IN96[4], w8252, w8253);
  FullAdder U2546 (w8253, w8156, IN97[3], w8254, w8255);
  FullAdder U2547 (w8255, w8158, IN98[2], w8256, w8257);
  FullAdder U2548 (w8257, w8160, IN99[1], w8258, w8259);
  FullAdder U2549 (w8259, w8161, IN100[0], w8260, w8261);
  HalfAdder U2550 (w8164, IN52[49], Out1[52], w8263);
  FullAdder U2551 (w8263, w8166, IN53[48], w8264, w8265);
  FullAdder U2552 (w8265, w8168, IN54[47], w8266, w8267);
  FullAdder U2553 (w8267, w8170, IN55[46], w8268, w8269);
  FullAdder U2554 (w8269, w8172, IN56[45], w8270, w8271);
  FullAdder U2555 (w8271, w8174, IN57[44], w8272, w8273);
  FullAdder U2556 (w8273, w8176, IN58[43], w8274, w8275);
  FullAdder U2557 (w8275, w8178, IN59[42], w8276, w8277);
  FullAdder U2558 (w8277, w8180, IN60[41], w8278, w8279);
  FullAdder U2559 (w8279, w8182, IN61[40], w8280, w8281);
  FullAdder U2560 (w8281, w8184, IN62[39], w8282, w8283);
  FullAdder U2561 (w8283, w8186, IN63[38], w8284, w8285);
  FullAdder U2562 (w8285, w8188, IN64[37], w8286, w8287);
  FullAdder U2563 (w8287, w8190, IN65[36], w8288, w8289);
  FullAdder U2564 (w8289, w8192, IN66[35], w8290, w8291);
  FullAdder U2565 (w8291, w8194, IN67[34], w8292, w8293);
  FullAdder U2566 (w8293, w8196, IN68[33], w8294, w8295);
  FullAdder U2567 (w8295, w8198, IN69[32], w8296, w8297);
  FullAdder U2568 (w8297, w8200, IN70[31], w8298, w8299);
  FullAdder U2569 (w8299, w8202, IN71[30], w8300, w8301);
  FullAdder U2570 (w8301, w8204, IN72[29], w8302, w8303);
  FullAdder U2571 (w8303, w8206, IN73[28], w8304, w8305);
  FullAdder U2572 (w8305, w8208, IN74[27], w8306, w8307);
  FullAdder U2573 (w8307, w8210, IN75[26], w8308, w8309);
  FullAdder U2574 (w8309, w8212, IN76[25], w8310, w8311);
  FullAdder U2575 (w8311, w8214, IN77[24], w8312, w8313);
  FullAdder U2576 (w8313, w8216, IN78[23], w8314, w8315);
  FullAdder U2577 (w8315, w8218, IN79[22], w8316, w8317);
  FullAdder U2578 (w8317, w8220, IN80[21], w8318, w8319);
  FullAdder U2579 (w8319, w8222, IN81[20], w8320, w8321);
  FullAdder U2580 (w8321, w8224, IN82[19], w8322, w8323);
  FullAdder U2581 (w8323, w8226, IN83[18], w8324, w8325);
  FullAdder U2582 (w8325, w8228, IN84[17], w8326, w8327);
  FullAdder U2583 (w8327, w8230, IN85[16], w8328, w8329);
  FullAdder U2584 (w8329, w8232, IN86[15], w8330, w8331);
  FullAdder U2585 (w8331, w8234, IN87[14], w8332, w8333);
  FullAdder U2586 (w8333, w8236, IN88[13], w8334, w8335);
  FullAdder U2587 (w8335, w8238, IN89[12], w8336, w8337);
  FullAdder U2588 (w8337, w8240, IN90[11], w8338, w8339);
  FullAdder U2589 (w8339, w8242, IN91[10], w8340, w8341);
  FullAdder U2590 (w8341, w8244, IN92[9], w8342, w8343);
  FullAdder U2591 (w8343, w8246, IN93[8], w8344, w8345);
  FullAdder U2592 (w8345, w8248, IN94[7], w8346, w8347);
  FullAdder U2593 (w8347, w8250, IN95[6], w8348, w8349);
  FullAdder U2594 (w8349, w8252, IN96[5], w8350, w8351);
  FullAdder U2595 (w8351, w8254, IN97[4], w8352, w8353);
  FullAdder U2596 (w8353, w8256, IN98[3], w8354, w8355);
  FullAdder U2597 (w8355, w8258, IN99[2], w8356, w8357);
  FullAdder U2598 (w8357, w8260, IN100[1], w8358, w8359);
  FullAdder U2599 (w8359, w8261, IN101[0], w8360, w8361);
  HalfAdder U2600 (w8264, IN53[49], Out1[53], w8363);
  FullAdder U2601 (w8363, w8266, IN54[48], w8364, w8365);
  FullAdder U2602 (w8365, w8268, IN55[47], w8366, w8367);
  FullAdder U2603 (w8367, w8270, IN56[46], w8368, w8369);
  FullAdder U2604 (w8369, w8272, IN57[45], w8370, w8371);
  FullAdder U2605 (w8371, w8274, IN58[44], w8372, w8373);
  FullAdder U2606 (w8373, w8276, IN59[43], w8374, w8375);
  FullAdder U2607 (w8375, w8278, IN60[42], w8376, w8377);
  FullAdder U2608 (w8377, w8280, IN61[41], w8378, w8379);
  FullAdder U2609 (w8379, w8282, IN62[40], w8380, w8381);
  FullAdder U2610 (w8381, w8284, IN63[39], w8382, w8383);
  FullAdder U2611 (w8383, w8286, IN64[38], w8384, w8385);
  FullAdder U2612 (w8385, w8288, IN65[37], w8386, w8387);
  FullAdder U2613 (w8387, w8290, IN66[36], w8388, w8389);
  FullAdder U2614 (w8389, w8292, IN67[35], w8390, w8391);
  FullAdder U2615 (w8391, w8294, IN68[34], w8392, w8393);
  FullAdder U2616 (w8393, w8296, IN69[33], w8394, w8395);
  FullAdder U2617 (w8395, w8298, IN70[32], w8396, w8397);
  FullAdder U2618 (w8397, w8300, IN71[31], w8398, w8399);
  FullAdder U2619 (w8399, w8302, IN72[30], w8400, w8401);
  FullAdder U2620 (w8401, w8304, IN73[29], w8402, w8403);
  FullAdder U2621 (w8403, w8306, IN74[28], w8404, w8405);
  FullAdder U2622 (w8405, w8308, IN75[27], w8406, w8407);
  FullAdder U2623 (w8407, w8310, IN76[26], w8408, w8409);
  FullAdder U2624 (w8409, w8312, IN77[25], w8410, w8411);
  FullAdder U2625 (w8411, w8314, IN78[24], w8412, w8413);
  FullAdder U2626 (w8413, w8316, IN79[23], w8414, w8415);
  FullAdder U2627 (w8415, w8318, IN80[22], w8416, w8417);
  FullAdder U2628 (w8417, w8320, IN81[21], w8418, w8419);
  FullAdder U2629 (w8419, w8322, IN82[20], w8420, w8421);
  FullAdder U2630 (w8421, w8324, IN83[19], w8422, w8423);
  FullAdder U2631 (w8423, w8326, IN84[18], w8424, w8425);
  FullAdder U2632 (w8425, w8328, IN85[17], w8426, w8427);
  FullAdder U2633 (w8427, w8330, IN86[16], w8428, w8429);
  FullAdder U2634 (w8429, w8332, IN87[15], w8430, w8431);
  FullAdder U2635 (w8431, w8334, IN88[14], w8432, w8433);
  FullAdder U2636 (w8433, w8336, IN89[13], w8434, w8435);
  FullAdder U2637 (w8435, w8338, IN90[12], w8436, w8437);
  FullAdder U2638 (w8437, w8340, IN91[11], w8438, w8439);
  FullAdder U2639 (w8439, w8342, IN92[10], w8440, w8441);
  FullAdder U2640 (w8441, w8344, IN93[9], w8442, w8443);
  FullAdder U2641 (w8443, w8346, IN94[8], w8444, w8445);
  FullAdder U2642 (w8445, w8348, IN95[7], w8446, w8447);
  FullAdder U2643 (w8447, w8350, IN96[6], w8448, w8449);
  FullAdder U2644 (w8449, w8352, IN97[5], w8450, w8451);
  FullAdder U2645 (w8451, w8354, IN98[4], w8452, w8453);
  FullAdder U2646 (w8453, w8356, IN99[3], w8454, w8455);
  FullAdder U2647 (w8455, w8358, IN100[2], w8456, w8457);
  FullAdder U2648 (w8457, w8360, IN101[1], w8458, w8459);
  FullAdder U2649 (w8459, w8361, IN102[0], w8460, w8461);
  HalfAdder U2650 (w8364, IN54[49], Out1[54], w8463);
  FullAdder U2651 (w8463, w8366, IN55[48], w8464, w8465);
  FullAdder U2652 (w8465, w8368, IN56[47], w8466, w8467);
  FullAdder U2653 (w8467, w8370, IN57[46], w8468, w8469);
  FullAdder U2654 (w8469, w8372, IN58[45], w8470, w8471);
  FullAdder U2655 (w8471, w8374, IN59[44], w8472, w8473);
  FullAdder U2656 (w8473, w8376, IN60[43], w8474, w8475);
  FullAdder U2657 (w8475, w8378, IN61[42], w8476, w8477);
  FullAdder U2658 (w8477, w8380, IN62[41], w8478, w8479);
  FullAdder U2659 (w8479, w8382, IN63[40], w8480, w8481);
  FullAdder U2660 (w8481, w8384, IN64[39], w8482, w8483);
  FullAdder U2661 (w8483, w8386, IN65[38], w8484, w8485);
  FullAdder U2662 (w8485, w8388, IN66[37], w8486, w8487);
  FullAdder U2663 (w8487, w8390, IN67[36], w8488, w8489);
  FullAdder U2664 (w8489, w8392, IN68[35], w8490, w8491);
  FullAdder U2665 (w8491, w8394, IN69[34], w8492, w8493);
  FullAdder U2666 (w8493, w8396, IN70[33], w8494, w8495);
  FullAdder U2667 (w8495, w8398, IN71[32], w8496, w8497);
  FullAdder U2668 (w8497, w8400, IN72[31], w8498, w8499);
  FullAdder U2669 (w8499, w8402, IN73[30], w8500, w8501);
  FullAdder U2670 (w8501, w8404, IN74[29], w8502, w8503);
  FullAdder U2671 (w8503, w8406, IN75[28], w8504, w8505);
  FullAdder U2672 (w8505, w8408, IN76[27], w8506, w8507);
  FullAdder U2673 (w8507, w8410, IN77[26], w8508, w8509);
  FullAdder U2674 (w8509, w8412, IN78[25], w8510, w8511);
  FullAdder U2675 (w8511, w8414, IN79[24], w8512, w8513);
  FullAdder U2676 (w8513, w8416, IN80[23], w8514, w8515);
  FullAdder U2677 (w8515, w8418, IN81[22], w8516, w8517);
  FullAdder U2678 (w8517, w8420, IN82[21], w8518, w8519);
  FullAdder U2679 (w8519, w8422, IN83[20], w8520, w8521);
  FullAdder U2680 (w8521, w8424, IN84[19], w8522, w8523);
  FullAdder U2681 (w8523, w8426, IN85[18], w8524, w8525);
  FullAdder U2682 (w8525, w8428, IN86[17], w8526, w8527);
  FullAdder U2683 (w8527, w8430, IN87[16], w8528, w8529);
  FullAdder U2684 (w8529, w8432, IN88[15], w8530, w8531);
  FullAdder U2685 (w8531, w8434, IN89[14], w8532, w8533);
  FullAdder U2686 (w8533, w8436, IN90[13], w8534, w8535);
  FullAdder U2687 (w8535, w8438, IN91[12], w8536, w8537);
  FullAdder U2688 (w8537, w8440, IN92[11], w8538, w8539);
  FullAdder U2689 (w8539, w8442, IN93[10], w8540, w8541);
  FullAdder U2690 (w8541, w8444, IN94[9], w8542, w8543);
  FullAdder U2691 (w8543, w8446, IN95[8], w8544, w8545);
  FullAdder U2692 (w8545, w8448, IN96[7], w8546, w8547);
  FullAdder U2693 (w8547, w8450, IN97[6], w8548, w8549);
  FullAdder U2694 (w8549, w8452, IN98[5], w8550, w8551);
  FullAdder U2695 (w8551, w8454, IN99[4], w8552, w8553);
  FullAdder U2696 (w8553, w8456, IN100[3], w8554, w8555);
  FullAdder U2697 (w8555, w8458, IN101[2], w8556, w8557);
  FullAdder U2698 (w8557, w8460, IN102[1], w8558, w8559);
  FullAdder U2699 (w8559, w8461, IN103[0], w8560, w8561);
  HalfAdder U2700 (w8464, IN55[49], Out1[55], w8563);
  FullAdder U2701 (w8563, w8466, IN56[48], w8564, w8565);
  FullAdder U2702 (w8565, w8468, IN57[47], w8566, w8567);
  FullAdder U2703 (w8567, w8470, IN58[46], w8568, w8569);
  FullAdder U2704 (w8569, w8472, IN59[45], w8570, w8571);
  FullAdder U2705 (w8571, w8474, IN60[44], w8572, w8573);
  FullAdder U2706 (w8573, w8476, IN61[43], w8574, w8575);
  FullAdder U2707 (w8575, w8478, IN62[42], w8576, w8577);
  FullAdder U2708 (w8577, w8480, IN63[41], w8578, w8579);
  FullAdder U2709 (w8579, w8482, IN64[40], w8580, w8581);
  FullAdder U2710 (w8581, w8484, IN65[39], w8582, w8583);
  FullAdder U2711 (w8583, w8486, IN66[38], w8584, w8585);
  FullAdder U2712 (w8585, w8488, IN67[37], w8586, w8587);
  FullAdder U2713 (w8587, w8490, IN68[36], w8588, w8589);
  FullAdder U2714 (w8589, w8492, IN69[35], w8590, w8591);
  FullAdder U2715 (w8591, w8494, IN70[34], w8592, w8593);
  FullAdder U2716 (w8593, w8496, IN71[33], w8594, w8595);
  FullAdder U2717 (w8595, w8498, IN72[32], w8596, w8597);
  FullAdder U2718 (w8597, w8500, IN73[31], w8598, w8599);
  FullAdder U2719 (w8599, w8502, IN74[30], w8600, w8601);
  FullAdder U2720 (w8601, w8504, IN75[29], w8602, w8603);
  FullAdder U2721 (w8603, w8506, IN76[28], w8604, w8605);
  FullAdder U2722 (w8605, w8508, IN77[27], w8606, w8607);
  FullAdder U2723 (w8607, w8510, IN78[26], w8608, w8609);
  FullAdder U2724 (w8609, w8512, IN79[25], w8610, w8611);
  FullAdder U2725 (w8611, w8514, IN80[24], w8612, w8613);
  FullAdder U2726 (w8613, w8516, IN81[23], w8614, w8615);
  FullAdder U2727 (w8615, w8518, IN82[22], w8616, w8617);
  FullAdder U2728 (w8617, w8520, IN83[21], w8618, w8619);
  FullAdder U2729 (w8619, w8522, IN84[20], w8620, w8621);
  FullAdder U2730 (w8621, w8524, IN85[19], w8622, w8623);
  FullAdder U2731 (w8623, w8526, IN86[18], w8624, w8625);
  FullAdder U2732 (w8625, w8528, IN87[17], w8626, w8627);
  FullAdder U2733 (w8627, w8530, IN88[16], w8628, w8629);
  FullAdder U2734 (w8629, w8532, IN89[15], w8630, w8631);
  FullAdder U2735 (w8631, w8534, IN90[14], w8632, w8633);
  FullAdder U2736 (w8633, w8536, IN91[13], w8634, w8635);
  FullAdder U2737 (w8635, w8538, IN92[12], w8636, w8637);
  FullAdder U2738 (w8637, w8540, IN93[11], w8638, w8639);
  FullAdder U2739 (w8639, w8542, IN94[10], w8640, w8641);
  FullAdder U2740 (w8641, w8544, IN95[9], w8642, w8643);
  FullAdder U2741 (w8643, w8546, IN96[8], w8644, w8645);
  FullAdder U2742 (w8645, w8548, IN97[7], w8646, w8647);
  FullAdder U2743 (w8647, w8550, IN98[6], w8648, w8649);
  FullAdder U2744 (w8649, w8552, IN99[5], w8650, w8651);
  FullAdder U2745 (w8651, w8554, IN100[4], w8652, w8653);
  FullAdder U2746 (w8653, w8556, IN101[3], w8654, w8655);
  FullAdder U2747 (w8655, w8558, IN102[2], w8656, w8657);
  FullAdder U2748 (w8657, w8560, IN103[1], w8658, w8659);
  FullAdder U2749 (w8659, w8561, IN104[0], w8660, w8661);
  HalfAdder U2750 (w8564, IN56[49], Out1[56], w8663);
  FullAdder U2751 (w8663, w8566, IN57[48], w8664, w8665);
  FullAdder U2752 (w8665, w8568, IN58[47], w8666, w8667);
  FullAdder U2753 (w8667, w8570, IN59[46], w8668, w8669);
  FullAdder U2754 (w8669, w8572, IN60[45], w8670, w8671);
  FullAdder U2755 (w8671, w8574, IN61[44], w8672, w8673);
  FullAdder U2756 (w8673, w8576, IN62[43], w8674, w8675);
  FullAdder U2757 (w8675, w8578, IN63[42], w8676, w8677);
  FullAdder U2758 (w8677, w8580, IN64[41], w8678, w8679);
  FullAdder U2759 (w8679, w8582, IN65[40], w8680, w8681);
  FullAdder U2760 (w8681, w8584, IN66[39], w8682, w8683);
  FullAdder U2761 (w8683, w8586, IN67[38], w8684, w8685);
  FullAdder U2762 (w8685, w8588, IN68[37], w8686, w8687);
  FullAdder U2763 (w8687, w8590, IN69[36], w8688, w8689);
  FullAdder U2764 (w8689, w8592, IN70[35], w8690, w8691);
  FullAdder U2765 (w8691, w8594, IN71[34], w8692, w8693);
  FullAdder U2766 (w8693, w8596, IN72[33], w8694, w8695);
  FullAdder U2767 (w8695, w8598, IN73[32], w8696, w8697);
  FullAdder U2768 (w8697, w8600, IN74[31], w8698, w8699);
  FullAdder U2769 (w8699, w8602, IN75[30], w8700, w8701);
  FullAdder U2770 (w8701, w8604, IN76[29], w8702, w8703);
  FullAdder U2771 (w8703, w8606, IN77[28], w8704, w8705);
  FullAdder U2772 (w8705, w8608, IN78[27], w8706, w8707);
  FullAdder U2773 (w8707, w8610, IN79[26], w8708, w8709);
  FullAdder U2774 (w8709, w8612, IN80[25], w8710, w8711);
  FullAdder U2775 (w8711, w8614, IN81[24], w8712, w8713);
  FullAdder U2776 (w8713, w8616, IN82[23], w8714, w8715);
  FullAdder U2777 (w8715, w8618, IN83[22], w8716, w8717);
  FullAdder U2778 (w8717, w8620, IN84[21], w8718, w8719);
  FullAdder U2779 (w8719, w8622, IN85[20], w8720, w8721);
  FullAdder U2780 (w8721, w8624, IN86[19], w8722, w8723);
  FullAdder U2781 (w8723, w8626, IN87[18], w8724, w8725);
  FullAdder U2782 (w8725, w8628, IN88[17], w8726, w8727);
  FullAdder U2783 (w8727, w8630, IN89[16], w8728, w8729);
  FullAdder U2784 (w8729, w8632, IN90[15], w8730, w8731);
  FullAdder U2785 (w8731, w8634, IN91[14], w8732, w8733);
  FullAdder U2786 (w8733, w8636, IN92[13], w8734, w8735);
  FullAdder U2787 (w8735, w8638, IN93[12], w8736, w8737);
  FullAdder U2788 (w8737, w8640, IN94[11], w8738, w8739);
  FullAdder U2789 (w8739, w8642, IN95[10], w8740, w8741);
  FullAdder U2790 (w8741, w8644, IN96[9], w8742, w8743);
  FullAdder U2791 (w8743, w8646, IN97[8], w8744, w8745);
  FullAdder U2792 (w8745, w8648, IN98[7], w8746, w8747);
  FullAdder U2793 (w8747, w8650, IN99[6], w8748, w8749);
  FullAdder U2794 (w8749, w8652, IN100[5], w8750, w8751);
  FullAdder U2795 (w8751, w8654, IN101[4], w8752, w8753);
  FullAdder U2796 (w8753, w8656, IN102[3], w8754, w8755);
  FullAdder U2797 (w8755, w8658, IN103[2], w8756, w8757);
  FullAdder U2798 (w8757, w8660, IN104[1], w8758, w8759);
  FullAdder U2799 (w8759, w8661, IN105[0], w8760, w8761);
  HalfAdder U2800 (w8664, IN57[49], Out1[57], w8763);
  FullAdder U2801 (w8763, w8666, IN58[48], w8764, w8765);
  FullAdder U2802 (w8765, w8668, IN59[47], w8766, w8767);
  FullAdder U2803 (w8767, w8670, IN60[46], w8768, w8769);
  FullAdder U2804 (w8769, w8672, IN61[45], w8770, w8771);
  FullAdder U2805 (w8771, w8674, IN62[44], w8772, w8773);
  FullAdder U2806 (w8773, w8676, IN63[43], w8774, w8775);
  FullAdder U2807 (w8775, w8678, IN64[42], w8776, w8777);
  FullAdder U2808 (w8777, w8680, IN65[41], w8778, w8779);
  FullAdder U2809 (w8779, w8682, IN66[40], w8780, w8781);
  FullAdder U2810 (w8781, w8684, IN67[39], w8782, w8783);
  FullAdder U2811 (w8783, w8686, IN68[38], w8784, w8785);
  FullAdder U2812 (w8785, w8688, IN69[37], w8786, w8787);
  FullAdder U2813 (w8787, w8690, IN70[36], w8788, w8789);
  FullAdder U2814 (w8789, w8692, IN71[35], w8790, w8791);
  FullAdder U2815 (w8791, w8694, IN72[34], w8792, w8793);
  FullAdder U2816 (w8793, w8696, IN73[33], w8794, w8795);
  FullAdder U2817 (w8795, w8698, IN74[32], w8796, w8797);
  FullAdder U2818 (w8797, w8700, IN75[31], w8798, w8799);
  FullAdder U2819 (w8799, w8702, IN76[30], w8800, w8801);
  FullAdder U2820 (w8801, w8704, IN77[29], w8802, w8803);
  FullAdder U2821 (w8803, w8706, IN78[28], w8804, w8805);
  FullAdder U2822 (w8805, w8708, IN79[27], w8806, w8807);
  FullAdder U2823 (w8807, w8710, IN80[26], w8808, w8809);
  FullAdder U2824 (w8809, w8712, IN81[25], w8810, w8811);
  FullAdder U2825 (w8811, w8714, IN82[24], w8812, w8813);
  FullAdder U2826 (w8813, w8716, IN83[23], w8814, w8815);
  FullAdder U2827 (w8815, w8718, IN84[22], w8816, w8817);
  FullAdder U2828 (w8817, w8720, IN85[21], w8818, w8819);
  FullAdder U2829 (w8819, w8722, IN86[20], w8820, w8821);
  FullAdder U2830 (w8821, w8724, IN87[19], w8822, w8823);
  FullAdder U2831 (w8823, w8726, IN88[18], w8824, w8825);
  FullAdder U2832 (w8825, w8728, IN89[17], w8826, w8827);
  FullAdder U2833 (w8827, w8730, IN90[16], w8828, w8829);
  FullAdder U2834 (w8829, w8732, IN91[15], w8830, w8831);
  FullAdder U2835 (w8831, w8734, IN92[14], w8832, w8833);
  FullAdder U2836 (w8833, w8736, IN93[13], w8834, w8835);
  FullAdder U2837 (w8835, w8738, IN94[12], w8836, w8837);
  FullAdder U2838 (w8837, w8740, IN95[11], w8838, w8839);
  FullAdder U2839 (w8839, w8742, IN96[10], w8840, w8841);
  FullAdder U2840 (w8841, w8744, IN97[9], w8842, w8843);
  FullAdder U2841 (w8843, w8746, IN98[8], w8844, w8845);
  FullAdder U2842 (w8845, w8748, IN99[7], w8846, w8847);
  FullAdder U2843 (w8847, w8750, IN100[6], w8848, w8849);
  FullAdder U2844 (w8849, w8752, IN101[5], w8850, w8851);
  FullAdder U2845 (w8851, w8754, IN102[4], w8852, w8853);
  FullAdder U2846 (w8853, w8756, IN103[3], w8854, w8855);
  FullAdder U2847 (w8855, w8758, IN104[2], w8856, w8857);
  FullAdder U2848 (w8857, w8760, IN105[1], w8858, w8859);
  FullAdder U2849 (w8859, w8761, IN106[0], w8860, w8861);
  HalfAdder U2850 (w8764, IN58[49], Out1[58], w8863);
  FullAdder U2851 (w8863, w8766, IN59[48], w8864, w8865);
  FullAdder U2852 (w8865, w8768, IN60[47], w8866, w8867);
  FullAdder U2853 (w8867, w8770, IN61[46], w8868, w8869);
  FullAdder U2854 (w8869, w8772, IN62[45], w8870, w8871);
  FullAdder U2855 (w8871, w8774, IN63[44], w8872, w8873);
  FullAdder U2856 (w8873, w8776, IN64[43], w8874, w8875);
  FullAdder U2857 (w8875, w8778, IN65[42], w8876, w8877);
  FullAdder U2858 (w8877, w8780, IN66[41], w8878, w8879);
  FullAdder U2859 (w8879, w8782, IN67[40], w8880, w8881);
  FullAdder U2860 (w8881, w8784, IN68[39], w8882, w8883);
  FullAdder U2861 (w8883, w8786, IN69[38], w8884, w8885);
  FullAdder U2862 (w8885, w8788, IN70[37], w8886, w8887);
  FullAdder U2863 (w8887, w8790, IN71[36], w8888, w8889);
  FullAdder U2864 (w8889, w8792, IN72[35], w8890, w8891);
  FullAdder U2865 (w8891, w8794, IN73[34], w8892, w8893);
  FullAdder U2866 (w8893, w8796, IN74[33], w8894, w8895);
  FullAdder U2867 (w8895, w8798, IN75[32], w8896, w8897);
  FullAdder U2868 (w8897, w8800, IN76[31], w8898, w8899);
  FullAdder U2869 (w8899, w8802, IN77[30], w8900, w8901);
  FullAdder U2870 (w8901, w8804, IN78[29], w8902, w8903);
  FullAdder U2871 (w8903, w8806, IN79[28], w8904, w8905);
  FullAdder U2872 (w8905, w8808, IN80[27], w8906, w8907);
  FullAdder U2873 (w8907, w8810, IN81[26], w8908, w8909);
  FullAdder U2874 (w8909, w8812, IN82[25], w8910, w8911);
  FullAdder U2875 (w8911, w8814, IN83[24], w8912, w8913);
  FullAdder U2876 (w8913, w8816, IN84[23], w8914, w8915);
  FullAdder U2877 (w8915, w8818, IN85[22], w8916, w8917);
  FullAdder U2878 (w8917, w8820, IN86[21], w8918, w8919);
  FullAdder U2879 (w8919, w8822, IN87[20], w8920, w8921);
  FullAdder U2880 (w8921, w8824, IN88[19], w8922, w8923);
  FullAdder U2881 (w8923, w8826, IN89[18], w8924, w8925);
  FullAdder U2882 (w8925, w8828, IN90[17], w8926, w8927);
  FullAdder U2883 (w8927, w8830, IN91[16], w8928, w8929);
  FullAdder U2884 (w8929, w8832, IN92[15], w8930, w8931);
  FullAdder U2885 (w8931, w8834, IN93[14], w8932, w8933);
  FullAdder U2886 (w8933, w8836, IN94[13], w8934, w8935);
  FullAdder U2887 (w8935, w8838, IN95[12], w8936, w8937);
  FullAdder U2888 (w8937, w8840, IN96[11], w8938, w8939);
  FullAdder U2889 (w8939, w8842, IN97[10], w8940, w8941);
  FullAdder U2890 (w8941, w8844, IN98[9], w8942, w8943);
  FullAdder U2891 (w8943, w8846, IN99[8], w8944, w8945);
  FullAdder U2892 (w8945, w8848, IN100[7], w8946, w8947);
  FullAdder U2893 (w8947, w8850, IN101[6], w8948, w8949);
  FullAdder U2894 (w8949, w8852, IN102[5], w8950, w8951);
  FullAdder U2895 (w8951, w8854, IN103[4], w8952, w8953);
  FullAdder U2896 (w8953, w8856, IN104[3], w8954, w8955);
  FullAdder U2897 (w8955, w8858, IN105[2], w8956, w8957);
  FullAdder U2898 (w8957, w8860, IN106[1], w8958, w8959);
  FullAdder U2899 (w8959, w8861, IN107[0], w8960, w8961);
  HalfAdder U2900 (w8864, IN59[49], Out1[59], w8963);
  FullAdder U2901 (w8963, w8866, IN60[48], w8964, w8965);
  FullAdder U2902 (w8965, w8868, IN61[47], w8966, w8967);
  FullAdder U2903 (w8967, w8870, IN62[46], w8968, w8969);
  FullAdder U2904 (w8969, w8872, IN63[45], w8970, w8971);
  FullAdder U2905 (w8971, w8874, IN64[44], w8972, w8973);
  FullAdder U2906 (w8973, w8876, IN65[43], w8974, w8975);
  FullAdder U2907 (w8975, w8878, IN66[42], w8976, w8977);
  FullAdder U2908 (w8977, w8880, IN67[41], w8978, w8979);
  FullAdder U2909 (w8979, w8882, IN68[40], w8980, w8981);
  FullAdder U2910 (w8981, w8884, IN69[39], w8982, w8983);
  FullAdder U2911 (w8983, w8886, IN70[38], w8984, w8985);
  FullAdder U2912 (w8985, w8888, IN71[37], w8986, w8987);
  FullAdder U2913 (w8987, w8890, IN72[36], w8988, w8989);
  FullAdder U2914 (w8989, w8892, IN73[35], w8990, w8991);
  FullAdder U2915 (w8991, w8894, IN74[34], w8992, w8993);
  FullAdder U2916 (w8993, w8896, IN75[33], w8994, w8995);
  FullAdder U2917 (w8995, w8898, IN76[32], w8996, w8997);
  FullAdder U2918 (w8997, w8900, IN77[31], w8998, w8999);
  FullAdder U2919 (w8999, w8902, IN78[30], w9000, w9001);
  FullAdder U2920 (w9001, w8904, IN79[29], w9002, w9003);
  FullAdder U2921 (w9003, w8906, IN80[28], w9004, w9005);
  FullAdder U2922 (w9005, w8908, IN81[27], w9006, w9007);
  FullAdder U2923 (w9007, w8910, IN82[26], w9008, w9009);
  FullAdder U2924 (w9009, w8912, IN83[25], w9010, w9011);
  FullAdder U2925 (w9011, w8914, IN84[24], w9012, w9013);
  FullAdder U2926 (w9013, w8916, IN85[23], w9014, w9015);
  FullAdder U2927 (w9015, w8918, IN86[22], w9016, w9017);
  FullAdder U2928 (w9017, w8920, IN87[21], w9018, w9019);
  FullAdder U2929 (w9019, w8922, IN88[20], w9020, w9021);
  FullAdder U2930 (w9021, w8924, IN89[19], w9022, w9023);
  FullAdder U2931 (w9023, w8926, IN90[18], w9024, w9025);
  FullAdder U2932 (w9025, w8928, IN91[17], w9026, w9027);
  FullAdder U2933 (w9027, w8930, IN92[16], w9028, w9029);
  FullAdder U2934 (w9029, w8932, IN93[15], w9030, w9031);
  FullAdder U2935 (w9031, w8934, IN94[14], w9032, w9033);
  FullAdder U2936 (w9033, w8936, IN95[13], w9034, w9035);
  FullAdder U2937 (w9035, w8938, IN96[12], w9036, w9037);
  FullAdder U2938 (w9037, w8940, IN97[11], w9038, w9039);
  FullAdder U2939 (w9039, w8942, IN98[10], w9040, w9041);
  FullAdder U2940 (w9041, w8944, IN99[9], w9042, w9043);
  FullAdder U2941 (w9043, w8946, IN100[8], w9044, w9045);
  FullAdder U2942 (w9045, w8948, IN101[7], w9046, w9047);
  FullAdder U2943 (w9047, w8950, IN102[6], w9048, w9049);
  FullAdder U2944 (w9049, w8952, IN103[5], w9050, w9051);
  FullAdder U2945 (w9051, w8954, IN104[4], w9052, w9053);
  FullAdder U2946 (w9053, w8956, IN105[3], w9054, w9055);
  FullAdder U2947 (w9055, w8958, IN106[2], w9056, w9057);
  FullAdder U2948 (w9057, w8960, IN107[1], w9058, w9059);
  FullAdder U2949 (w9059, w8961, IN108[0], w9060, w9061);
  HalfAdder U2950 (w8964, IN60[49], Out1[60], w9063);
  FullAdder U2951 (w9063, w8966, IN61[48], w9064, w9065);
  FullAdder U2952 (w9065, w8968, IN62[47], w9066, w9067);
  FullAdder U2953 (w9067, w8970, IN63[46], w9068, w9069);
  FullAdder U2954 (w9069, w8972, IN64[45], w9070, w9071);
  FullAdder U2955 (w9071, w8974, IN65[44], w9072, w9073);
  FullAdder U2956 (w9073, w8976, IN66[43], w9074, w9075);
  FullAdder U2957 (w9075, w8978, IN67[42], w9076, w9077);
  FullAdder U2958 (w9077, w8980, IN68[41], w9078, w9079);
  FullAdder U2959 (w9079, w8982, IN69[40], w9080, w9081);
  FullAdder U2960 (w9081, w8984, IN70[39], w9082, w9083);
  FullAdder U2961 (w9083, w8986, IN71[38], w9084, w9085);
  FullAdder U2962 (w9085, w8988, IN72[37], w9086, w9087);
  FullAdder U2963 (w9087, w8990, IN73[36], w9088, w9089);
  FullAdder U2964 (w9089, w8992, IN74[35], w9090, w9091);
  FullAdder U2965 (w9091, w8994, IN75[34], w9092, w9093);
  FullAdder U2966 (w9093, w8996, IN76[33], w9094, w9095);
  FullAdder U2967 (w9095, w8998, IN77[32], w9096, w9097);
  FullAdder U2968 (w9097, w9000, IN78[31], w9098, w9099);
  FullAdder U2969 (w9099, w9002, IN79[30], w9100, w9101);
  FullAdder U2970 (w9101, w9004, IN80[29], w9102, w9103);
  FullAdder U2971 (w9103, w9006, IN81[28], w9104, w9105);
  FullAdder U2972 (w9105, w9008, IN82[27], w9106, w9107);
  FullAdder U2973 (w9107, w9010, IN83[26], w9108, w9109);
  FullAdder U2974 (w9109, w9012, IN84[25], w9110, w9111);
  FullAdder U2975 (w9111, w9014, IN85[24], w9112, w9113);
  FullAdder U2976 (w9113, w9016, IN86[23], w9114, w9115);
  FullAdder U2977 (w9115, w9018, IN87[22], w9116, w9117);
  FullAdder U2978 (w9117, w9020, IN88[21], w9118, w9119);
  FullAdder U2979 (w9119, w9022, IN89[20], w9120, w9121);
  FullAdder U2980 (w9121, w9024, IN90[19], w9122, w9123);
  FullAdder U2981 (w9123, w9026, IN91[18], w9124, w9125);
  FullAdder U2982 (w9125, w9028, IN92[17], w9126, w9127);
  FullAdder U2983 (w9127, w9030, IN93[16], w9128, w9129);
  FullAdder U2984 (w9129, w9032, IN94[15], w9130, w9131);
  FullAdder U2985 (w9131, w9034, IN95[14], w9132, w9133);
  FullAdder U2986 (w9133, w9036, IN96[13], w9134, w9135);
  FullAdder U2987 (w9135, w9038, IN97[12], w9136, w9137);
  FullAdder U2988 (w9137, w9040, IN98[11], w9138, w9139);
  FullAdder U2989 (w9139, w9042, IN99[10], w9140, w9141);
  FullAdder U2990 (w9141, w9044, IN100[9], w9142, w9143);
  FullAdder U2991 (w9143, w9046, IN101[8], w9144, w9145);
  FullAdder U2992 (w9145, w9048, IN102[7], w9146, w9147);
  FullAdder U2993 (w9147, w9050, IN103[6], w9148, w9149);
  FullAdder U2994 (w9149, w9052, IN104[5], w9150, w9151);
  FullAdder U2995 (w9151, w9054, IN105[4], w9152, w9153);
  FullAdder U2996 (w9153, w9056, IN106[3], w9154, w9155);
  FullAdder U2997 (w9155, w9058, IN107[2], w9156, w9157);
  FullAdder U2998 (w9157, w9060, IN108[1], w9158, w9159);
  FullAdder U2999 (w9159, w9061, IN109[0], w9160, w9161);
  HalfAdder U3000 (w9064, IN61[49], Out1[61], w9163);
  FullAdder U3001 (w9163, w9066, IN62[48], Out1[62], w9165);
  FullAdder U3002 (w9165, w9068, IN63[47], Out1[63], w9167);
  FullAdder U3003 (w9167, w9070, IN64[46], Out1[64], w9169);
  FullAdder U3004 (w9169, w9072, IN65[45], Out1[65], w9171);
  FullAdder U3005 (w9171, w9074, IN66[44], Out1[66], w9173);
  FullAdder U3006 (w9173, w9076, IN67[43], Out1[67], w9175);
  FullAdder U3007 (w9175, w9078, IN68[42], Out1[68], w9177);
  FullAdder U3008 (w9177, w9080, IN69[41], Out1[69], w9179);
  FullAdder U3009 (w9179, w9082, IN70[40], Out1[70], w9181);
  FullAdder U3010 (w9181, w9084, IN71[39], Out1[71], w9183);
  FullAdder U3011 (w9183, w9086, IN72[38], Out1[72], w9185);
  FullAdder U3012 (w9185, w9088, IN73[37], Out1[73], w9187);
  FullAdder U3013 (w9187, w9090, IN74[36], Out1[74], w9189);
  FullAdder U3014 (w9189, w9092, IN75[35], Out1[75], w9191);
  FullAdder U3015 (w9191, w9094, IN76[34], Out1[76], w9193);
  FullAdder U3016 (w9193, w9096, IN77[33], Out1[77], w9195);
  FullAdder U3017 (w9195, w9098, IN78[32], Out1[78], w9197);
  FullAdder U3018 (w9197, w9100, IN79[31], Out1[79], w9199);
  FullAdder U3019 (w9199, w9102, IN80[30], Out1[80], w9201);
  FullAdder U3020 (w9201, w9104, IN81[29], Out1[81], w9203);
  FullAdder U3021 (w9203, w9106, IN82[28], Out1[82], w9205);
  FullAdder U3022 (w9205, w9108, IN83[27], Out1[83], w9207);
  FullAdder U3023 (w9207, w9110, IN84[26], Out1[84], w9209);
  FullAdder U3024 (w9209, w9112, IN85[25], Out1[85], w9211);
  FullAdder U3025 (w9211, w9114, IN86[24], Out1[86], w9213);
  FullAdder U3026 (w9213, w9116, IN87[23], Out1[87], w9215);
  FullAdder U3027 (w9215, w9118, IN88[22], Out1[88], w9217);
  FullAdder U3028 (w9217, w9120, IN89[21], Out1[89], w9219);
  FullAdder U3029 (w9219, w9122, IN90[20], Out1[90], w9221);
  FullAdder U3030 (w9221, w9124, IN91[19], Out1[91], w9223);
  FullAdder U3031 (w9223, w9126, IN92[18], Out1[92], w9225);
  FullAdder U3032 (w9225, w9128, IN93[17], Out1[93], w9227);
  FullAdder U3033 (w9227, w9130, IN94[16], Out1[94], w9229);
  FullAdder U3034 (w9229, w9132, IN95[15], Out1[95], w9231);
  FullAdder U3035 (w9231, w9134, IN96[14], Out1[96], w9233);
  FullAdder U3036 (w9233, w9136, IN97[13], Out1[97], w9235);
  FullAdder U3037 (w9235, w9138, IN98[12], Out1[98], w9237);
  FullAdder U3038 (w9237, w9140, IN99[11], Out1[99], w9239);
  FullAdder U3039 (w9239, w9142, IN100[10], Out1[100], w9241);
  FullAdder U3040 (w9241, w9144, IN101[9], Out1[101], w9243);
  FullAdder U3041 (w9243, w9146, IN102[8], Out1[102], w9245);
  FullAdder U3042 (w9245, w9148, IN103[7], Out1[103], w9247);
  FullAdder U3043 (w9247, w9150, IN104[6], Out1[104], w9249);
  FullAdder U3044 (w9249, w9152, IN105[5], Out1[105], w9251);
  FullAdder U3045 (w9251, w9154, IN106[4], Out1[106], w9253);
  FullAdder U3046 (w9253, w9156, IN107[3], Out1[107], w9255);
  FullAdder U3047 (w9255, w9158, IN108[2], Out1[108], w9257);
  FullAdder U3048 (w9257, w9160, IN109[1], Out1[109], w9259);
  FullAdder U3049 (w9259, w9161, IN110[0], Out1[110], Out1[111]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN51[50];
  assign Out2[1] = IN52[50];
  assign Out2[2] = IN53[50];
  assign Out2[3] = IN54[50];
  assign Out2[4] = IN55[50];
  assign Out2[5] = IN56[50];
  assign Out2[6] = IN57[50];
  assign Out2[7] = IN58[50];
  assign Out2[8] = IN59[50];
  assign Out2[9] = IN60[50];
  assign Out2[10] = IN61[50];
  assign Out2[11] = IN62[49];
  assign Out2[12] = IN63[48];
  assign Out2[13] = IN64[47];
  assign Out2[14] = IN65[46];
  assign Out2[15] = IN66[45];
  assign Out2[16] = IN67[44];
  assign Out2[17] = IN68[43];
  assign Out2[18] = IN69[42];
  assign Out2[19] = IN70[41];
  assign Out2[20] = IN71[40];
  assign Out2[21] = IN72[39];
  assign Out2[22] = IN73[38];
  assign Out2[23] = IN74[37];
  assign Out2[24] = IN75[36];
  assign Out2[25] = IN76[35];
  assign Out2[26] = IN77[34];
  assign Out2[27] = IN78[33];
  assign Out2[28] = IN79[32];
  assign Out2[29] = IN80[31];
  assign Out2[30] = IN81[30];
  assign Out2[31] = IN82[29];
  assign Out2[32] = IN83[28];
  assign Out2[33] = IN84[27];
  assign Out2[34] = IN85[26];
  assign Out2[35] = IN86[25];
  assign Out2[36] = IN87[24];
  assign Out2[37] = IN88[23];
  assign Out2[38] = IN89[22];
  assign Out2[39] = IN90[21];
  assign Out2[40] = IN91[20];
  assign Out2[41] = IN92[19];
  assign Out2[42] = IN93[18];
  assign Out2[43] = IN94[17];
  assign Out2[44] = IN95[16];
  assign Out2[45] = IN96[15];
  assign Out2[46] = IN97[14];
  assign Out2[47] = IN98[13];
  assign Out2[48] = IN99[12];
  assign Out2[49] = IN100[11];
  assign Out2[50] = IN101[10];
  assign Out2[51] = IN102[9];
  assign Out2[52] = IN103[8];
  assign Out2[53] = IN104[7];
  assign Out2[54] = IN105[6];
  assign Out2[55] = IN106[5];
  assign Out2[56] = IN107[4];
  assign Out2[57] = IN108[3];
  assign Out2[58] = IN109[2];
  assign Out2[59] = IN110[1];
  assign Out2[60] = IN111[0];

endmodule
module RC_61_61(IN1, IN2, Out);
  input [60:0] IN1;
  input [60:0] IN2;
  output [61:0] Out;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  wire w231;
  wire w233;
  wire w235;
  wire w237;
  wire w239;
  wire w241;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w123);
  FullAdder U1 (IN1[1], IN2[1], w123, Out[1], w125);
  FullAdder U2 (IN1[2], IN2[2], w125, Out[2], w127);
  FullAdder U3 (IN1[3], IN2[3], w127, Out[3], w129);
  FullAdder U4 (IN1[4], IN2[4], w129, Out[4], w131);
  FullAdder U5 (IN1[5], IN2[5], w131, Out[5], w133);
  FullAdder U6 (IN1[6], IN2[6], w133, Out[6], w135);
  FullAdder U7 (IN1[7], IN2[7], w135, Out[7], w137);
  FullAdder U8 (IN1[8], IN2[8], w137, Out[8], w139);
  FullAdder U9 (IN1[9], IN2[9], w139, Out[9], w141);
  FullAdder U10 (IN1[10], IN2[10], w141, Out[10], w143);
  FullAdder U11 (IN1[11], IN2[11], w143, Out[11], w145);
  FullAdder U12 (IN1[12], IN2[12], w145, Out[12], w147);
  FullAdder U13 (IN1[13], IN2[13], w147, Out[13], w149);
  FullAdder U14 (IN1[14], IN2[14], w149, Out[14], w151);
  FullAdder U15 (IN1[15], IN2[15], w151, Out[15], w153);
  FullAdder U16 (IN1[16], IN2[16], w153, Out[16], w155);
  FullAdder U17 (IN1[17], IN2[17], w155, Out[17], w157);
  FullAdder U18 (IN1[18], IN2[18], w157, Out[18], w159);
  FullAdder U19 (IN1[19], IN2[19], w159, Out[19], w161);
  FullAdder U20 (IN1[20], IN2[20], w161, Out[20], w163);
  FullAdder U21 (IN1[21], IN2[21], w163, Out[21], w165);
  FullAdder U22 (IN1[22], IN2[22], w165, Out[22], w167);
  FullAdder U23 (IN1[23], IN2[23], w167, Out[23], w169);
  FullAdder U24 (IN1[24], IN2[24], w169, Out[24], w171);
  FullAdder U25 (IN1[25], IN2[25], w171, Out[25], w173);
  FullAdder U26 (IN1[26], IN2[26], w173, Out[26], w175);
  FullAdder U27 (IN1[27], IN2[27], w175, Out[27], w177);
  FullAdder U28 (IN1[28], IN2[28], w177, Out[28], w179);
  FullAdder U29 (IN1[29], IN2[29], w179, Out[29], w181);
  FullAdder U30 (IN1[30], IN2[30], w181, Out[30], w183);
  FullAdder U31 (IN1[31], IN2[31], w183, Out[31], w185);
  FullAdder U32 (IN1[32], IN2[32], w185, Out[32], w187);
  FullAdder U33 (IN1[33], IN2[33], w187, Out[33], w189);
  FullAdder U34 (IN1[34], IN2[34], w189, Out[34], w191);
  FullAdder U35 (IN1[35], IN2[35], w191, Out[35], w193);
  FullAdder U36 (IN1[36], IN2[36], w193, Out[36], w195);
  FullAdder U37 (IN1[37], IN2[37], w195, Out[37], w197);
  FullAdder U38 (IN1[38], IN2[38], w197, Out[38], w199);
  FullAdder U39 (IN1[39], IN2[39], w199, Out[39], w201);
  FullAdder U40 (IN1[40], IN2[40], w201, Out[40], w203);
  FullAdder U41 (IN1[41], IN2[41], w203, Out[41], w205);
  FullAdder U42 (IN1[42], IN2[42], w205, Out[42], w207);
  FullAdder U43 (IN1[43], IN2[43], w207, Out[43], w209);
  FullAdder U44 (IN1[44], IN2[44], w209, Out[44], w211);
  FullAdder U45 (IN1[45], IN2[45], w211, Out[45], w213);
  FullAdder U46 (IN1[46], IN2[46], w213, Out[46], w215);
  FullAdder U47 (IN1[47], IN2[47], w215, Out[47], w217);
  FullAdder U48 (IN1[48], IN2[48], w217, Out[48], w219);
  FullAdder U49 (IN1[49], IN2[49], w219, Out[49], w221);
  FullAdder U50 (IN1[50], IN2[50], w221, Out[50], w223);
  FullAdder U51 (IN1[51], IN2[51], w223, Out[51], w225);
  FullAdder U52 (IN1[52], IN2[52], w225, Out[52], w227);
  FullAdder U53 (IN1[53], IN2[53], w227, Out[53], w229);
  FullAdder U54 (IN1[54], IN2[54], w229, Out[54], w231);
  FullAdder U55 (IN1[55], IN2[55], w231, Out[55], w233);
  FullAdder U56 (IN1[56], IN2[56], w233, Out[56], w235);
  FullAdder U57 (IN1[57], IN2[57], w235, Out[57], w237);
  FullAdder U58 (IN1[58], IN2[58], w237, Out[58], w239);
  FullAdder U59 (IN1[59], IN2[59], w239, Out[59], w241);
  FullAdder U60 (IN1[60], IN2[60], w241, Out[60], Out[61]);

endmodule
module NR_51_62(IN1, IN2, Out);
  input [50:0] IN1;
  input [61:0] IN2;
  output [112:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [29:0] P29;
  wire [30:0] P30;
  wire [31:0] P31;
  wire [32:0] P32;
  wire [33:0] P33;
  wire [34:0] P34;
  wire [35:0] P35;
  wire [36:0] P36;
  wire [37:0] P37;
  wire [38:0] P38;
  wire [39:0] P39;
  wire [40:0] P40;
  wire [41:0] P41;
  wire [42:0] P42;
  wire [43:0] P43;
  wire [44:0] P44;
  wire [45:0] P45;
  wire [46:0] P46;
  wire [47:0] P47;
  wire [48:0] P48;
  wire [49:0] P49;
  wire [50:0] P50;
  wire [50:0] P51;
  wire [50:0] P52;
  wire [50:0] P53;
  wire [50:0] P54;
  wire [50:0] P55;
  wire [50:0] P56;
  wire [50:0] P57;
  wire [50:0] P58;
  wire [50:0] P59;
  wire [50:0] P60;
  wire [50:0] P61;
  wire [49:0] P62;
  wire [48:0] P63;
  wire [47:0] P64;
  wire [46:0] P65;
  wire [45:0] P66;
  wire [44:0] P67;
  wire [43:0] P68;
  wire [42:0] P69;
  wire [41:0] P70;
  wire [40:0] P71;
  wire [39:0] P72;
  wire [38:0] P73;
  wire [37:0] P74;
  wire [36:0] P75;
  wire [35:0] P76;
  wire [34:0] P77;
  wire [33:0] P78;
  wire [32:0] P79;
  wire [31:0] P80;
  wire [30:0] P81;
  wire [29:0] P82;
  wire [28:0] P83;
  wire [27:0] P84;
  wire [26:0] P85;
  wire [25:0] P86;
  wire [24:0] P87;
  wire [23:0] P88;
  wire [22:0] P89;
  wire [21:0] P90;
  wire [20:0] P91;
  wire [19:0] P92;
  wire [18:0] P93;
  wire [17:0] P94;
  wire [16:0] P95;
  wire [15:0] P96;
  wire [14:0] P97;
  wire [13:0] P98;
  wire [12:0] P99;
  wire [11:0] P100;
  wire [10:0] P101;
  wire [9:0] P102;
  wire [8:0] P103;
  wire [7:0] P104;
  wire [6:0] P105;
  wire [5:0] P106;
  wire [4:0] P107;
  wire [3:0] P108;
  wire [2:0] P109;
  wire [1:0] P110;
  wire [0:0] P111;
  wire [111:0] R1;
  wire [60:0] R2;
  wire [112:0] aOut;
  U_SP_51_62 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, R1, R2);
  RC_61_61 S2 (R1[111:51], R2, aOut[112:51]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign Out = aOut[112:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
