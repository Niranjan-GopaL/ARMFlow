//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 33
  second input length: 6
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_33_6(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37);
  input [32:0] IN1;
  input [5:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [5:0] P6;
  output [5:0] P7;
  output [5:0] P8;
  output [5:0] P9;
  output [5:0] P10;
  output [5:0] P11;
  output [5:0] P12;
  output [5:0] P13;
  output [5:0] P14;
  output [5:0] P15;
  output [5:0] P16;
  output [5:0] P17;
  output [5:0] P18;
  output [5:0] P19;
  output [5:0] P20;
  output [5:0] P21;
  output [5:0] P22;
  output [5:0] P23;
  output [5:0] P24;
  output [5:0] P25;
  output [5:0] P26;
  output [5:0] P27;
  output [5:0] P28;
  output [5:0] P29;
  output [5:0] P30;
  output [5:0] P31;
  output [5:0] P32;
  output [4:0] P33;
  output [3:0] P34;
  output [2:0] P35;
  output [1:0] P36;
  output [0:0] P37;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[0] = IN1[1]&IN2[5];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[1] = IN1[2]&IN2[4];
  assign P7[0] = IN1[2]&IN2[5];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[2] = IN1[3]&IN2[3];
  assign P7[1] = IN1[3]&IN2[4];
  assign P8[0] = IN1[3]&IN2[5];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[3] = IN1[4]&IN2[2];
  assign P7[2] = IN1[4]&IN2[3];
  assign P8[1] = IN1[4]&IN2[4];
  assign P9[0] = IN1[4]&IN2[5];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[4] = IN1[5]&IN2[1];
  assign P7[3] = IN1[5]&IN2[2];
  assign P8[2] = IN1[5]&IN2[3];
  assign P9[1] = IN1[5]&IN2[4];
  assign P10[0] = IN1[5]&IN2[5];
  assign P6[5] = IN1[6]&IN2[0];
  assign P7[4] = IN1[6]&IN2[1];
  assign P8[3] = IN1[6]&IN2[2];
  assign P9[2] = IN1[6]&IN2[3];
  assign P10[1] = IN1[6]&IN2[4];
  assign P11[0] = IN1[6]&IN2[5];
  assign P7[5] = IN1[7]&IN2[0];
  assign P8[4] = IN1[7]&IN2[1];
  assign P9[3] = IN1[7]&IN2[2];
  assign P10[2] = IN1[7]&IN2[3];
  assign P11[1] = IN1[7]&IN2[4];
  assign P12[0] = IN1[7]&IN2[5];
  assign P8[5] = IN1[8]&IN2[0];
  assign P9[4] = IN1[8]&IN2[1];
  assign P10[3] = IN1[8]&IN2[2];
  assign P11[2] = IN1[8]&IN2[3];
  assign P12[1] = IN1[8]&IN2[4];
  assign P13[0] = IN1[8]&IN2[5];
  assign P9[5] = IN1[9]&IN2[0];
  assign P10[4] = IN1[9]&IN2[1];
  assign P11[3] = IN1[9]&IN2[2];
  assign P12[2] = IN1[9]&IN2[3];
  assign P13[1] = IN1[9]&IN2[4];
  assign P14[0] = IN1[9]&IN2[5];
  assign P10[5] = IN1[10]&IN2[0];
  assign P11[4] = IN1[10]&IN2[1];
  assign P12[3] = IN1[10]&IN2[2];
  assign P13[2] = IN1[10]&IN2[3];
  assign P14[1] = IN1[10]&IN2[4];
  assign P15[0] = IN1[10]&IN2[5];
  assign P11[5] = IN1[11]&IN2[0];
  assign P12[4] = IN1[11]&IN2[1];
  assign P13[3] = IN1[11]&IN2[2];
  assign P14[2] = IN1[11]&IN2[3];
  assign P15[1] = IN1[11]&IN2[4];
  assign P16[0] = IN1[11]&IN2[5];
  assign P12[5] = IN1[12]&IN2[0];
  assign P13[4] = IN1[12]&IN2[1];
  assign P14[3] = IN1[12]&IN2[2];
  assign P15[2] = IN1[12]&IN2[3];
  assign P16[1] = IN1[12]&IN2[4];
  assign P17[0] = IN1[12]&IN2[5];
  assign P13[5] = IN1[13]&IN2[0];
  assign P14[4] = IN1[13]&IN2[1];
  assign P15[3] = IN1[13]&IN2[2];
  assign P16[2] = IN1[13]&IN2[3];
  assign P17[1] = IN1[13]&IN2[4];
  assign P18[0] = IN1[13]&IN2[5];
  assign P14[5] = IN1[14]&IN2[0];
  assign P15[4] = IN1[14]&IN2[1];
  assign P16[3] = IN1[14]&IN2[2];
  assign P17[2] = IN1[14]&IN2[3];
  assign P18[1] = IN1[14]&IN2[4];
  assign P19[0] = IN1[14]&IN2[5];
  assign P15[5] = IN1[15]&IN2[0];
  assign P16[4] = IN1[15]&IN2[1];
  assign P17[3] = IN1[15]&IN2[2];
  assign P18[2] = IN1[15]&IN2[3];
  assign P19[1] = IN1[15]&IN2[4];
  assign P20[0] = IN1[15]&IN2[5];
  assign P16[5] = IN1[16]&IN2[0];
  assign P17[4] = IN1[16]&IN2[1];
  assign P18[3] = IN1[16]&IN2[2];
  assign P19[2] = IN1[16]&IN2[3];
  assign P20[1] = IN1[16]&IN2[4];
  assign P21[0] = IN1[16]&IN2[5];
  assign P17[5] = IN1[17]&IN2[0];
  assign P18[4] = IN1[17]&IN2[1];
  assign P19[3] = IN1[17]&IN2[2];
  assign P20[2] = IN1[17]&IN2[3];
  assign P21[1] = IN1[17]&IN2[4];
  assign P22[0] = IN1[17]&IN2[5];
  assign P18[5] = IN1[18]&IN2[0];
  assign P19[4] = IN1[18]&IN2[1];
  assign P20[3] = IN1[18]&IN2[2];
  assign P21[2] = IN1[18]&IN2[3];
  assign P22[1] = IN1[18]&IN2[4];
  assign P23[0] = IN1[18]&IN2[5];
  assign P19[5] = IN1[19]&IN2[0];
  assign P20[4] = IN1[19]&IN2[1];
  assign P21[3] = IN1[19]&IN2[2];
  assign P22[2] = IN1[19]&IN2[3];
  assign P23[1] = IN1[19]&IN2[4];
  assign P24[0] = IN1[19]&IN2[5];
  assign P20[5] = IN1[20]&IN2[0];
  assign P21[4] = IN1[20]&IN2[1];
  assign P22[3] = IN1[20]&IN2[2];
  assign P23[2] = IN1[20]&IN2[3];
  assign P24[1] = IN1[20]&IN2[4];
  assign P25[0] = IN1[20]&IN2[5];
  assign P21[5] = IN1[21]&IN2[0];
  assign P22[4] = IN1[21]&IN2[1];
  assign P23[3] = IN1[21]&IN2[2];
  assign P24[2] = IN1[21]&IN2[3];
  assign P25[1] = IN1[21]&IN2[4];
  assign P26[0] = IN1[21]&IN2[5];
  assign P22[5] = IN1[22]&IN2[0];
  assign P23[4] = IN1[22]&IN2[1];
  assign P24[3] = IN1[22]&IN2[2];
  assign P25[2] = IN1[22]&IN2[3];
  assign P26[1] = IN1[22]&IN2[4];
  assign P27[0] = IN1[22]&IN2[5];
  assign P23[5] = IN1[23]&IN2[0];
  assign P24[4] = IN1[23]&IN2[1];
  assign P25[3] = IN1[23]&IN2[2];
  assign P26[2] = IN1[23]&IN2[3];
  assign P27[1] = IN1[23]&IN2[4];
  assign P28[0] = IN1[23]&IN2[5];
  assign P24[5] = IN1[24]&IN2[0];
  assign P25[4] = IN1[24]&IN2[1];
  assign P26[3] = IN1[24]&IN2[2];
  assign P27[2] = IN1[24]&IN2[3];
  assign P28[1] = IN1[24]&IN2[4];
  assign P29[0] = IN1[24]&IN2[5];
  assign P25[5] = IN1[25]&IN2[0];
  assign P26[4] = IN1[25]&IN2[1];
  assign P27[3] = IN1[25]&IN2[2];
  assign P28[2] = IN1[25]&IN2[3];
  assign P29[1] = IN1[25]&IN2[4];
  assign P30[0] = IN1[25]&IN2[5];
  assign P26[5] = IN1[26]&IN2[0];
  assign P27[4] = IN1[26]&IN2[1];
  assign P28[3] = IN1[26]&IN2[2];
  assign P29[2] = IN1[26]&IN2[3];
  assign P30[1] = IN1[26]&IN2[4];
  assign P31[0] = IN1[26]&IN2[5];
  assign P27[5] = IN1[27]&IN2[0];
  assign P28[4] = IN1[27]&IN2[1];
  assign P29[3] = IN1[27]&IN2[2];
  assign P30[2] = IN1[27]&IN2[3];
  assign P31[1] = IN1[27]&IN2[4];
  assign P32[0] = IN1[27]&IN2[5];
  assign P28[5] = IN1[28]&IN2[0];
  assign P29[4] = IN1[28]&IN2[1];
  assign P30[3] = IN1[28]&IN2[2];
  assign P31[2] = IN1[28]&IN2[3];
  assign P32[1] = IN1[28]&IN2[4];
  assign P33[0] = IN1[28]&IN2[5];
  assign P29[5] = IN1[29]&IN2[0];
  assign P30[4] = IN1[29]&IN2[1];
  assign P31[3] = IN1[29]&IN2[2];
  assign P32[2] = IN1[29]&IN2[3];
  assign P33[1] = IN1[29]&IN2[4];
  assign P34[0] = IN1[29]&IN2[5];
  assign P30[5] = IN1[30]&IN2[0];
  assign P31[4] = IN1[30]&IN2[1];
  assign P32[3] = IN1[30]&IN2[2];
  assign P33[2] = IN1[30]&IN2[3];
  assign P34[1] = IN1[30]&IN2[4];
  assign P35[0] = IN1[30]&IN2[5];
  assign P31[5] = IN1[31]&IN2[0];
  assign P32[4] = IN1[31]&IN2[1];
  assign P33[3] = IN1[31]&IN2[2];
  assign P34[2] = IN1[31]&IN2[3];
  assign P35[1] = IN1[31]&IN2[4];
  assign P36[0] = IN1[31]&IN2[5];
  assign P32[5] = IN1[32]&IN2[0];
  assign P33[4] = IN1[32]&IN2[1];
  assign P34[3] = IN1[32]&IN2[2];
  assign P35[2] = IN1[32]&IN2[3];
  assign P36[1] = IN1[32]&IN2[4];
  assign P37[0] = IN1[32]&IN2[5];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [5:0] IN6;
  input [5:0] IN7;
  input [5:0] IN8;
  input [5:0] IN9;
  input [5:0] IN10;
  input [5:0] IN11;
  input [5:0] IN12;
  input [5:0] IN13;
  input [5:0] IN14;
  input [5:0] IN15;
  input [5:0] IN16;
  input [5:0] IN17;
  input [5:0] IN18;
  input [5:0] IN19;
  input [5:0] IN20;
  input [5:0] IN21;
  input [5:0] IN22;
  input [5:0] IN23;
  input [5:0] IN24;
  input [5:0] IN25;
  input [5:0] IN26;
  input [5:0] IN27;
  input [5:0] IN28;
  input [5:0] IN29;
  input [5:0] IN30;
  input [5:0] IN31;
  input [5:0] IN32;
  input [4:0] IN33;
  input [3:0] IN34;
  input [2:0] IN35;
  input [1:0] IN36;
  input [0:0] IN37;
  output [37:0] Out1;
  output [4:0] Out2;
  wire w199;
  wire w200;
  wire w201;
  wire w202;
  wire w203;
  wire w204;
  wire w205;
  wire w206;
  wire w207;
  wire w208;
  wire w209;
  wire w210;
  wire w211;
  wire w212;
  wire w213;
  wire w214;
  wire w215;
  wire w216;
  wire w217;
  wire w218;
  wire w219;
  wire w220;
  wire w221;
  wire w222;
  wire w223;
  wire w224;
  wire w225;
  wire w226;
  wire w227;
  wire w228;
  wire w229;
  wire w230;
  wire w231;
  wire w232;
  wire w233;
  wire w234;
  wire w235;
  wire w236;
  wire w237;
  wire w238;
  wire w239;
  wire w240;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w246;
  wire w247;
  wire w248;
  wire w249;
  wire w250;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w455;
  wire w457;
  wire w459;
  wire w461;
  wire w463;
  wire w465;
  wire w467;
  wire w469;
  wire w471;
  wire w473;
  wire w475;
  wire w477;
  wire w479;
  wire w481;
  wire w483;
  wire w485;
  wire w487;
  wire w489;
  wire w491;
  wire w493;
  wire w495;
  wire w497;
  wire w499;
  wire w501;
  wire w503;
  wire w505;
  wire w507;
  wire w509;
  wire w511;
  wire w513;
  wire w515;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w199);
  FullAdder U1 (w199, IN2[0], IN2[1], w200, w201);
  FullAdder U2 (w201, IN3[0], IN3[1], w202, w203);
  FullAdder U3 (w203, IN4[0], IN4[1], w204, w205);
  FullAdder U4 (w205, IN5[0], IN5[1], w206, w207);
  FullAdder U5 (w207, IN6[0], IN6[1], w208, w209);
  FullAdder U6 (w209, IN7[0], IN7[1], w210, w211);
  FullAdder U7 (w211, IN8[0], IN8[1], w212, w213);
  FullAdder U8 (w213, IN9[0], IN9[1], w214, w215);
  FullAdder U9 (w215, IN10[0], IN10[1], w216, w217);
  FullAdder U10 (w217, IN11[0], IN11[1], w218, w219);
  FullAdder U11 (w219, IN12[0], IN12[1], w220, w221);
  FullAdder U12 (w221, IN13[0], IN13[1], w222, w223);
  FullAdder U13 (w223, IN14[0], IN14[1], w224, w225);
  FullAdder U14 (w225, IN15[0], IN15[1], w226, w227);
  FullAdder U15 (w227, IN16[0], IN16[1], w228, w229);
  FullAdder U16 (w229, IN17[0], IN17[1], w230, w231);
  FullAdder U17 (w231, IN18[0], IN18[1], w232, w233);
  FullAdder U18 (w233, IN19[0], IN19[1], w234, w235);
  FullAdder U19 (w235, IN20[0], IN20[1], w236, w237);
  FullAdder U20 (w237, IN21[0], IN21[1], w238, w239);
  FullAdder U21 (w239, IN22[0], IN22[1], w240, w241);
  FullAdder U22 (w241, IN23[0], IN23[1], w242, w243);
  FullAdder U23 (w243, IN24[0], IN24[1], w244, w245);
  FullAdder U24 (w245, IN25[0], IN25[1], w246, w247);
  FullAdder U25 (w247, IN26[0], IN26[1], w248, w249);
  FullAdder U26 (w249, IN27[0], IN27[1], w250, w251);
  FullAdder U27 (w251, IN28[0], IN28[1], w252, w253);
  FullAdder U28 (w253, IN29[0], IN29[1], w254, w255);
  FullAdder U29 (w255, IN30[0], IN30[1], w256, w257);
  FullAdder U30 (w257, IN31[0], IN31[1], w258, w259);
  FullAdder U31 (w259, IN32[0], IN32[1], w260, w261);
  HalfAdder U32 (w200, IN2[2], Out1[2], w263);
  FullAdder U33 (w263, w202, IN3[2], w264, w265);
  FullAdder U34 (w265, w204, IN4[2], w266, w267);
  FullAdder U35 (w267, w206, IN5[2], w268, w269);
  FullAdder U36 (w269, w208, IN6[2], w270, w271);
  FullAdder U37 (w271, w210, IN7[2], w272, w273);
  FullAdder U38 (w273, w212, IN8[2], w274, w275);
  FullAdder U39 (w275, w214, IN9[2], w276, w277);
  FullAdder U40 (w277, w216, IN10[2], w278, w279);
  FullAdder U41 (w279, w218, IN11[2], w280, w281);
  FullAdder U42 (w281, w220, IN12[2], w282, w283);
  FullAdder U43 (w283, w222, IN13[2], w284, w285);
  FullAdder U44 (w285, w224, IN14[2], w286, w287);
  FullAdder U45 (w287, w226, IN15[2], w288, w289);
  FullAdder U46 (w289, w228, IN16[2], w290, w291);
  FullAdder U47 (w291, w230, IN17[2], w292, w293);
  FullAdder U48 (w293, w232, IN18[2], w294, w295);
  FullAdder U49 (w295, w234, IN19[2], w296, w297);
  FullAdder U50 (w297, w236, IN20[2], w298, w299);
  FullAdder U51 (w299, w238, IN21[2], w300, w301);
  FullAdder U52 (w301, w240, IN22[2], w302, w303);
  FullAdder U53 (w303, w242, IN23[2], w304, w305);
  FullAdder U54 (w305, w244, IN24[2], w306, w307);
  FullAdder U55 (w307, w246, IN25[2], w308, w309);
  FullAdder U56 (w309, w248, IN26[2], w310, w311);
  FullAdder U57 (w311, w250, IN27[2], w312, w313);
  FullAdder U58 (w313, w252, IN28[2], w314, w315);
  FullAdder U59 (w315, w254, IN29[2], w316, w317);
  FullAdder U60 (w317, w256, IN30[2], w318, w319);
  FullAdder U61 (w319, w258, IN31[2], w320, w321);
  FullAdder U62 (w321, w260, IN32[2], w322, w323);
  FullAdder U63 (w323, w261, IN33[0], w324, w325);
  HalfAdder U64 (w264, IN3[3], Out1[3], w327);
  FullAdder U65 (w327, w266, IN4[3], w328, w329);
  FullAdder U66 (w329, w268, IN5[3], w330, w331);
  FullAdder U67 (w331, w270, IN6[3], w332, w333);
  FullAdder U68 (w333, w272, IN7[3], w334, w335);
  FullAdder U69 (w335, w274, IN8[3], w336, w337);
  FullAdder U70 (w337, w276, IN9[3], w338, w339);
  FullAdder U71 (w339, w278, IN10[3], w340, w341);
  FullAdder U72 (w341, w280, IN11[3], w342, w343);
  FullAdder U73 (w343, w282, IN12[3], w344, w345);
  FullAdder U74 (w345, w284, IN13[3], w346, w347);
  FullAdder U75 (w347, w286, IN14[3], w348, w349);
  FullAdder U76 (w349, w288, IN15[3], w350, w351);
  FullAdder U77 (w351, w290, IN16[3], w352, w353);
  FullAdder U78 (w353, w292, IN17[3], w354, w355);
  FullAdder U79 (w355, w294, IN18[3], w356, w357);
  FullAdder U80 (w357, w296, IN19[3], w358, w359);
  FullAdder U81 (w359, w298, IN20[3], w360, w361);
  FullAdder U82 (w361, w300, IN21[3], w362, w363);
  FullAdder U83 (w363, w302, IN22[3], w364, w365);
  FullAdder U84 (w365, w304, IN23[3], w366, w367);
  FullAdder U85 (w367, w306, IN24[3], w368, w369);
  FullAdder U86 (w369, w308, IN25[3], w370, w371);
  FullAdder U87 (w371, w310, IN26[3], w372, w373);
  FullAdder U88 (w373, w312, IN27[3], w374, w375);
  FullAdder U89 (w375, w314, IN28[3], w376, w377);
  FullAdder U90 (w377, w316, IN29[3], w378, w379);
  FullAdder U91 (w379, w318, IN30[3], w380, w381);
  FullAdder U92 (w381, w320, IN31[3], w382, w383);
  FullAdder U93 (w383, w322, IN32[3], w384, w385);
  FullAdder U94 (w385, w324, IN33[1], w386, w387);
  FullAdder U95 (w387, w325, IN34[0], w388, w389);
  HalfAdder U96 (w328, IN4[4], Out1[4], w391);
  FullAdder U97 (w391, w330, IN5[4], w392, w393);
  FullAdder U98 (w393, w332, IN6[4], w394, w395);
  FullAdder U99 (w395, w334, IN7[4], w396, w397);
  FullAdder U100 (w397, w336, IN8[4], w398, w399);
  FullAdder U101 (w399, w338, IN9[4], w400, w401);
  FullAdder U102 (w401, w340, IN10[4], w402, w403);
  FullAdder U103 (w403, w342, IN11[4], w404, w405);
  FullAdder U104 (w405, w344, IN12[4], w406, w407);
  FullAdder U105 (w407, w346, IN13[4], w408, w409);
  FullAdder U106 (w409, w348, IN14[4], w410, w411);
  FullAdder U107 (w411, w350, IN15[4], w412, w413);
  FullAdder U108 (w413, w352, IN16[4], w414, w415);
  FullAdder U109 (w415, w354, IN17[4], w416, w417);
  FullAdder U110 (w417, w356, IN18[4], w418, w419);
  FullAdder U111 (w419, w358, IN19[4], w420, w421);
  FullAdder U112 (w421, w360, IN20[4], w422, w423);
  FullAdder U113 (w423, w362, IN21[4], w424, w425);
  FullAdder U114 (w425, w364, IN22[4], w426, w427);
  FullAdder U115 (w427, w366, IN23[4], w428, w429);
  FullAdder U116 (w429, w368, IN24[4], w430, w431);
  FullAdder U117 (w431, w370, IN25[4], w432, w433);
  FullAdder U118 (w433, w372, IN26[4], w434, w435);
  FullAdder U119 (w435, w374, IN27[4], w436, w437);
  FullAdder U120 (w437, w376, IN28[4], w438, w439);
  FullAdder U121 (w439, w378, IN29[4], w440, w441);
  FullAdder U122 (w441, w380, IN30[4], w442, w443);
  FullAdder U123 (w443, w382, IN31[4], w444, w445);
  FullAdder U124 (w445, w384, IN32[4], w446, w447);
  FullAdder U125 (w447, w386, IN33[2], w448, w449);
  FullAdder U126 (w449, w388, IN34[1], w450, w451);
  FullAdder U127 (w451, w389, IN35[0], w452, w453);
  HalfAdder U128 (w392, IN5[5], Out1[5], w455);
  FullAdder U129 (w455, w394, IN6[5], Out1[6], w457);
  FullAdder U130 (w457, w396, IN7[5], Out1[7], w459);
  FullAdder U131 (w459, w398, IN8[5], Out1[8], w461);
  FullAdder U132 (w461, w400, IN9[5], Out1[9], w463);
  FullAdder U133 (w463, w402, IN10[5], Out1[10], w465);
  FullAdder U134 (w465, w404, IN11[5], Out1[11], w467);
  FullAdder U135 (w467, w406, IN12[5], Out1[12], w469);
  FullAdder U136 (w469, w408, IN13[5], Out1[13], w471);
  FullAdder U137 (w471, w410, IN14[5], Out1[14], w473);
  FullAdder U138 (w473, w412, IN15[5], Out1[15], w475);
  FullAdder U139 (w475, w414, IN16[5], Out1[16], w477);
  FullAdder U140 (w477, w416, IN17[5], Out1[17], w479);
  FullAdder U141 (w479, w418, IN18[5], Out1[18], w481);
  FullAdder U142 (w481, w420, IN19[5], Out1[19], w483);
  FullAdder U143 (w483, w422, IN20[5], Out1[20], w485);
  FullAdder U144 (w485, w424, IN21[5], Out1[21], w487);
  FullAdder U145 (w487, w426, IN22[5], Out1[22], w489);
  FullAdder U146 (w489, w428, IN23[5], Out1[23], w491);
  FullAdder U147 (w491, w430, IN24[5], Out1[24], w493);
  FullAdder U148 (w493, w432, IN25[5], Out1[25], w495);
  FullAdder U149 (w495, w434, IN26[5], Out1[26], w497);
  FullAdder U150 (w497, w436, IN27[5], Out1[27], w499);
  FullAdder U151 (w499, w438, IN28[5], Out1[28], w501);
  FullAdder U152 (w501, w440, IN29[5], Out1[29], w503);
  FullAdder U153 (w503, w442, IN30[5], Out1[30], w505);
  FullAdder U154 (w505, w444, IN31[5], Out1[31], w507);
  FullAdder U155 (w507, w446, IN32[5], Out1[32], w509);
  FullAdder U156 (w509, w448, IN33[3], Out1[33], w511);
  FullAdder U157 (w511, w450, IN34[2], Out1[34], w513);
  FullAdder U158 (w513, w452, IN35[1], Out1[35], w515);
  FullAdder U159 (w515, w453, IN36[0], Out1[36], Out1[37]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN33[4];
  assign Out2[1] = IN34[3];
  assign Out2[2] = IN35[2];
  assign Out2[3] = IN36[1];
  assign Out2[4] = IN37[0];

endmodule
module RC_5_5(IN1, IN2, Out);
  input [4:0] IN1;
  input [4:0] IN2;
  output [5:0] Out;
  wire w11;
  wire w13;
  wire w15;
  wire w17;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w11);
  FullAdder U1 (IN1[1], IN2[1], w11, Out[1], w13);
  FullAdder U2 (IN1[2], IN2[2], w13, Out[2], w15);
  FullAdder U3 (IN1[3], IN2[3], w15, Out[3], w17);
  FullAdder U4 (IN1[4], IN2[4], w17, Out[4], Out[5]);

endmodule
module NR_33_6(IN1, IN2, Out);
  input [32:0] IN1;
  input [5:0] IN2;
  output [38:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [5:0] P6;
  wire [5:0] P7;
  wire [5:0] P8;
  wire [5:0] P9;
  wire [5:0] P10;
  wire [5:0] P11;
  wire [5:0] P12;
  wire [5:0] P13;
  wire [5:0] P14;
  wire [5:0] P15;
  wire [5:0] P16;
  wire [5:0] P17;
  wire [5:0] P18;
  wire [5:0] P19;
  wire [5:0] P20;
  wire [5:0] P21;
  wire [5:0] P22;
  wire [5:0] P23;
  wire [5:0] P24;
  wire [5:0] P25;
  wire [5:0] P26;
  wire [5:0] P27;
  wire [5:0] P28;
  wire [5:0] P29;
  wire [5:0] P30;
  wire [5:0] P31;
  wire [5:0] P32;
  wire [4:0] P33;
  wire [3:0] P34;
  wire [2:0] P35;
  wire [1:0] P36;
  wire [0:0] P37;
  wire [37:0] R1;
  wire [4:0] R2;
  wire [38:0] aOut;
  U_SP_33_6 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, R1, R2);
  RC_5_5 S2 (R1[37:33], R2, aOut[38:33]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign Out = aOut[38:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
