//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 57
  second input length: 5
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_57_5(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60);
  input [56:0] IN1;
  input [4:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [4:0] P5;
  output [4:0] P6;
  output [4:0] P7;
  output [4:0] P8;
  output [4:0] P9;
  output [4:0] P10;
  output [4:0] P11;
  output [4:0] P12;
  output [4:0] P13;
  output [4:0] P14;
  output [4:0] P15;
  output [4:0] P16;
  output [4:0] P17;
  output [4:0] P18;
  output [4:0] P19;
  output [4:0] P20;
  output [4:0] P21;
  output [4:0] P22;
  output [4:0] P23;
  output [4:0] P24;
  output [4:0] P25;
  output [4:0] P26;
  output [4:0] P27;
  output [4:0] P28;
  output [4:0] P29;
  output [4:0] P30;
  output [4:0] P31;
  output [4:0] P32;
  output [4:0] P33;
  output [4:0] P34;
  output [4:0] P35;
  output [4:0] P36;
  output [4:0] P37;
  output [4:0] P38;
  output [4:0] P39;
  output [4:0] P40;
  output [4:0] P41;
  output [4:0] P42;
  output [4:0] P43;
  output [4:0] P44;
  output [4:0] P45;
  output [4:0] P46;
  output [4:0] P47;
  output [4:0] P48;
  output [4:0] P49;
  output [4:0] P50;
  output [4:0] P51;
  output [4:0] P52;
  output [4:0] P53;
  output [4:0] P54;
  output [4:0] P55;
  output [4:0] P56;
  output [3:0] P57;
  output [2:0] P58;
  output [1:0] P59;
  output [0:0] P60;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[0] = IN1[1]&IN2[4];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[1] = IN1[2]&IN2[3];
  assign P6[0] = IN1[2]&IN2[4];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[2] = IN1[3]&IN2[2];
  assign P6[1] = IN1[3]&IN2[3];
  assign P7[0] = IN1[3]&IN2[4];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[3] = IN1[4]&IN2[1];
  assign P6[2] = IN1[4]&IN2[2];
  assign P7[1] = IN1[4]&IN2[3];
  assign P8[0] = IN1[4]&IN2[4];
  assign P5[4] = IN1[5]&IN2[0];
  assign P6[3] = IN1[5]&IN2[1];
  assign P7[2] = IN1[5]&IN2[2];
  assign P8[1] = IN1[5]&IN2[3];
  assign P9[0] = IN1[5]&IN2[4];
  assign P6[4] = IN1[6]&IN2[0];
  assign P7[3] = IN1[6]&IN2[1];
  assign P8[2] = IN1[6]&IN2[2];
  assign P9[1] = IN1[6]&IN2[3];
  assign P10[0] = IN1[6]&IN2[4];
  assign P7[4] = IN1[7]&IN2[0];
  assign P8[3] = IN1[7]&IN2[1];
  assign P9[2] = IN1[7]&IN2[2];
  assign P10[1] = IN1[7]&IN2[3];
  assign P11[0] = IN1[7]&IN2[4];
  assign P8[4] = IN1[8]&IN2[0];
  assign P9[3] = IN1[8]&IN2[1];
  assign P10[2] = IN1[8]&IN2[2];
  assign P11[1] = IN1[8]&IN2[3];
  assign P12[0] = IN1[8]&IN2[4];
  assign P9[4] = IN1[9]&IN2[0];
  assign P10[3] = IN1[9]&IN2[1];
  assign P11[2] = IN1[9]&IN2[2];
  assign P12[1] = IN1[9]&IN2[3];
  assign P13[0] = IN1[9]&IN2[4];
  assign P10[4] = IN1[10]&IN2[0];
  assign P11[3] = IN1[10]&IN2[1];
  assign P12[2] = IN1[10]&IN2[2];
  assign P13[1] = IN1[10]&IN2[3];
  assign P14[0] = IN1[10]&IN2[4];
  assign P11[4] = IN1[11]&IN2[0];
  assign P12[3] = IN1[11]&IN2[1];
  assign P13[2] = IN1[11]&IN2[2];
  assign P14[1] = IN1[11]&IN2[3];
  assign P15[0] = IN1[11]&IN2[4];
  assign P12[4] = IN1[12]&IN2[0];
  assign P13[3] = IN1[12]&IN2[1];
  assign P14[2] = IN1[12]&IN2[2];
  assign P15[1] = IN1[12]&IN2[3];
  assign P16[0] = IN1[12]&IN2[4];
  assign P13[4] = IN1[13]&IN2[0];
  assign P14[3] = IN1[13]&IN2[1];
  assign P15[2] = IN1[13]&IN2[2];
  assign P16[1] = IN1[13]&IN2[3];
  assign P17[0] = IN1[13]&IN2[4];
  assign P14[4] = IN1[14]&IN2[0];
  assign P15[3] = IN1[14]&IN2[1];
  assign P16[2] = IN1[14]&IN2[2];
  assign P17[1] = IN1[14]&IN2[3];
  assign P18[0] = IN1[14]&IN2[4];
  assign P15[4] = IN1[15]&IN2[0];
  assign P16[3] = IN1[15]&IN2[1];
  assign P17[2] = IN1[15]&IN2[2];
  assign P18[1] = IN1[15]&IN2[3];
  assign P19[0] = IN1[15]&IN2[4];
  assign P16[4] = IN1[16]&IN2[0];
  assign P17[3] = IN1[16]&IN2[1];
  assign P18[2] = IN1[16]&IN2[2];
  assign P19[1] = IN1[16]&IN2[3];
  assign P20[0] = IN1[16]&IN2[4];
  assign P17[4] = IN1[17]&IN2[0];
  assign P18[3] = IN1[17]&IN2[1];
  assign P19[2] = IN1[17]&IN2[2];
  assign P20[1] = IN1[17]&IN2[3];
  assign P21[0] = IN1[17]&IN2[4];
  assign P18[4] = IN1[18]&IN2[0];
  assign P19[3] = IN1[18]&IN2[1];
  assign P20[2] = IN1[18]&IN2[2];
  assign P21[1] = IN1[18]&IN2[3];
  assign P22[0] = IN1[18]&IN2[4];
  assign P19[4] = IN1[19]&IN2[0];
  assign P20[3] = IN1[19]&IN2[1];
  assign P21[2] = IN1[19]&IN2[2];
  assign P22[1] = IN1[19]&IN2[3];
  assign P23[0] = IN1[19]&IN2[4];
  assign P20[4] = IN1[20]&IN2[0];
  assign P21[3] = IN1[20]&IN2[1];
  assign P22[2] = IN1[20]&IN2[2];
  assign P23[1] = IN1[20]&IN2[3];
  assign P24[0] = IN1[20]&IN2[4];
  assign P21[4] = IN1[21]&IN2[0];
  assign P22[3] = IN1[21]&IN2[1];
  assign P23[2] = IN1[21]&IN2[2];
  assign P24[1] = IN1[21]&IN2[3];
  assign P25[0] = IN1[21]&IN2[4];
  assign P22[4] = IN1[22]&IN2[0];
  assign P23[3] = IN1[22]&IN2[1];
  assign P24[2] = IN1[22]&IN2[2];
  assign P25[1] = IN1[22]&IN2[3];
  assign P26[0] = IN1[22]&IN2[4];
  assign P23[4] = IN1[23]&IN2[0];
  assign P24[3] = IN1[23]&IN2[1];
  assign P25[2] = IN1[23]&IN2[2];
  assign P26[1] = IN1[23]&IN2[3];
  assign P27[0] = IN1[23]&IN2[4];
  assign P24[4] = IN1[24]&IN2[0];
  assign P25[3] = IN1[24]&IN2[1];
  assign P26[2] = IN1[24]&IN2[2];
  assign P27[1] = IN1[24]&IN2[3];
  assign P28[0] = IN1[24]&IN2[4];
  assign P25[4] = IN1[25]&IN2[0];
  assign P26[3] = IN1[25]&IN2[1];
  assign P27[2] = IN1[25]&IN2[2];
  assign P28[1] = IN1[25]&IN2[3];
  assign P29[0] = IN1[25]&IN2[4];
  assign P26[4] = IN1[26]&IN2[0];
  assign P27[3] = IN1[26]&IN2[1];
  assign P28[2] = IN1[26]&IN2[2];
  assign P29[1] = IN1[26]&IN2[3];
  assign P30[0] = IN1[26]&IN2[4];
  assign P27[4] = IN1[27]&IN2[0];
  assign P28[3] = IN1[27]&IN2[1];
  assign P29[2] = IN1[27]&IN2[2];
  assign P30[1] = IN1[27]&IN2[3];
  assign P31[0] = IN1[27]&IN2[4];
  assign P28[4] = IN1[28]&IN2[0];
  assign P29[3] = IN1[28]&IN2[1];
  assign P30[2] = IN1[28]&IN2[2];
  assign P31[1] = IN1[28]&IN2[3];
  assign P32[0] = IN1[28]&IN2[4];
  assign P29[4] = IN1[29]&IN2[0];
  assign P30[3] = IN1[29]&IN2[1];
  assign P31[2] = IN1[29]&IN2[2];
  assign P32[1] = IN1[29]&IN2[3];
  assign P33[0] = IN1[29]&IN2[4];
  assign P30[4] = IN1[30]&IN2[0];
  assign P31[3] = IN1[30]&IN2[1];
  assign P32[2] = IN1[30]&IN2[2];
  assign P33[1] = IN1[30]&IN2[3];
  assign P34[0] = IN1[30]&IN2[4];
  assign P31[4] = IN1[31]&IN2[0];
  assign P32[3] = IN1[31]&IN2[1];
  assign P33[2] = IN1[31]&IN2[2];
  assign P34[1] = IN1[31]&IN2[3];
  assign P35[0] = IN1[31]&IN2[4];
  assign P32[4] = IN1[32]&IN2[0];
  assign P33[3] = IN1[32]&IN2[1];
  assign P34[2] = IN1[32]&IN2[2];
  assign P35[1] = IN1[32]&IN2[3];
  assign P36[0] = IN1[32]&IN2[4];
  assign P33[4] = IN1[33]&IN2[0];
  assign P34[3] = IN1[33]&IN2[1];
  assign P35[2] = IN1[33]&IN2[2];
  assign P36[1] = IN1[33]&IN2[3];
  assign P37[0] = IN1[33]&IN2[4];
  assign P34[4] = IN1[34]&IN2[0];
  assign P35[3] = IN1[34]&IN2[1];
  assign P36[2] = IN1[34]&IN2[2];
  assign P37[1] = IN1[34]&IN2[3];
  assign P38[0] = IN1[34]&IN2[4];
  assign P35[4] = IN1[35]&IN2[0];
  assign P36[3] = IN1[35]&IN2[1];
  assign P37[2] = IN1[35]&IN2[2];
  assign P38[1] = IN1[35]&IN2[3];
  assign P39[0] = IN1[35]&IN2[4];
  assign P36[4] = IN1[36]&IN2[0];
  assign P37[3] = IN1[36]&IN2[1];
  assign P38[2] = IN1[36]&IN2[2];
  assign P39[1] = IN1[36]&IN2[3];
  assign P40[0] = IN1[36]&IN2[4];
  assign P37[4] = IN1[37]&IN2[0];
  assign P38[3] = IN1[37]&IN2[1];
  assign P39[2] = IN1[37]&IN2[2];
  assign P40[1] = IN1[37]&IN2[3];
  assign P41[0] = IN1[37]&IN2[4];
  assign P38[4] = IN1[38]&IN2[0];
  assign P39[3] = IN1[38]&IN2[1];
  assign P40[2] = IN1[38]&IN2[2];
  assign P41[1] = IN1[38]&IN2[3];
  assign P42[0] = IN1[38]&IN2[4];
  assign P39[4] = IN1[39]&IN2[0];
  assign P40[3] = IN1[39]&IN2[1];
  assign P41[2] = IN1[39]&IN2[2];
  assign P42[1] = IN1[39]&IN2[3];
  assign P43[0] = IN1[39]&IN2[4];
  assign P40[4] = IN1[40]&IN2[0];
  assign P41[3] = IN1[40]&IN2[1];
  assign P42[2] = IN1[40]&IN2[2];
  assign P43[1] = IN1[40]&IN2[3];
  assign P44[0] = IN1[40]&IN2[4];
  assign P41[4] = IN1[41]&IN2[0];
  assign P42[3] = IN1[41]&IN2[1];
  assign P43[2] = IN1[41]&IN2[2];
  assign P44[1] = IN1[41]&IN2[3];
  assign P45[0] = IN1[41]&IN2[4];
  assign P42[4] = IN1[42]&IN2[0];
  assign P43[3] = IN1[42]&IN2[1];
  assign P44[2] = IN1[42]&IN2[2];
  assign P45[1] = IN1[42]&IN2[3];
  assign P46[0] = IN1[42]&IN2[4];
  assign P43[4] = IN1[43]&IN2[0];
  assign P44[3] = IN1[43]&IN2[1];
  assign P45[2] = IN1[43]&IN2[2];
  assign P46[1] = IN1[43]&IN2[3];
  assign P47[0] = IN1[43]&IN2[4];
  assign P44[4] = IN1[44]&IN2[0];
  assign P45[3] = IN1[44]&IN2[1];
  assign P46[2] = IN1[44]&IN2[2];
  assign P47[1] = IN1[44]&IN2[3];
  assign P48[0] = IN1[44]&IN2[4];
  assign P45[4] = IN1[45]&IN2[0];
  assign P46[3] = IN1[45]&IN2[1];
  assign P47[2] = IN1[45]&IN2[2];
  assign P48[1] = IN1[45]&IN2[3];
  assign P49[0] = IN1[45]&IN2[4];
  assign P46[4] = IN1[46]&IN2[0];
  assign P47[3] = IN1[46]&IN2[1];
  assign P48[2] = IN1[46]&IN2[2];
  assign P49[1] = IN1[46]&IN2[3];
  assign P50[0] = IN1[46]&IN2[4];
  assign P47[4] = IN1[47]&IN2[0];
  assign P48[3] = IN1[47]&IN2[1];
  assign P49[2] = IN1[47]&IN2[2];
  assign P50[1] = IN1[47]&IN2[3];
  assign P51[0] = IN1[47]&IN2[4];
  assign P48[4] = IN1[48]&IN2[0];
  assign P49[3] = IN1[48]&IN2[1];
  assign P50[2] = IN1[48]&IN2[2];
  assign P51[1] = IN1[48]&IN2[3];
  assign P52[0] = IN1[48]&IN2[4];
  assign P49[4] = IN1[49]&IN2[0];
  assign P50[3] = IN1[49]&IN2[1];
  assign P51[2] = IN1[49]&IN2[2];
  assign P52[1] = IN1[49]&IN2[3];
  assign P53[0] = IN1[49]&IN2[4];
  assign P50[4] = IN1[50]&IN2[0];
  assign P51[3] = IN1[50]&IN2[1];
  assign P52[2] = IN1[50]&IN2[2];
  assign P53[1] = IN1[50]&IN2[3];
  assign P54[0] = IN1[50]&IN2[4];
  assign P51[4] = IN1[51]&IN2[0];
  assign P52[3] = IN1[51]&IN2[1];
  assign P53[2] = IN1[51]&IN2[2];
  assign P54[1] = IN1[51]&IN2[3];
  assign P55[0] = IN1[51]&IN2[4];
  assign P52[4] = IN1[52]&IN2[0];
  assign P53[3] = IN1[52]&IN2[1];
  assign P54[2] = IN1[52]&IN2[2];
  assign P55[1] = IN1[52]&IN2[3];
  assign P56[0] = IN1[52]&IN2[4];
  assign P53[4] = IN1[53]&IN2[0];
  assign P54[3] = IN1[53]&IN2[1];
  assign P55[2] = IN1[53]&IN2[2];
  assign P56[1] = IN1[53]&IN2[3];
  assign P57[0] = IN1[53]&IN2[4];
  assign P54[4] = IN1[54]&IN2[0];
  assign P55[3] = IN1[54]&IN2[1];
  assign P56[2] = IN1[54]&IN2[2];
  assign P57[1] = IN1[54]&IN2[3];
  assign P58[0] = IN1[54]&IN2[4];
  assign P55[4] = IN1[55]&IN2[0];
  assign P56[3] = IN1[55]&IN2[1];
  assign P57[2] = IN1[55]&IN2[2];
  assign P58[1] = IN1[55]&IN2[3];
  assign P59[0] = IN1[55]&IN2[4];
  assign P56[4] = IN1[56]&IN2[0];
  assign P57[3] = IN1[56]&IN2[1];
  assign P58[2] = IN1[56]&IN2[2];
  assign P59[1] = IN1[56]&IN2[3];
  assign P60[0] = IN1[56]&IN2[4];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [4:0] IN5;
  input [4:0] IN6;
  input [4:0] IN7;
  input [4:0] IN8;
  input [4:0] IN9;
  input [4:0] IN10;
  input [4:0] IN11;
  input [4:0] IN12;
  input [4:0] IN13;
  input [4:0] IN14;
  input [4:0] IN15;
  input [4:0] IN16;
  input [4:0] IN17;
  input [4:0] IN18;
  input [4:0] IN19;
  input [4:0] IN20;
  input [4:0] IN21;
  input [4:0] IN22;
  input [4:0] IN23;
  input [4:0] IN24;
  input [4:0] IN25;
  input [4:0] IN26;
  input [4:0] IN27;
  input [4:0] IN28;
  input [4:0] IN29;
  input [4:0] IN30;
  input [4:0] IN31;
  input [4:0] IN32;
  input [4:0] IN33;
  input [4:0] IN34;
  input [4:0] IN35;
  input [4:0] IN36;
  input [4:0] IN37;
  input [4:0] IN38;
  input [4:0] IN39;
  input [4:0] IN40;
  input [4:0] IN41;
  input [4:0] IN42;
  input [4:0] IN43;
  input [4:0] IN44;
  input [4:0] IN45;
  input [4:0] IN46;
  input [4:0] IN47;
  input [4:0] IN48;
  input [4:0] IN49;
  input [4:0] IN50;
  input [4:0] IN51;
  input [4:0] IN52;
  input [4:0] IN53;
  input [4:0] IN54;
  input [4:0] IN55;
  input [4:0] IN56;
  input [3:0] IN57;
  input [2:0] IN58;
  input [1:0] IN59;
  input [0:0] IN60;
  output [60:0] Out1;
  output [3:0] Out2;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w622;
  wire w624;
  wire w626;
  wire w628;
  wire w630;
  wire w632;
  wire w634;
  wire w636;
  wire w638;
  wire w640;
  wire w642;
  wire w644;
  wire w646;
  wire w648;
  wire w650;
  wire w652;
  wire w654;
  wire w656;
  wire w658;
  wire w660;
  wire w662;
  wire w664;
  wire w666;
  wire w668;
  wire w670;
  wire w672;
  wire w674;
  wire w676;
  wire w678;
  wire w680;
  wire w682;
  wire w684;
  wire w686;
  wire w688;
  wire w690;
  wire w692;
  wire w694;
  wire w696;
  wire w698;
  wire w700;
  wire w702;
  wire w704;
  wire w706;
  wire w708;
  wire w710;
  wire w712;
  wire w714;
  wire w716;
  wire w718;
  wire w720;
  wire w722;
  wire w724;
  wire w726;
  wire w728;
  wire w730;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w286);
  FullAdder U1 (w286, IN2[0], IN2[1], w287, w288);
  FullAdder U2 (w288, IN3[0], IN3[1], w289, w290);
  FullAdder U3 (w290, IN4[0], IN4[1], w291, w292);
  FullAdder U4 (w292, IN5[0], IN5[1], w293, w294);
  FullAdder U5 (w294, IN6[0], IN6[1], w295, w296);
  FullAdder U6 (w296, IN7[0], IN7[1], w297, w298);
  FullAdder U7 (w298, IN8[0], IN8[1], w299, w300);
  FullAdder U8 (w300, IN9[0], IN9[1], w301, w302);
  FullAdder U9 (w302, IN10[0], IN10[1], w303, w304);
  FullAdder U10 (w304, IN11[0], IN11[1], w305, w306);
  FullAdder U11 (w306, IN12[0], IN12[1], w307, w308);
  FullAdder U12 (w308, IN13[0], IN13[1], w309, w310);
  FullAdder U13 (w310, IN14[0], IN14[1], w311, w312);
  FullAdder U14 (w312, IN15[0], IN15[1], w313, w314);
  FullAdder U15 (w314, IN16[0], IN16[1], w315, w316);
  FullAdder U16 (w316, IN17[0], IN17[1], w317, w318);
  FullAdder U17 (w318, IN18[0], IN18[1], w319, w320);
  FullAdder U18 (w320, IN19[0], IN19[1], w321, w322);
  FullAdder U19 (w322, IN20[0], IN20[1], w323, w324);
  FullAdder U20 (w324, IN21[0], IN21[1], w325, w326);
  FullAdder U21 (w326, IN22[0], IN22[1], w327, w328);
  FullAdder U22 (w328, IN23[0], IN23[1], w329, w330);
  FullAdder U23 (w330, IN24[0], IN24[1], w331, w332);
  FullAdder U24 (w332, IN25[0], IN25[1], w333, w334);
  FullAdder U25 (w334, IN26[0], IN26[1], w335, w336);
  FullAdder U26 (w336, IN27[0], IN27[1], w337, w338);
  FullAdder U27 (w338, IN28[0], IN28[1], w339, w340);
  FullAdder U28 (w340, IN29[0], IN29[1], w341, w342);
  FullAdder U29 (w342, IN30[0], IN30[1], w343, w344);
  FullAdder U30 (w344, IN31[0], IN31[1], w345, w346);
  FullAdder U31 (w346, IN32[0], IN32[1], w347, w348);
  FullAdder U32 (w348, IN33[0], IN33[1], w349, w350);
  FullAdder U33 (w350, IN34[0], IN34[1], w351, w352);
  FullAdder U34 (w352, IN35[0], IN35[1], w353, w354);
  FullAdder U35 (w354, IN36[0], IN36[1], w355, w356);
  FullAdder U36 (w356, IN37[0], IN37[1], w357, w358);
  FullAdder U37 (w358, IN38[0], IN38[1], w359, w360);
  FullAdder U38 (w360, IN39[0], IN39[1], w361, w362);
  FullAdder U39 (w362, IN40[0], IN40[1], w363, w364);
  FullAdder U40 (w364, IN41[0], IN41[1], w365, w366);
  FullAdder U41 (w366, IN42[0], IN42[1], w367, w368);
  FullAdder U42 (w368, IN43[0], IN43[1], w369, w370);
  FullAdder U43 (w370, IN44[0], IN44[1], w371, w372);
  FullAdder U44 (w372, IN45[0], IN45[1], w373, w374);
  FullAdder U45 (w374, IN46[0], IN46[1], w375, w376);
  FullAdder U46 (w376, IN47[0], IN47[1], w377, w378);
  FullAdder U47 (w378, IN48[0], IN48[1], w379, w380);
  FullAdder U48 (w380, IN49[0], IN49[1], w381, w382);
  FullAdder U49 (w382, IN50[0], IN50[1], w383, w384);
  FullAdder U50 (w384, IN51[0], IN51[1], w385, w386);
  FullAdder U51 (w386, IN52[0], IN52[1], w387, w388);
  FullAdder U52 (w388, IN53[0], IN53[1], w389, w390);
  FullAdder U53 (w390, IN54[0], IN54[1], w391, w392);
  FullAdder U54 (w392, IN55[0], IN55[1], w393, w394);
  FullAdder U55 (w394, IN56[0], IN56[1], w395, w396);
  HalfAdder U56 (w287, IN2[2], Out1[2], w398);
  FullAdder U57 (w398, w289, IN3[2], w399, w400);
  FullAdder U58 (w400, w291, IN4[2], w401, w402);
  FullAdder U59 (w402, w293, IN5[2], w403, w404);
  FullAdder U60 (w404, w295, IN6[2], w405, w406);
  FullAdder U61 (w406, w297, IN7[2], w407, w408);
  FullAdder U62 (w408, w299, IN8[2], w409, w410);
  FullAdder U63 (w410, w301, IN9[2], w411, w412);
  FullAdder U64 (w412, w303, IN10[2], w413, w414);
  FullAdder U65 (w414, w305, IN11[2], w415, w416);
  FullAdder U66 (w416, w307, IN12[2], w417, w418);
  FullAdder U67 (w418, w309, IN13[2], w419, w420);
  FullAdder U68 (w420, w311, IN14[2], w421, w422);
  FullAdder U69 (w422, w313, IN15[2], w423, w424);
  FullAdder U70 (w424, w315, IN16[2], w425, w426);
  FullAdder U71 (w426, w317, IN17[2], w427, w428);
  FullAdder U72 (w428, w319, IN18[2], w429, w430);
  FullAdder U73 (w430, w321, IN19[2], w431, w432);
  FullAdder U74 (w432, w323, IN20[2], w433, w434);
  FullAdder U75 (w434, w325, IN21[2], w435, w436);
  FullAdder U76 (w436, w327, IN22[2], w437, w438);
  FullAdder U77 (w438, w329, IN23[2], w439, w440);
  FullAdder U78 (w440, w331, IN24[2], w441, w442);
  FullAdder U79 (w442, w333, IN25[2], w443, w444);
  FullAdder U80 (w444, w335, IN26[2], w445, w446);
  FullAdder U81 (w446, w337, IN27[2], w447, w448);
  FullAdder U82 (w448, w339, IN28[2], w449, w450);
  FullAdder U83 (w450, w341, IN29[2], w451, w452);
  FullAdder U84 (w452, w343, IN30[2], w453, w454);
  FullAdder U85 (w454, w345, IN31[2], w455, w456);
  FullAdder U86 (w456, w347, IN32[2], w457, w458);
  FullAdder U87 (w458, w349, IN33[2], w459, w460);
  FullAdder U88 (w460, w351, IN34[2], w461, w462);
  FullAdder U89 (w462, w353, IN35[2], w463, w464);
  FullAdder U90 (w464, w355, IN36[2], w465, w466);
  FullAdder U91 (w466, w357, IN37[2], w467, w468);
  FullAdder U92 (w468, w359, IN38[2], w469, w470);
  FullAdder U93 (w470, w361, IN39[2], w471, w472);
  FullAdder U94 (w472, w363, IN40[2], w473, w474);
  FullAdder U95 (w474, w365, IN41[2], w475, w476);
  FullAdder U96 (w476, w367, IN42[2], w477, w478);
  FullAdder U97 (w478, w369, IN43[2], w479, w480);
  FullAdder U98 (w480, w371, IN44[2], w481, w482);
  FullAdder U99 (w482, w373, IN45[2], w483, w484);
  FullAdder U100 (w484, w375, IN46[2], w485, w486);
  FullAdder U101 (w486, w377, IN47[2], w487, w488);
  FullAdder U102 (w488, w379, IN48[2], w489, w490);
  FullAdder U103 (w490, w381, IN49[2], w491, w492);
  FullAdder U104 (w492, w383, IN50[2], w493, w494);
  FullAdder U105 (w494, w385, IN51[2], w495, w496);
  FullAdder U106 (w496, w387, IN52[2], w497, w498);
  FullAdder U107 (w498, w389, IN53[2], w499, w500);
  FullAdder U108 (w500, w391, IN54[2], w501, w502);
  FullAdder U109 (w502, w393, IN55[2], w503, w504);
  FullAdder U110 (w504, w395, IN56[2], w505, w506);
  FullAdder U111 (w506, w396, IN57[0], w507, w508);
  HalfAdder U112 (w399, IN3[3], Out1[3], w510);
  FullAdder U113 (w510, w401, IN4[3], w511, w512);
  FullAdder U114 (w512, w403, IN5[3], w513, w514);
  FullAdder U115 (w514, w405, IN6[3], w515, w516);
  FullAdder U116 (w516, w407, IN7[3], w517, w518);
  FullAdder U117 (w518, w409, IN8[3], w519, w520);
  FullAdder U118 (w520, w411, IN9[3], w521, w522);
  FullAdder U119 (w522, w413, IN10[3], w523, w524);
  FullAdder U120 (w524, w415, IN11[3], w525, w526);
  FullAdder U121 (w526, w417, IN12[3], w527, w528);
  FullAdder U122 (w528, w419, IN13[3], w529, w530);
  FullAdder U123 (w530, w421, IN14[3], w531, w532);
  FullAdder U124 (w532, w423, IN15[3], w533, w534);
  FullAdder U125 (w534, w425, IN16[3], w535, w536);
  FullAdder U126 (w536, w427, IN17[3], w537, w538);
  FullAdder U127 (w538, w429, IN18[3], w539, w540);
  FullAdder U128 (w540, w431, IN19[3], w541, w542);
  FullAdder U129 (w542, w433, IN20[3], w543, w544);
  FullAdder U130 (w544, w435, IN21[3], w545, w546);
  FullAdder U131 (w546, w437, IN22[3], w547, w548);
  FullAdder U132 (w548, w439, IN23[3], w549, w550);
  FullAdder U133 (w550, w441, IN24[3], w551, w552);
  FullAdder U134 (w552, w443, IN25[3], w553, w554);
  FullAdder U135 (w554, w445, IN26[3], w555, w556);
  FullAdder U136 (w556, w447, IN27[3], w557, w558);
  FullAdder U137 (w558, w449, IN28[3], w559, w560);
  FullAdder U138 (w560, w451, IN29[3], w561, w562);
  FullAdder U139 (w562, w453, IN30[3], w563, w564);
  FullAdder U140 (w564, w455, IN31[3], w565, w566);
  FullAdder U141 (w566, w457, IN32[3], w567, w568);
  FullAdder U142 (w568, w459, IN33[3], w569, w570);
  FullAdder U143 (w570, w461, IN34[3], w571, w572);
  FullAdder U144 (w572, w463, IN35[3], w573, w574);
  FullAdder U145 (w574, w465, IN36[3], w575, w576);
  FullAdder U146 (w576, w467, IN37[3], w577, w578);
  FullAdder U147 (w578, w469, IN38[3], w579, w580);
  FullAdder U148 (w580, w471, IN39[3], w581, w582);
  FullAdder U149 (w582, w473, IN40[3], w583, w584);
  FullAdder U150 (w584, w475, IN41[3], w585, w586);
  FullAdder U151 (w586, w477, IN42[3], w587, w588);
  FullAdder U152 (w588, w479, IN43[3], w589, w590);
  FullAdder U153 (w590, w481, IN44[3], w591, w592);
  FullAdder U154 (w592, w483, IN45[3], w593, w594);
  FullAdder U155 (w594, w485, IN46[3], w595, w596);
  FullAdder U156 (w596, w487, IN47[3], w597, w598);
  FullAdder U157 (w598, w489, IN48[3], w599, w600);
  FullAdder U158 (w600, w491, IN49[3], w601, w602);
  FullAdder U159 (w602, w493, IN50[3], w603, w604);
  FullAdder U160 (w604, w495, IN51[3], w605, w606);
  FullAdder U161 (w606, w497, IN52[3], w607, w608);
  FullAdder U162 (w608, w499, IN53[3], w609, w610);
  FullAdder U163 (w610, w501, IN54[3], w611, w612);
  FullAdder U164 (w612, w503, IN55[3], w613, w614);
  FullAdder U165 (w614, w505, IN56[3], w615, w616);
  FullAdder U166 (w616, w507, IN57[1], w617, w618);
  FullAdder U167 (w618, w508, IN58[0], w619, w620);
  HalfAdder U168 (w511, IN4[4], Out1[4], w622);
  FullAdder U169 (w622, w513, IN5[4], Out1[5], w624);
  FullAdder U170 (w624, w515, IN6[4], Out1[6], w626);
  FullAdder U171 (w626, w517, IN7[4], Out1[7], w628);
  FullAdder U172 (w628, w519, IN8[4], Out1[8], w630);
  FullAdder U173 (w630, w521, IN9[4], Out1[9], w632);
  FullAdder U174 (w632, w523, IN10[4], Out1[10], w634);
  FullAdder U175 (w634, w525, IN11[4], Out1[11], w636);
  FullAdder U176 (w636, w527, IN12[4], Out1[12], w638);
  FullAdder U177 (w638, w529, IN13[4], Out1[13], w640);
  FullAdder U178 (w640, w531, IN14[4], Out1[14], w642);
  FullAdder U179 (w642, w533, IN15[4], Out1[15], w644);
  FullAdder U180 (w644, w535, IN16[4], Out1[16], w646);
  FullAdder U181 (w646, w537, IN17[4], Out1[17], w648);
  FullAdder U182 (w648, w539, IN18[4], Out1[18], w650);
  FullAdder U183 (w650, w541, IN19[4], Out1[19], w652);
  FullAdder U184 (w652, w543, IN20[4], Out1[20], w654);
  FullAdder U185 (w654, w545, IN21[4], Out1[21], w656);
  FullAdder U186 (w656, w547, IN22[4], Out1[22], w658);
  FullAdder U187 (w658, w549, IN23[4], Out1[23], w660);
  FullAdder U188 (w660, w551, IN24[4], Out1[24], w662);
  FullAdder U189 (w662, w553, IN25[4], Out1[25], w664);
  FullAdder U190 (w664, w555, IN26[4], Out1[26], w666);
  FullAdder U191 (w666, w557, IN27[4], Out1[27], w668);
  FullAdder U192 (w668, w559, IN28[4], Out1[28], w670);
  FullAdder U193 (w670, w561, IN29[4], Out1[29], w672);
  FullAdder U194 (w672, w563, IN30[4], Out1[30], w674);
  FullAdder U195 (w674, w565, IN31[4], Out1[31], w676);
  FullAdder U196 (w676, w567, IN32[4], Out1[32], w678);
  FullAdder U197 (w678, w569, IN33[4], Out1[33], w680);
  FullAdder U198 (w680, w571, IN34[4], Out1[34], w682);
  FullAdder U199 (w682, w573, IN35[4], Out1[35], w684);
  FullAdder U200 (w684, w575, IN36[4], Out1[36], w686);
  FullAdder U201 (w686, w577, IN37[4], Out1[37], w688);
  FullAdder U202 (w688, w579, IN38[4], Out1[38], w690);
  FullAdder U203 (w690, w581, IN39[4], Out1[39], w692);
  FullAdder U204 (w692, w583, IN40[4], Out1[40], w694);
  FullAdder U205 (w694, w585, IN41[4], Out1[41], w696);
  FullAdder U206 (w696, w587, IN42[4], Out1[42], w698);
  FullAdder U207 (w698, w589, IN43[4], Out1[43], w700);
  FullAdder U208 (w700, w591, IN44[4], Out1[44], w702);
  FullAdder U209 (w702, w593, IN45[4], Out1[45], w704);
  FullAdder U210 (w704, w595, IN46[4], Out1[46], w706);
  FullAdder U211 (w706, w597, IN47[4], Out1[47], w708);
  FullAdder U212 (w708, w599, IN48[4], Out1[48], w710);
  FullAdder U213 (w710, w601, IN49[4], Out1[49], w712);
  FullAdder U214 (w712, w603, IN50[4], Out1[50], w714);
  FullAdder U215 (w714, w605, IN51[4], Out1[51], w716);
  FullAdder U216 (w716, w607, IN52[4], Out1[52], w718);
  FullAdder U217 (w718, w609, IN53[4], Out1[53], w720);
  FullAdder U218 (w720, w611, IN54[4], Out1[54], w722);
  FullAdder U219 (w722, w613, IN55[4], Out1[55], w724);
  FullAdder U220 (w724, w615, IN56[4], Out1[56], w726);
  FullAdder U221 (w726, w617, IN57[2], Out1[57], w728);
  FullAdder U222 (w728, w619, IN58[1], Out1[58], w730);
  FullAdder U223 (w730, w620, IN59[0], Out1[59], Out1[60]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN57[3];
  assign Out2[1] = IN58[2];
  assign Out2[2] = IN59[1];
  assign Out2[3] = IN60[0];

endmodule
module RC_4_4(IN1, IN2, Out);
  input [3:0] IN1;
  input [3:0] IN2;
  output [4:0] Out;
  wire w9;
  wire w11;
  wire w13;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w9);
  FullAdder U1 (IN1[1], IN2[1], w9, Out[1], w11);
  FullAdder U2 (IN1[2], IN2[2], w11, Out[2], w13);
  FullAdder U3 (IN1[3], IN2[3], w13, Out[3], Out[4]);

endmodule
module NR_57_5(IN1, IN2, Out);
  input [56:0] IN1;
  input [4:0] IN2;
  output [61:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [4:0] P5;
  wire [4:0] P6;
  wire [4:0] P7;
  wire [4:0] P8;
  wire [4:0] P9;
  wire [4:0] P10;
  wire [4:0] P11;
  wire [4:0] P12;
  wire [4:0] P13;
  wire [4:0] P14;
  wire [4:0] P15;
  wire [4:0] P16;
  wire [4:0] P17;
  wire [4:0] P18;
  wire [4:0] P19;
  wire [4:0] P20;
  wire [4:0] P21;
  wire [4:0] P22;
  wire [4:0] P23;
  wire [4:0] P24;
  wire [4:0] P25;
  wire [4:0] P26;
  wire [4:0] P27;
  wire [4:0] P28;
  wire [4:0] P29;
  wire [4:0] P30;
  wire [4:0] P31;
  wire [4:0] P32;
  wire [4:0] P33;
  wire [4:0] P34;
  wire [4:0] P35;
  wire [4:0] P36;
  wire [4:0] P37;
  wire [4:0] P38;
  wire [4:0] P39;
  wire [4:0] P40;
  wire [4:0] P41;
  wire [4:0] P42;
  wire [4:0] P43;
  wire [4:0] P44;
  wire [4:0] P45;
  wire [4:0] P46;
  wire [4:0] P47;
  wire [4:0] P48;
  wire [4:0] P49;
  wire [4:0] P50;
  wire [4:0] P51;
  wire [4:0] P52;
  wire [4:0] P53;
  wire [4:0] P54;
  wire [4:0] P55;
  wire [4:0] P56;
  wire [3:0] P57;
  wire [2:0] P58;
  wire [1:0] P59;
  wire [0:0] P60;
  wire [60:0] R1;
  wire [3:0] R2;
  wire [61:0] aOut;
  U_SP_57_5 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, R1, R2);
  RC_4_4 S2 (R1[60:57], R2, aOut[61:57]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign Out = aOut[61:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
