//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 17
  second input length: 38
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_17_38(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53);
  input [16:0] IN1;
  input [37:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [16:0] P17;
  output [16:0] P18;
  output [16:0] P19;
  output [16:0] P20;
  output [16:0] P21;
  output [16:0] P22;
  output [16:0] P23;
  output [16:0] P24;
  output [16:0] P25;
  output [16:0] P26;
  output [16:0] P27;
  output [16:0] P28;
  output [16:0] P29;
  output [16:0] P30;
  output [16:0] P31;
  output [16:0] P32;
  output [16:0] P33;
  output [16:0] P34;
  output [16:0] P35;
  output [16:0] P36;
  output [16:0] P37;
  output [15:0] P38;
  output [14:0] P39;
  output [13:0] P40;
  output [12:0] P41;
  output [11:0] P42;
  output [10:0] P43;
  output [9:0] P44;
  output [8:0] P45;
  output [7:0] P46;
  output [6:0] P47;
  output [5:0] P48;
  output [4:0] P49;
  output [3:0] P50;
  output [2:0] P51;
  output [1:0] P52;
  output [0:0] P53;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[0] = IN1[1]&IN2[37];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[1] = IN1[2]&IN2[36];
  assign P39[0] = IN1[2]&IN2[37];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[2] = IN1[3]&IN2[35];
  assign P39[1] = IN1[3]&IN2[36];
  assign P40[0] = IN1[3]&IN2[37];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[3] = IN1[4]&IN2[34];
  assign P39[2] = IN1[4]&IN2[35];
  assign P40[1] = IN1[4]&IN2[36];
  assign P41[0] = IN1[4]&IN2[37];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[4] = IN1[5]&IN2[33];
  assign P39[3] = IN1[5]&IN2[34];
  assign P40[2] = IN1[5]&IN2[35];
  assign P41[1] = IN1[5]&IN2[36];
  assign P42[0] = IN1[5]&IN2[37];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[5] = IN1[6]&IN2[32];
  assign P39[4] = IN1[6]&IN2[33];
  assign P40[3] = IN1[6]&IN2[34];
  assign P41[2] = IN1[6]&IN2[35];
  assign P42[1] = IN1[6]&IN2[36];
  assign P43[0] = IN1[6]&IN2[37];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[6] = IN1[7]&IN2[31];
  assign P39[5] = IN1[7]&IN2[32];
  assign P40[4] = IN1[7]&IN2[33];
  assign P41[3] = IN1[7]&IN2[34];
  assign P42[2] = IN1[7]&IN2[35];
  assign P43[1] = IN1[7]&IN2[36];
  assign P44[0] = IN1[7]&IN2[37];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[7] = IN1[8]&IN2[30];
  assign P39[6] = IN1[8]&IN2[31];
  assign P40[5] = IN1[8]&IN2[32];
  assign P41[4] = IN1[8]&IN2[33];
  assign P42[3] = IN1[8]&IN2[34];
  assign P43[2] = IN1[8]&IN2[35];
  assign P44[1] = IN1[8]&IN2[36];
  assign P45[0] = IN1[8]&IN2[37];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[8] = IN1[9]&IN2[29];
  assign P39[7] = IN1[9]&IN2[30];
  assign P40[6] = IN1[9]&IN2[31];
  assign P41[5] = IN1[9]&IN2[32];
  assign P42[4] = IN1[9]&IN2[33];
  assign P43[3] = IN1[9]&IN2[34];
  assign P44[2] = IN1[9]&IN2[35];
  assign P45[1] = IN1[9]&IN2[36];
  assign P46[0] = IN1[9]&IN2[37];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[9] = IN1[10]&IN2[28];
  assign P39[8] = IN1[10]&IN2[29];
  assign P40[7] = IN1[10]&IN2[30];
  assign P41[6] = IN1[10]&IN2[31];
  assign P42[5] = IN1[10]&IN2[32];
  assign P43[4] = IN1[10]&IN2[33];
  assign P44[3] = IN1[10]&IN2[34];
  assign P45[2] = IN1[10]&IN2[35];
  assign P46[1] = IN1[10]&IN2[36];
  assign P47[0] = IN1[10]&IN2[37];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[10] = IN1[11]&IN2[27];
  assign P39[9] = IN1[11]&IN2[28];
  assign P40[8] = IN1[11]&IN2[29];
  assign P41[7] = IN1[11]&IN2[30];
  assign P42[6] = IN1[11]&IN2[31];
  assign P43[5] = IN1[11]&IN2[32];
  assign P44[4] = IN1[11]&IN2[33];
  assign P45[3] = IN1[11]&IN2[34];
  assign P46[2] = IN1[11]&IN2[35];
  assign P47[1] = IN1[11]&IN2[36];
  assign P48[0] = IN1[11]&IN2[37];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[11] = IN1[12]&IN2[26];
  assign P39[10] = IN1[12]&IN2[27];
  assign P40[9] = IN1[12]&IN2[28];
  assign P41[8] = IN1[12]&IN2[29];
  assign P42[7] = IN1[12]&IN2[30];
  assign P43[6] = IN1[12]&IN2[31];
  assign P44[5] = IN1[12]&IN2[32];
  assign P45[4] = IN1[12]&IN2[33];
  assign P46[3] = IN1[12]&IN2[34];
  assign P47[2] = IN1[12]&IN2[35];
  assign P48[1] = IN1[12]&IN2[36];
  assign P49[0] = IN1[12]&IN2[37];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[12] = IN1[13]&IN2[25];
  assign P39[11] = IN1[13]&IN2[26];
  assign P40[10] = IN1[13]&IN2[27];
  assign P41[9] = IN1[13]&IN2[28];
  assign P42[8] = IN1[13]&IN2[29];
  assign P43[7] = IN1[13]&IN2[30];
  assign P44[6] = IN1[13]&IN2[31];
  assign P45[5] = IN1[13]&IN2[32];
  assign P46[4] = IN1[13]&IN2[33];
  assign P47[3] = IN1[13]&IN2[34];
  assign P48[2] = IN1[13]&IN2[35];
  assign P49[1] = IN1[13]&IN2[36];
  assign P50[0] = IN1[13]&IN2[37];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[13] = IN1[14]&IN2[24];
  assign P39[12] = IN1[14]&IN2[25];
  assign P40[11] = IN1[14]&IN2[26];
  assign P41[10] = IN1[14]&IN2[27];
  assign P42[9] = IN1[14]&IN2[28];
  assign P43[8] = IN1[14]&IN2[29];
  assign P44[7] = IN1[14]&IN2[30];
  assign P45[6] = IN1[14]&IN2[31];
  assign P46[5] = IN1[14]&IN2[32];
  assign P47[4] = IN1[14]&IN2[33];
  assign P48[3] = IN1[14]&IN2[34];
  assign P49[2] = IN1[14]&IN2[35];
  assign P50[1] = IN1[14]&IN2[36];
  assign P51[0] = IN1[14]&IN2[37];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[14] = IN1[15]&IN2[23];
  assign P39[13] = IN1[15]&IN2[24];
  assign P40[12] = IN1[15]&IN2[25];
  assign P41[11] = IN1[15]&IN2[26];
  assign P42[10] = IN1[15]&IN2[27];
  assign P43[9] = IN1[15]&IN2[28];
  assign P44[8] = IN1[15]&IN2[29];
  assign P45[7] = IN1[15]&IN2[30];
  assign P46[6] = IN1[15]&IN2[31];
  assign P47[5] = IN1[15]&IN2[32];
  assign P48[4] = IN1[15]&IN2[33];
  assign P49[3] = IN1[15]&IN2[34];
  assign P50[2] = IN1[15]&IN2[35];
  assign P51[1] = IN1[15]&IN2[36];
  assign P52[0] = IN1[15]&IN2[37];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[15] = IN1[16]&IN2[22];
  assign P39[14] = IN1[16]&IN2[23];
  assign P40[13] = IN1[16]&IN2[24];
  assign P41[12] = IN1[16]&IN2[25];
  assign P42[11] = IN1[16]&IN2[26];
  assign P43[10] = IN1[16]&IN2[27];
  assign P44[9] = IN1[16]&IN2[28];
  assign P45[8] = IN1[16]&IN2[29];
  assign P46[7] = IN1[16]&IN2[30];
  assign P47[6] = IN1[16]&IN2[31];
  assign P48[5] = IN1[16]&IN2[32];
  assign P49[4] = IN1[16]&IN2[33];
  assign P50[3] = IN1[16]&IN2[34];
  assign P51[2] = IN1[16]&IN2[35];
  assign P52[1] = IN1[16]&IN2[36];
  assign P53[0] = IN1[16]&IN2[37];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [16:0] IN17;
  input [16:0] IN18;
  input [16:0] IN19;
  input [16:0] IN20;
  input [16:0] IN21;
  input [16:0] IN22;
  input [16:0] IN23;
  input [16:0] IN24;
  input [16:0] IN25;
  input [16:0] IN26;
  input [16:0] IN27;
  input [16:0] IN28;
  input [16:0] IN29;
  input [16:0] IN30;
  input [16:0] IN31;
  input [16:0] IN32;
  input [16:0] IN33;
  input [16:0] IN34;
  input [16:0] IN35;
  input [16:0] IN36;
  input [16:0] IN37;
  input [15:0] IN38;
  input [14:0] IN39;
  input [13:0] IN40;
  input [12:0] IN41;
  input [11:0] IN42;
  input [10:0] IN43;
  input [9:0] IN44;
  input [8:0] IN45;
  input [7:0] IN46;
  input [6:0] IN47;
  input [5:0] IN48;
  input [4:0] IN49;
  input [3:0] IN50;
  input [2:0] IN51;
  input [1:0] IN52;
  input [0:0] IN53;
  output [53:0] Out1;
  output [36:0] Out2;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1799;
  wire w1801;
  wire w1803;
  wire w1805;
  wire w1807;
  wire w1809;
  wire w1811;
  wire w1813;
  wire w1815;
  wire w1817;
  wire w1819;
  wire w1821;
  wire w1823;
  wire w1825;
  wire w1827;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w647);
  FullAdder U1 (w647, IN2[0], IN2[1], w648, w649);
  FullAdder U2 (w649, IN3[0], IN3[1], w650, w651);
  FullAdder U3 (w651, IN4[0], IN4[1], w652, w653);
  FullAdder U4 (w653, IN5[0], IN5[1], w654, w655);
  FullAdder U5 (w655, IN6[0], IN6[1], w656, w657);
  FullAdder U6 (w657, IN7[0], IN7[1], w658, w659);
  FullAdder U7 (w659, IN8[0], IN8[1], w660, w661);
  FullAdder U8 (w661, IN9[0], IN9[1], w662, w663);
  FullAdder U9 (w663, IN10[0], IN10[1], w664, w665);
  FullAdder U10 (w665, IN11[0], IN11[1], w666, w667);
  FullAdder U11 (w667, IN12[0], IN12[1], w668, w669);
  FullAdder U12 (w669, IN13[0], IN13[1], w670, w671);
  FullAdder U13 (w671, IN14[0], IN14[1], w672, w673);
  FullAdder U14 (w673, IN15[0], IN15[1], w674, w675);
  FullAdder U15 (w675, IN16[0], IN16[1], w676, w677);
  HalfAdder U16 (w648, IN2[2], Out1[2], w679);
  FullAdder U17 (w679, w650, IN3[2], w680, w681);
  FullAdder U18 (w681, w652, IN4[2], w682, w683);
  FullAdder U19 (w683, w654, IN5[2], w684, w685);
  FullAdder U20 (w685, w656, IN6[2], w686, w687);
  FullAdder U21 (w687, w658, IN7[2], w688, w689);
  FullAdder U22 (w689, w660, IN8[2], w690, w691);
  FullAdder U23 (w691, w662, IN9[2], w692, w693);
  FullAdder U24 (w693, w664, IN10[2], w694, w695);
  FullAdder U25 (w695, w666, IN11[2], w696, w697);
  FullAdder U26 (w697, w668, IN12[2], w698, w699);
  FullAdder U27 (w699, w670, IN13[2], w700, w701);
  FullAdder U28 (w701, w672, IN14[2], w702, w703);
  FullAdder U29 (w703, w674, IN15[2], w704, w705);
  FullAdder U30 (w705, w676, IN16[2], w706, w707);
  FullAdder U31 (w707, w677, IN17[0], w708, w709);
  HalfAdder U32 (w680, IN3[3], Out1[3], w711);
  FullAdder U33 (w711, w682, IN4[3], w712, w713);
  FullAdder U34 (w713, w684, IN5[3], w714, w715);
  FullAdder U35 (w715, w686, IN6[3], w716, w717);
  FullAdder U36 (w717, w688, IN7[3], w718, w719);
  FullAdder U37 (w719, w690, IN8[3], w720, w721);
  FullAdder U38 (w721, w692, IN9[3], w722, w723);
  FullAdder U39 (w723, w694, IN10[3], w724, w725);
  FullAdder U40 (w725, w696, IN11[3], w726, w727);
  FullAdder U41 (w727, w698, IN12[3], w728, w729);
  FullAdder U42 (w729, w700, IN13[3], w730, w731);
  FullAdder U43 (w731, w702, IN14[3], w732, w733);
  FullAdder U44 (w733, w704, IN15[3], w734, w735);
  FullAdder U45 (w735, w706, IN16[3], w736, w737);
  FullAdder U46 (w737, w708, IN17[1], w738, w739);
  FullAdder U47 (w739, w709, IN18[0], w740, w741);
  HalfAdder U48 (w712, IN4[4], Out1[4], w743);
  FullAdder U49 (w743, w714, IN5[4], w744, w745);
  FullAdder U50 (w745, w716, IN6[4], w746, w747);
  FullAdder U51 (w747, w718, IN7[4], w748, w749);
  FullAdder U52 (w749, w720, IN8[4], w750, w751);
  FullAdder U53 (w751, w722, IN9[4], w752, w753);
  FullAdder U54 (w753, w724, IN10[4], w754, w755);
  FullAdder U55 (w755, w726, IN11[4], w756, w757);
  FullAdder U56 (w757, w728, IN12[4], w758, w759);
  FullAdder U57 (w759, w730, IN13[4], w760, w761);
  FullAdder U58 (w761, w732, IN14[4], w762, w763);
  FullAdder U59 (w763, w734, IN15[4], w764, w765);
  FullAdder U60 (w765, w736, IN16[4], w766, w767);
  FullAdder U61 (w767, w738, IN17[2], w768, w769);
  FullAdder U62 (w769, w740, IN18[1], w770, w771);
  FullAdder U63 (w771, w741, IN19[0], w772, w773);
  HalfAdder U64 (w744, IN5[5], Out1[5], w775);
  FullAdder U65 (w775, w746, IN6[5], w776, w777);
  FullAdder U66 (w777, w748, IN7[5], w778, w779);
  FullAdder U67 (w779, w750, IN8[5], w780, w781);
  FullAdder U68 (w781, w752, IN9[5], w782, w783);
  FullAdder U69 (w783, w754, IN10[5], w784, w785);
  FullAdder U70 (w785, w756, IN11[5], w786, w787);
  FullAdder U71 (w787, w758, IN12[5], w788, w789);
  FullAdder U72 (w789, w760, IN13[5], w790, w791);
  FullAdder U73 (w791, w762, IN14[5], w792, w793);
  FullAdder U74 (w793, w764, IN15[5], w794, w795);
  FullAdder U75 (w795, w766, IN16[5], w796, w797);
  FullAdder U76 (w797, w768, IN17[3], w798, w799);
  FullAdder U77 (w799, w770, IN18[2], w800, w801);
  FullAdder U78 (w801, w772, IN19[1], w802, w803);
  FullAdder U79 (w803, w773, IN20[0], w804, w805);
  HalfAdder U80 (w776, IN6[6], Out1[6], w807);
  FullAdder U81 (w807, w778, IN7[6], w808, w809);
  FullAdder U82 (w809, w780, IN8[6], w810, w811);
  FullAdder U83 (w811, w782, IN9[6], w812, w813);
  FullAdder U84 (w813, w784, IN10[6], w814, w815);
  FullAdder U85 (w815, w786, IN11[6], w816, w817);
  FullAdder U86 (w817, w788, IN12[6], w818, w819);
  FullAdder U87 (w819, w790, IN13[6], w820, w821);
  FullAdder U88 (w821, w792, IN14[6], w822, w823);
  FullAdder U89 (w823, w794, IN15[6], w824, w825);
  FullAdder U90 (w825, w796, IN16[6], w826, w827);
  FullAdder U91 (w827, w798, IN17[4], w828, w829);
  FullAdder U92 (w829, w800, IN18[3], w830, w831);
  FullAdder U93 (w831, w802, IN19[2], w832, w833);
  FullAdder U94 (w833, w804, IN20[1], w834, w835);
  FullAdder U95 (w835, w805, IN21[0], w836, w837);
  HalfAdder U96 (w808, IN7[7], Out1[7], w839);
  FullAdder U97 (w839, w810, IN8[7], w840, w841);
  FullAdder U98 (w841, w812, IN9[7], w842, w843);
  FullAdder U99 (w843, w814, IN10[7], w844, w845);
  FullAdder U100 (w845, w816, IN11[7], w846, w847);
  FullAdder U101 (w847, w818, IN12[7], w848, w849);
  FullAdder U102 (w849, w820, IN13[7], w850, w851);
  FullAdder U103 (w851, w822, IN14[7], w852, w853);
  FullAdder U104 (w853, w824, IN15[7], w854, w855);
  FullAdder U105 (w855, w826, IN16[7], w856, w857);
  FullAdder U106 (w857, w828, IN17[5], w858, w859);
  FullAdder U107 (w859, w830, IN18[4], w860, w861);
  FullAdder U108 (w861, w832, IN19[3], w862, w863);
  FullAdder U109 (w863, w834, IN20[2], w864, w865);
  FullAdder U110 (w865, w836, IN21[1], w866, w867);
  FullAdder U111 (w867, w837, IN22[0], w868, w869);
  HalfAdder U112 (w840, IN8[8], Out1[8], w871);
  FullAdder U113 (w871, w842, IN9[8], w872, w873);
  FullAdder U114 (w873, w844, IN10[8], w874, w875);
  FullAdder U115 (w875, w846, IN11[8], w876, w877);
  FullAdder U116 (w877, w848, IN12[8], w878, w879);
  FullAdder U117 (w879, w850, IN13[8], w880, w881);
  FullAdder U118 (w881, w852, IN14[8], w882, w883);
  FullAdder U119 (w883, w854, IN15[8], w884, w885);
  FullAdder U120 (w885, w856, IN16[8], w886, w887);
  FullAdder U121 (w887, w858, IN17[6], w888, w889);
  FullAdder U122 (w889, w860, IN18[5], w890, w891);
  FullAdder U123 (w891, w862, IN19[4], w892, w893);
  FullAdder U124 (w893, w864, IN20[3], w894, w895);
  FullAdder U125 (w895, w866, IN21[2], w896, w897);
  FullAdder U126 (w897, w868, IN22[1], w898, w899);
  FullAdder U127 (w899, w869, IN23[0], w900, w901);
  HalfAdder U128 (w872, IN9[9], Out1[9], w903);
  FullAdder U129 (w903, w874, IN10[9], w904, w905);
  FullAdder U130 (w905, w876, IN11[9], w906, w907);
  FullAdder U131 (w907, w878, IN12[9], w908, w909);
  FullAdder U132 (w909, w880, IN13[9], w910, w911);
  FullAdder U133 (w911, w882, IN14[9], w912, w913);
  FullAdder U134 (w913, w884, IN15[9], w914, w915);
  FullAdder U135 (w915, w886, IN16[9], w916, w917);
  FullAdder U136 (w917, w888, IN17[7], w918, w919);
  FullAdder U137 (w919, w890, IN18[6], w920, w921);
  FullAdder U138 (w921, w892, IN19[5], w922, w923);
  FullAdder U139 (w923, w894, IN20[4], w924, w925);
  FullAdder U140 (w925, w896, IN21[3], w926, w927);
  FullAdder U141 (w927, w898, IN22[2], w928, w929);
  FullAdder U142 (w929, w900, IN23[1], w930, w931);
  FullAdder U143 (w931, w901, IN24[0], w932, w933);
  HalfAdder U144 (w904, IN10[10], Out1[10], w935);
  FullAdder U145 (w935, w906, IN11[10], w936, w937);
  FullAdder U146 (w937, w908, IN12[10], w938, w939);
  FullAdder U147 (w939, w910, IN13[10], w940, w941);
  FullAdder U148 (w941, w912, IN14[10], w942, w943);
  FullAdder U149 (w943, w914, IN15[10], w944, w945);
  FullAdder U150 (w945, w916, IN16[10], w946, w947);
  FullAdder U151 (w947, w918, IN17[8], w948, w949);
  FullAdder U152 (w949, w920, IN18[7], w950, w951);
  FullAdder U153 (w951, w922, IN19[6], w952, w953);
  FullAdder U154 (w953, w924, IN20[5], w954, w955);
  FullAdder U155 (w955, w926, IN21[4], w956, w957);
  FullAdder U156 (w957, w928, IN22[3], w958, w959);
  FullAdder U157 (w959, w930, IN23[2], w960, w961);
  FullAdder U158 (w961, w932, IN24[1], w962, w963);
  FullAdder U159 (w963, w933, IN25[0], w964, w965);
  HalfAdder U160 (w936, IN11[11], Out1[11], w967);
  FullAdder U161 (w967, w938, IN12[11], w968, w969);
  FullAdder U162 (w969, w940, IN13[11], w970, w971);
  FullAdder U163 (w971, w942, IN14[11], w972, w973);
  FullAdder U164 (w973, w944, IN15[11], w974, w975);
  FullAdder U165 (w975, w946, IN16[11], w976, w977);
  FullAdder U166 (w977, w948, IN17[9], w978, w979);
  FullAdder U167 (w979, w950, IN18[8], w980, w981);
  FullAdder U168 (w981, w952, IN19[7], w982, w983);
  FullAdder U169 (w983, w954, IN20[6], w984, w985);
  FullAdder U170 (w985, w956, IN21[5], w986, w987);
  FullAdder U171 (w987, w958, IN22[4], w988, w989);
  FullAdder U172 (w989, w960, IN23[3], w990, w991);
  FullAdder U173 (w991, w962, IN24[2], w992, w993);
  FullAdder U174 (w993, w964, IN25[1], w994, w995);
  FullAdder U175 (w995, w965, IN26[0], w996, w997);
  HalfAdder U176 (w968, IN12[12], Out1[12], w999);
  FullAdder U177 (w999, w970, IN13[12], w1000, w1001);
  FullAdder U178 (w1001, w972, IN14[12], w1002, w1003);
  FullAdder U179 (w1003, w974, IN15[12], w1004, w1005);
  FullAdder U180 (w1005, w976, IN16[12], w1006, w1007);
  FullAdder U181 (w1007, w978, IN17[10], w1008, w1009);
  FullAdder U182 (w1009, w980, IN18[9], w1010, w1011);
  FullAdder U183 (w1011, w982, IN19[8], w1012, w1013);
  FullAdder U184 (w1013, w984, IN20[7], w1014, w1015);
  FullAdder U185 (w1015, w986, IN21[6], w1016, w1017);
  FullAdder U186 (w1017, w988, IN22[5], w1018, w1019);
  FullAdder U187 (w1019, w990, IN23[4], w1020, w1021);
  FullAdder U188 (w1021, w992, IN24[3], w1022, w1023);
  FullAdder U189 (w1023, w994, IN25[2], w1024, w1025);
  FullAdder U190 (w1025, w996, IN26[1], w1026, w1027);
  FullAdder U191 (w1027, w997, IN27[0], w1028, w1029);
  HalfAdder U192 (w1000, IN13[13], Out1[13], w1031);
  FullAdder U193 (w1031, w1002, IN14[13], w1032, w1033);
  FullAdder U194 (w1033, w1004, IN15[13], w1034, w1035);
  FullAdder U195 (w1035, w1006, IN16[13], w1036, w1037);
  FullAdder U196 (w1037, w1008, IN17[11], w1038, w1039);
  FullAdder U197 (w1039, w1010, IN18[10], w1040, w1041);
  FullAdder U198 (w1041, w1012, IN19[9], w1042, w1043);
  FullAdder U199 (w1043, w1014, IN20[8], w1044, w1045);
  FullAdder U200 (w1045, w1016, IN21[7], w1046, w1047);
  FullAdder U201 (w1047, w1018, IN22[6], w1048, w1049);
  FullAdder U202 (w1049, w1020, IN23[5], w1050, w1051);
  FullAdder U203 (w1051, w1022, IN24[4], w1052, w1053);
  FullAdder U204 (w1053, w1024, IN25[3], w1054, w1055);
  FullAdder U205 (w1055, w1026, IN26[2], w1056, w1057);
  FullAdder U206 (w1057, w1028, IN27[1], w1058, w1059);
  FullAdder U207 (w1059, w1029, IN28[0], w1060, w1061);
  HalfAdder U208 (w1032, IN14[14], Out1[14], w1063);
  FullAdder U209 (w1063, w1034, IN15[14], w1064, w1065);
  FullAdder U210 (w1065, w1036, IN16[14], w1066, w1067);
  FullAdder U211 (w1067, w1038, IN17[12], w1068, w1069);
  FullAdder U212 (w1069, w1040, IN18[11], w1070, w1071);
  FullAdder U213 (w1071, w1042, IN19[10], w1072, w1073);
  FullAdder U214 (w1073, w1044, IN20[9], w1074, w1075);
  FullAdder U215 (w1075, w1046, IN21[8], w1076, w1077);
  FullAdder U216 (w1077, w1048, IN22[7], w1078, w1079);
  FullAdder U217 (w1079, w1050, IN23[6], w1080, w1081);
  FullAdder U218 (w1081, w1052, IN24[5], w1082, w1083);
  FullAdder U219 (w1083, w1054, IN25[4], w1084, w1085);
  FullAdder U220 (w1085, w1056, IN26[3], w1086, w1087);
  FullAdder U221 (w1087, w1058, IN27[2], w1088, w1089);
  FullAdder U222 (w1089, w1060, IN28[1], w1090, w1091);
  FullAdder U223 (w1091, w1061, IN29[0], w1092, w1093);
  HalfAdder U224 (w1064, IN15[15], Out1[15], w1095);
  FullAdder U225 (w1095, w1066, IN16[15], w1096, w1097);
  FullAdder U226 (w1097, w1068, IN17[13], w1098, w1099);
  FullAdder U227 (w1099, w1070, IN18[12], w1100, w1101);
  FullAdder U228 (w1101, w1072, IN19[11], w1102, w1103);
  FullAdder U229 (w1103, w1074, IN20[10], w1104, w1105);
  FullAdder U230 (w1105, w1076, IN21[9], w1106, w1107);
  FullAdder U231 (w1107, w1078, IN22[8], w1108, w1109);
  FullAdder U232 (w1109, w1080, IN23[7], w1110, w1111);
  FullAdder U233 (w1111, w1082, IN24[6], w1112, w1113);
  FullAdder U234 (w1113, w1084, IN25[5], w1114, w1115);
  FullAdder U235 (w1115, w1086, IN26[4], w1116, w1117);
  FullAdder U236 (w1117, w1088, IN27[3], w1118, w1119);
  FullAdder U237 (w1119, w1090, IN28[2], w1120, w1121);
  FullAdder U238 (w1121, w1092, IN29[1], w1122, w1123);
  FullAdder U239 (w1123, w1093, IN30[0], w1124, w1125);
  HalfAdder U240 (w1096, IN16[16], Out1[16], w1127);
  FullAdder U241 (w1127, w1098, IN17[14], w1128, w1129);
  FullAdder U242 (w1129, w1100, IN18[13], w1130, w1131);
  FullAdder U243 (w1131, w1102, IN19[12], w1132, w1133);
  FullAdder U244 (w1133, w1104, IN20[11], w1134, w1135);
  FullAdder U245 (w1135, w1106, IN21[10], w1136, w1137);
  FullAdder U246 (w1137, w1108, IN22[9], w1138, w1139);
  FullAdder U247 (w1139, w1110, IN23[8], w1140, w1141);
  FullAdder U248 (w1141, w1112, IN24[7], w1142, w1143);
  FullAdder U249 (w1143, w1114, IN25[6], w1144, w1145);
  FullAdder U250 (w1145, w1116, IN26[5], w1146, w1147);
  FullAdder U251 (w1147, w1118, IN27[4], w1148, w1149);
  FullAdder U252 (w1149, w1120, IN28[3], w1150, w1151);
  FullAdder U253 (w1151, w1122, IN29[2], w1152, w1153);
  FullAdder U254 (w1153, w1124, IN30[1], w1154, w1155);
  FullAdder U255 (w1155, w1125, IN31[0], w1156, w1157);
  HalfAdder U256 (w1128, IN17[15], Out1[17], w1159);
  FullAdder U257 (w1159, w1130, IN18[14], w1160, w1161);
  FullAdder U258 (w1161, w1132, IN19[13], w1162, w1163);
  FullAdder U259 (w1163, w1134, IN20[12], w1164, w1165);
  FullAdder U260 (w1165, w1136, IN21[11], w1166, w1167);
  FullAdder U261 (w1167, w1138, IN22[10], w1168, w1169);
  FullAdder U262 (w1169, w1140, IN23[9], w1170, w1171);
  FullAdder U263 (w1171, w1142, IN24[8], w1172, w1173);
  FullAdder U264 (w1173, w1144, IN25[7], w1174, w1175);
  FullAdder U265 (w1175, w1146, IN26[6], w1176, w1177);
  FullAdder U266 (w1177, w1148, IN27[5], w1178, w1179);
  FullAdder U267 (w1179, w1150, IN28[4], w1180, w1181);
  FullAdder U268 (w1181, w1152, IN29[3], w1182, w1183);
  FullAdder U269 (w1183, w1154, IN30[2], w1184, w1185);
  FullAdder U270 (w1185, w1156, IN31[1], w1186, w1187);
  FullAdder U271 (w1187, w1157, IN32[0], w1188, w1189);
  HalfAdder U272 (w1160, IN18[15], Out1[18], w1191);
  FullAdder U273 (w1191, w1162, IN19[14], w1192, w1193);
  FullAdder U274 (w1193, w1164, IN20[13], w1194, w1195);
  FullAdder U275 (w1195, w1166, IN21[12], w1196, w1197);
  FullAdder U276 (w1197, w1168, IN22[11], w1198, w1199);
  FullAdder U277 (w1199, w1170, IN23[10], w1200, w1201);
  FullAdder U278 (w1201, w1172, IN24[9], w1202, w1203);
  FullAdder U279 (w1203, w1174, IN25[8], w1204, w1205);
  FullAdder U280 (w1205, w1176, IN26[7], w1206, w1207);
  FullAdder U281 (w1207, w1178, IN27[6], w1208, w1209);
  FullAdder U282 (w1209, w1180, IN28[5], w1210, w1211);
  FullAdder U283 (w1211, w1182, IN29[4], w1212, w1213);
  FullAdder U284 (w1213, w1184, IN30[3], w1214, w1215);
  FullAdder U285 (w1215, w1186, IN31[2], w1216, w1217);
  FullAdder U286 (w1217, w1188, IN32[1], w1218, w1219);
  FullAdder U287 (w1219, w1189, IN33[0], w1220, w1221);
  HalfAdder U288 (w1192, IN19[15], Out1[19], w1223);
  FullAdder U289 (w1223, w1194, IN20[14], w1224, w1225);
  FullAdder U290 (w1225, w1196, IN21[13], w1226, w1227);
  FullAdder U291 (w1227, w1198, IN22[12], w1228, w1229);
  FullAdder U292 (w1229, w1200, IN23[11], w1230, w1231);
  FullAdder U293 (w1231, w1202, IN24[10], w1232, w1233);
  FullAdder U294 (w1233, w1204, IN25[9], w1234, w1235);
  FullAdder U295 (w1235, w1206, IN26[8], w1236, w1237);
  FullAdder U296 (w1237, w1208, IN27[7], w1238, w1239);
  FullAdder U297 (w1239, w1210, IN28[6], w1240, w1241);
  FullAdder U298 (w1241, w1212, IN29[5], w1242, w1243);
  FullAdder U299 (w1243, w1214, IN30[4], w1244, w1245);
  FullAdder U300 (w1245, w1216, IN31[3], w1246, w1247);
  FullAdder U301 (w1247, w1218, IN32[2], w1248, w1249);
  FullAdder U302 (w1249, w1220, IN33[1], w1250, w1251);
  FullAdder U303 (w1251, w1221, IN34[0], w1252, w1253);
  HalfAdder U304 (w1224, IN20[15], Out1[20], w1255);
  FullAdder U305 (w1255, w1226, IN21[14], w1256, w1257);
  FullAdder U306 (w1257, w1228, IN22[13], w1258, w1259);
  FullAdder U307 (w1259, w1230, IN23[12], w1260, w1261);
  FullAdder U308 (w1261, w1232, IN24[11], w1262, w1263);
  FullAdder U309 (w1263, w1234, IN25[10], w1264, w1265);
  FullAdder U310 (w1265, w1236, IN26[9], w1266, w1267);
  FullAdder U311 (w1267, w1238, IN27[8], w1268, w1269);
  FullAdder U312 (w1269, w1240, IN28[7], w1270, w1271);
  FullAdder U313 (w1271, w1242, IN29[6], w1272, w1273);
  FullAdder U314 (w1273, w1244, IN30[5], w1274, w1275);
  FullAdder U315 (w1275, w1246, IN31[4], w1276, w1277);
  FullAdder U316 (w1277, w1248, IN32[3], w1278, w1279);
  FullAdder U317 (w1279, w1250, IN33[2], w1280, w1281);
  FullAdder U318 (w1281, w1252, IN34[1], w1282, w1283);
  FullAdder U319 (w1283, w1253, IN35[0], w1284, w1285);
  HalfAdder U320 (w1256, IN21[15], Out1[21], w1287);
  FullAdder U321 (w1287, w1258, IN22[14], w1288, w1289);
  FullAdder U322 (w1289, w1260, IN23[13], w1290, w1291);
  FullAdder U323 (w1291, w1262, IN24[12], w1292, w1293);
  FullAdder U324 (w1293, w1264, IN25[11], w1294, w1295);
  FullAdder U325 (w1295, w1266, IN26[10], w1296, w1297);
  FullAdder U326 (w1297, w1268, IN27[9], w1298, w1299);
  FullAdder U327 (w1299, w1270, IN28[8], w1300, w1301);
  FullAdder U328 (w1301, w1272, IN29[7], w1302, w1303);
  FullAdder U329 (w1303, w1274, IN30[6], w1304, w1305);
  FullAdder U330 (w1305, w1276, IN31[5], w1306, w1307);
  FullAdder U331 (w1307, w1278, IN32[4], w1308, w1309);
  FullAdder U332 (w1309, w1280, IN33[3], w1310, w1311);
  FullAdder U333 (w1311, w1282, IN34[2], w1312, w1313);
  FullAdder U334 (w1313, w1284, IN35[1], w1314, w1315);
  FullAdder U335 (w1315, w1285, IN36[0], w1316, w1317);
  HalfAdder U336 (w1288, IN22[15], Out1[22], w1319);
  FullAdder U337 (w1319, w1290, IN23[14], w1320, w1321);
  FullAdder U338 (w1321, w1292, IN24[13], w1322, w1323);
  FullAdder U339 (w1323, w1294, IN25[12], w1324, w1325);
  FullAdder U340 (w1325, w1296, IN26[11], w1326, w1327);
  FullAdder U341 (w1327, w1298, IN27[10], w1328, w1329);
  FullAdder U342 (w1329, w1300, IN28[9], w1330, w1331);
  FullAdder U343 (w1331, w1302, IN29[8], w1332, w1333);
  FullAdder U344 (w1333, w1304, IN30[7], w1334, w1335);
  FullAdder U345 (w1335, w1306, IN31[6], w1336, w1337);
  FullAdder U346 (w1337, w1308, IN32[5], w1338, w1339);
  FullAdder U347 (w1339, w1310, IN33[4], w1340, w1341);
  FullAdder U348 (w1341, w1312, IN34[3], w1342, w1343);
  FullAdder U349 (w1343, w1314, IN35[2], w1344, w1345);
  FullAdder U350 (w1345, w1316, IN36[1], w1346, w1347);
  FullAdder U351 (w1347, w1317, IN37[0], w1348, w1349);
  HalfAdder U352 (w1320, IN23[15], Out1[23], w1351);
  FullAdder U353 (w1351, w1322, IN24[14], w1352, w1353);
  FullAdder U354 (w1353, w1324, IN25[13], w1354, w1355);
  FullAdder U355 (w1355, w1326, IN26[12], w1356, w1357);
  FullAdder U356 (w1357, w1328, IN27[11], w1358, w1359);
  FullAdder U357 (w1359, w1330, IN28[10], w1360, w1361);
  FullAdder U358 (w1361, w1332, IN29[9], w1362, w1363);
  FullAdder U359 (w1363, w1334, IN30[8], w1364, w1365);
  FullAdder U360 (w1365, w1336, IN31[7], w1366, w1367);
  FullAdder U361 (w1367, w1338, IN32[6], w1368, w1369);
  FullAdder U362 (w1369, w1340, IN33[5], w1370, w1371);
  FullAdder U363 (w1371, w1342, IN34[4], w1372, w1373);
  FullAdder U364 (w1373, w1344, IN35[3], w1374, w1375);
  FullAdder U365 (w1375, w1346, IN36[2], w1376, w1377);
  FullAdder U366 (w1377, w1348, IN37[1], w1378, w1379);
  FullAdder U367 (w1379, w1349, IN38[0], w1380, w1381);
  HalfAdder U368 (w1352, IN24[15], Out1[24], w1383);
  FullAdder U369 (w1383, w1354, IN25[14], w1384, w1385);
  FullAdder U370 (w1385, w1356, IN26[13], w1386, w1387);
  FullAdder U371 (w1387, w1358, IN27[12], w1388, w1389);
  FullAdder U372 (w1389, w1360, IN28[11], w1390, w1391);
  FullAdder U373 (w1391, w1362, IN29[10], w1392, w1393);
  FullAdder U374 (w1393, w1364, IN30[9], w1394, w1395);
  FullAdder U375 (w1395, w1366, IN31[8], w1396, w1397);
  FullAdder U376 (w1397, w1368, IN32[7], w1398, w1399);
  FullAdder U377 (w1399, w1370, IN33[6], w1400, w1401);
  FullAdder U378 (w1401, w1372, IN34[5], w1402, w1403);
  FullAdder U379 (w1403, w1374, IN35[4], w1404, w1405);
  FullAdder U380 (w1405, w1376, IN36[3], w1406, w1407);
  FullAdder U381 (w1407, w1378, IN37[2], w1408, w1409);
  FullAdder U382 (w1409, w1380, IN38[1], w1410, w1411);
  FullAdder U383 (w1411, w1381, IN39[0], w1412, w1413);
  HalfAdder U384 (w1384, IN25[15], Out1[25], w1415);
  FullAdder U385 (w1415, w1386, IN26[14], w1416, w1417);
  FullAdder U386 (w1417, w1388, IN27[13], w1418, w1419);
  FullAdder U387 (w1419, w1390, IN28[12], w1420, w1421);
  FullAdder U388 (w1421, w1392, IN29[11], w1422, w1423);
  FullAdder U389 (w1423, w1394, IN30[10], w1424, w1425);
  FullAdder U390 (w1425, w1396, IN31[9], w1426, w1427);
  FullAdder U391 (w1427, w1398, IN32[8], w1428, w1429);
  FullAdder U392 (w1429, w1400, IN33[7], w1430, w1431);
  FullAdder U393 (w1431, w1402, IN34[6], w1432, w1433);
  FullAdder U394 (w1433, w1404, IN35[5], w1434, w1435);
  FullAdder U395 (w1435, w1406, IN36[4], w1436, w1437);
  FullAdder U396 (w1437, w1408, IN37[3], w1438, w1439);
  FullAdder U397 (w1439, w1410, IN38[2], w1440, w1441);
  FullAdder U398 (w1441, w1412, IN39[1], w1442, w1443);
  FullAdder U399 (w1443, w1413, IN40[0], w1444, w1445);
  HalfAdder U400 (w1416, IN26[15], Out1[26], w1447);
  FullAdder U401 (w1447, w1418, IN27[14], w1448, w1449);
  FullAdder U402 (w1449, w1420, IN28[13], w1450, w1451);
  FullAdder U403 (w1451, w1422, IN29[12], w1452, w1453);
  FullAdder U404 (w1453, w1424, IN30[11], w1454, w1455);
  FullAdder U405 (w1455, w1426, IN31[10], w1456, w1457);
  FullAdder U406 (w1457, w1428, IN32[9], w1458, w1459);
  FullAdder U407 (w1459, w1430, IN33[8], w1460, w1461);
  FullAdder U408 (w1461, w1432, IN34[7], w1462, w1463);
  FullAdder U409 (w1463, w1434, IN35[6], w1464, w1465);
  FullAdder U410 (w1465, w1436, IN36[5], w1466, w1467);
  FullAdder U411 (w1467, w1438, IN37[4], w1468, w1469);
  FullAdder U412 (w1469, w1440, IN38[3], w1470, w1471);
  FullAdder U413 (w1471, w1442, IN39[2], w1472, w1473);
  FullAdder U414 (w1473, w1444, IN40[1], w1474, w1475);
  FullAdder U415 (w1475, w1445, IN41[0], w1476, w1477);
  HalfAdder U416 (w1448, IN27[15], Out1[27], w1479);
  FullAdder U417 (w1479, w1450, IN28[14], w1480, w1481);
  FullAdder U418 (w1481, w1452, IN29[13], w1482, w1483);
  FullAdder U419 (w1483, w1454, IN30[12], w1484, w1485);
  FullAdder U420 (w1485, w1456, IN31[11], w1486, w1487);
  FullAdder U421 (w1487, w1458, IN32[10], w1488, w1489);
  FullAdder U422 (w1489, w1460, IN33[9], w1490, w1491);
  FullAdder U423 (w1491, w1462, IN34[8], w1492, w1493);
  FullAdder U424 (w1493, w1464, IN35[7], w1494, w1495);
  FullAdder U425 (w1495, w1466, IN36[6], w1496, w1497);
  FullAdder U426 (w1497, w1468, IN37[5], w1498, w1499);
  FullAdder U427 (w1499, w1470, IN38[4], w1500, w1501);
  FullAdder U428 (w1501, w1472, IN39[3], w1502, w1503);
  FullAdder U429 (w1503, w1474, IN40[2], w1504, w1505);
  FullAdder U430 (w1505, w1476, IN41[1], w1506, w1507);
  FullAdder U431 (w1507, w1477, IN42[0], w1508, w1509);
  HalfAdder U432 (w1480, IN28[15], Out1[28], w1511);
  FullAdder U433 (w1511, w1482, IN29[14], w1512, w1513);
  FullAdder U434 (w1513, w1484, IN30[13], w1514, w1515);
  FullAdder U435 (w1515, w1486, IN31[12], w1516, w1517);
  FullAdder U436 (w1517, w1488, IN32[11], w1518, w1519);
  FullAdder U437 (w1519, w1490, IN33[10], w1520, w1521);
  FullAdder U438 (w1521, w1492, IN34[9], w1522, w1523);
  FullAdder U439 (w1523, w1494, IN35[8], w1524, w1525);
  FullAdder U440 (w1525, w1496, IN36[7], w1526, w1527);
  FullAdder U441 (w1527, w1498, IN37[6], w1528, w1529);
  FullAdder U442 (w1529, w1500, IN38[5], w1530, w1531);
  FullAdder U443 (w1531, w1502, IN39[4], w1532, w1533);
  FullAdder U444 (w1533, w1504, IN40[3], w1534, w1535);
  FullAdder U445 (w1535, w1506, IN41[2], w1536, w1537);
  FullAdder U446 (w1537, w1508, IN42[1], w1538, w1539);
  FullAdder U447 (w1539, w1509, IN43[0], w1540, w1541);
  HalfAdder U448 (w1512, IN29[15], Out1[29], w1543);
  FullAdder U449 (w1543, w1514, IN30[14], w1544, w1545);
  FullAdder U450 (w1545, w1516, IN31[13], w1546, w1547);
  FullAdder U451 (w1547, w1518, IN32[12], w1548, w1549);
  FullAdder U452 (w1549, w1520, IN33[11], w1550, w1551);
  FullAdder U453 (w1551, w1522, IN34[10], w1552, w1553);
  FullAdder U454 (w1553, w1524, IN35[9], w1554, w1555);
  FullAdder U455 (w1555, w1526, IN36[8], w1556, w1557);
  FullAdder U456 (w1557, w1528, IN37[7], w1558, w1559);
  FullAdder U457 (w1559, w1530, IN38[6], w1560, w1561);
  FullAdder U458 (w1561, w1532, IN39[5], w1562, w1563);
  FullAdder U459 (w1563, w1534, IN40[4], w1564, w1565);
  FullAdder U460 (w1565, w1536, IN41[3], w1566, w1567);
  FullAdder U461 (w1567, w1538, IN42[2], w1568, w1569);
  FullAdder U462 (w1569, w1540, IN43[1], w1570, w1571);
  FullAdder U463 (w1571, w1541, IN44[0], w1572, w1573);
  HalfAdder U464 (w1544, IN30[15], Out1[30], w1575);
  FullAdder U465 (w1575, w1546, IN31[14], w1576, w1577);
  FullAdder U466 (w1577, w1548, IN32[13], w1578, w1579);
  FullAdder U467 (w1579, w1550, IN33[12], w1580, w1581);
  FullAdder U468 (w1581, w1552, IN34[11], w1582, w1583);
  FullAdder U469 (w1583, w1554, IN35[10], w1584, w1585);
  FullAdder U470 (w1585, w1556, IN36[9], w1586, w1587);
  FullAdder U471 (w1587, w1558, IN37[8], w1588, w1589);
  FullAdder U472 (w1589, w1560, IN38[7], w1590, w1591);
  FullAdder U473 (w1591, w1562, IN39[6], w1592, w1593);
  FullAdder U474 (w1593, w1564, IN40[5], w1594, w1595);
  FullAdder U475 (w1595, w1566, IN41[4], w1596, w1597);
  FullAdder U476 (w1597, w1568, IN42[3], w1598, w1599);
  FullAdder U477 (w1599, w1570, IN43[2], w1600, w1601);
  FullAdder U478 (w1601, w1572, IN44[1], w1602, w1603);
  FullAdder U479 (w1603, w1573, IN45[0], w1604, w1605);
  HalfAdder U480 (w1576, IN31[15], Out1[31], w1607);
  FullAdder U481 (w1607, w1578, IN32[14], w1608, w1609);
  FullAdder U482 (w1609, w1580, IN33[13], w1610, w1611);
  FullAdder U483 (w1611, w1582, IN34[12], w1612, w1613);
  FullAdder U484 (w1613, w1584, IN35[11], w1614, w1615);
  FullAdder U485 (w1615, w1586, IN36[10], w1616, w1617);
  FullAdder U486 (w1617, w1588, IN37[9], w1618, w1619);
  FullAdder U487 (w1619, w1590, IN38[8], w1620, w1621);
  FullAdder U488 (w1621, w1592, IN39[7], w1622, w1623);
  FullAdder U489 (w1623, w1594, IN40[6], w1624, w1625);
  FullAdder U490 (w1625, w1596, IN41[5], w1626, w1627);
  FullAdder U491 (w1627, w1598, IN42[4], w1628, w1629);
  FullAdder U492 (w1629, w1600, IN43[3], w1630, w1631);
  FullAdder U493 (w1631, w1602, IN44[2], w1632, w1633);
  FullAdder U494 (w1633, w1604, IN45[1], w1634, w1635);
  FullAdder U495 (w1635, w1605, IN46[0], w1636, w1637);
  HalfAdder U496 (w1608, IN32[15], Out1[32], w1639);
  FullAdder U497 (w1639, w1610, IN33[14], w1640, w1641);
  FullAdder U498 (w1641, w1612, IN34[13], w1642, w1643);
  FullAdder U499 (w1643, w1614, IN35[12], w1644, w1645);
  FullAdder U500 (w1645, w1616, IN36[11], w1646, w1647);
  FullAdder U501 (w1647, w1618, IN37[10], w1648, w1649);
  FullAdder U502 (w1649, w1620, IN38[9], w1650, w1651);
  FullAdder U503 (w1651, w1622, IN39[8], w1652, w1653);
  FullAdder U504 (w1653, w1624, IN40[7], w1654, w1655);
  FullAdder U505 (w1655, w1626, IN41[6], w1656, w1657);
  FullAdder U506 (w1657, w1628, IN42[5], w1658, w1659);
  FullAdder U507 (w1659, w1630, IN43[4], w1660, w1661);
  FullAdder U508 (w1661, w1632, IN44[3], w1662, w1663);
  FullAdder U509 (w1663, w1634, IN45[2], w1664, w1665);
  FullAdder U510 (w1665, w1636, IN46[1], w1666, w1667);
  FullAdder U511 (w1667, w1637, IN47[0], w1668, w1669);
  HalfAdder U512 (w1640, IN33[15], Out1[33], w1671);
  FullAdder U513 (w1671, w1642, IN34[14], w1672, w1673);
  FullAdder U514 (w1673, w1644, IN35[13], w1674, w1675);
  FullAdder U515 (w1675, w1646, IN36[12], w1676, w1677);
  FullAdder U516 (w1677, w1648, IN37[11], w1678, w1679);
  FullAdder U517 (w1679, w1650, IN38[10], w1680, w1681);
  FullAdder U518 (w1681, w1652, IN39[9], w1682, w1683);
  FullAdder U519 (w1683, w1654, IN40[8], w1684, w1685);
  FullAdder U520 (w1685, w1656, IN41[7], w1686, w1687);
  FullAdder U521 (w1687, w1658, IN42[6], w1688, w1689);
  FullAdder U522 (w1689, w1660, IN43[5], w1690, w1691);
  FullAdder U523 (w1691, w1662, IN44[4], w1692, w1693);
  FullAdder U524 (w1693, w1664, IN45[3], w1694, w1695);
  FullAdder U525 (w1695, w1666, IN46[2], w1696, w1697);
  FullAdder U526 (w1697, w1668, IN47[1], w1698, w1699);
  FullAdder U527 (w1699, w1669, IN48[0], w1700, w1701);
  HalfAdder U528 (w1672, IN34[15], Out1[34], w1703);
  FullAdder U529 (w1703, w1674, IN35[14], w1704, w1705);
  FullAdder U530 (w1705, w1676, IN36[13], w1706, w1707);
  FullAdder U531 (w1707, w1678, IN37[12], w1708, w1709);
  FullAdder U532 (w1709, w1680, IN38[11], w1710, w1711);
  FullAdder U533 (w1711, w1682, IN39[10], w1712, w1713);
  FullAdder U534 (w1713, w1684, IN40[9], w1714, w1715);
  FullAdder U535 (w1715, w1686, IN41[8], w1716, w1717);
  FullAdder U536 (w1717, w1688, IN42[7], w1718, w1719);
  FullAdder U537 (w1719, w1690, IN43[6], w1720, w1721);
  FullAdder U538 (w1721, w1692, IN44[5], w1722, w1723);
  FullAdder U539 (w1723, w1694, IN45[4], w1724, w1725);
  FullAdder U540 (w1725, w1696, IN46[3], w1726, w1727);
  FullAdder U541 (w1727, w1698, IN47[2], w1728, w1729);
  FullAdder U542 (w1729, w1700, IN48[1], w1730, w1731);
  FullAdder U543 (w1731, w1701, IN49[0], w1732, w1733);
  HalfAdder U544 (w1704, IN35[15], Out1[35], w1735);
  FullAdder U545 (w1735, w1706, IN36[14], w1736, w1737);
  FullAdder U546 (w1737, w1708, IN37[13], w1738, w1739);
  FullAdder U547 (w1739, w1710, IN38[12], w1740, w1741);
  FullAdder U548 (w1741, w1712, IN39[11], w1742, w1743);
  FullAdder U549 (w1743, w1714, IN40[10], w1744, w1745);
  FullAdder U550 (w1745, w1716, IN41[9], w1746, w1747);
  FullAdder U551 (w1747, w1718, IN42[8], w1748, w1749);
  FullAdder U552 (w1749, w1720, IN43[7], w1750, w1751);
  FullAdder U553 (w1751, w1722, IN44[6], w1752, w1753);
  FullAdder U554 (w1753, w1724, IN45[5], w1754, w1755);
  FullAdder U555 (w1755, w1726, IN46[4], w1756, w1757);
  FullAdder U556 (w1757, w1728, IN47[3], w1758, w1759);
  FullAdder U557 (w1759, w1730, IN48[2], w1760, w1761);
  FullAdder U558 (w1761, w1732, IN49[1], w1762, w1763);
  FullAdder U559 (w1763, w1733, IN50[0], w1764, w1765);
  HalfAdder U560 (w1736, IN36[15], Out1[36], w1767);
  FullAdder U561 (w1767, w1738, IN37[14], w1768, w1769);
  FullAdder U562 (w1769, w1740, IN38[13], w1770, w1771);
  FullAdder U563 (w1771, w1742, IN39[12], w1772, w1773);
  FullAdder U564 (w1773, w1744, IN40[11], w1774, w1775);
  FullAdder U565 (w1775, w1746, IN41[10], w1776, w1777);
  FullAdder U566 (w1777, w1748, IN42[9], w1778, w1779);
  FullAdder U567 (w1779, w1750, IN43[8], w1780, w1781);
  FullAdder U568 (w1781, w1752, IN44[7], w1782, w1783);
  FullAdder U569 (w1783, w1754, IN45[6], w1784, w1785);
  FullAdder U570 (w1785, w1756, IN46[5], w1786, w1787);
  FullAdder U571 (w1787, w1758, IN47[4], w1788, w1789);
  FullAdder U572 (w1789, w1760, IN48[3], w1790, w1791);
  FullAdder U573 (w1791, w1762, IN49[2], w1792, w1793);
  FullAdder U574 (w1793, w1764, IN50[1], w1794, w1795);
  FullAdder U575 (w1795, w1765, IN51[0], w1796, w1797);
  HalfAdder U576 (w1768, IN37[15], Out1[37], w1799);
  FullAdder U577 (w1799, w1770, IN38[14], Out1[38], w1801);
  FullAdder U578 (w1801, w1772, IN39[13], Out1[39], w1803);
  FullAdder U579 (w1803, w1774, IN40[12], Out1[40], w1805);
  FullAdder U580 (w1805, w1776, IN41[11], Out1[41], w1807);
  FullAdder U581 (w1807, w1778, IN42[10], Out1[42], w1809);
  FullAdder U582 (w1809, w1780, IN43[9], Out1[43], w1811);
  FullAdder U583 (w1811, w1782, IN44[8], Out1[44], w1813);
  FullAdder U584 (w1813, w1784, IN45[7], Out1[45], w1815);
  FullAdder U585 (w1815, w1786, IN46[6], Out1[46], w1817);
  FullAdder U586 (w1817, w1788, IN47[5], Out1[47], w1819);
  FullAdder U587 (w1819, w1790, IN48[4], Out1[48], w1821);
  FullAdder U588 (w1821, w1792, IN49[3], Out1[49], w1823);
  FullAdder U589 (w1823, w1794, IN50[2], Out1[50], w1825);
  FullAdder U590 (w1825, w1796, IN51[1], Out1[51], w1827);
  FullAdder U591 (w1827, w1797, IN52[0], Out1[52], Out1[53]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN17[16];
  assign Out2[1] = IN18[16];
  assign Out2[2] = IN19[16];
  assign Out2[3] = IN20[16];
  assign Out2[4] = IN21[16];
  assign Out2[5] = IN22[16];
  assign Out2[6] = IN23[16];
  assign Out2[7] = IN24[16];
  assign Out2[8] = IN25[16];
  assign Out2[9] = IN26[16];
  assign Out2[10] = IN27[16];
  assign Out2[11] = IN28[16];
  assign Out2[12] = IN29[16];
  assign Out2[13] = IN30[16];
  assign Out2[14] = IN31[16];
  assign Out2[15] = IN32[16];
  assign Out2[16] = IN33[16];
  assign Out2[17] = IN34[16];
  assign Out2[18] = IN35[16];
  assign Out2[19] = IN36[16];
  assign Out2[20] = IN37[16];
  assign Out2[21] = IN38[15];
  assign Out2[22] = IN39[14];
  assign Out2[23] = IN40[13];
  assign Out2[24] = IN41[12];
  assign Out2[25] = IN42[11];
  assign Out2[26] = IN43[10];
  assign Out2[27] = IN44[9];
  assign Out2[28] = IN45[8];
  assign Out2[29] = IN46[7];
  assign Out2[30] = IN47[6];
  assign Out2[31] = IN48[5];
  assign Out2[32] = IN49[4];
  assign Out2[33] = IN50[3];
  assign Out2[34] = IN51[2];
  assign Out2[35] = IN52[1];
  assign Out2[36] = IN53[0];

endmodule
module RC_37_37(IN1, IN2, Out);
  input [36:0] IN1;
  input [36:0] IN2;
  output [37:0] Out;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w75);
  FullAdder U1 (IN1[1], IN2[1], w75, Out[1], w77);
  FullAdder U2 (IN1[2], IN2[2], w77, Out[2], w79);
  FullAdder U3 (IN1[3], IN2[3], w79, Out[3], w81);
  FullAdder U4 (IN1[4], IN2[4], w81, Out[4], w83);
  FullAdder U5 (IN1[5], IN2[5], w83, Out[5], w85);
  FullAdder U6 (IN1[6], IN2[6], w85, Out[6], w87);
  FullAdder U7 (IN1[7], IN2[7], w87, Out[7], w89);
  FullAdder U8 (IN1[8], IN2[8], w89, Out[8], w91);
  FullAdder U9 (IN1[9], IN2[9], w91, Out[9], w93);
  FullAdder U10 (IN1[10], IN2[10], w93, Out[10], w95);
  FullAdder U11 (IN1[11], IN2[11], w95, Out[11], w97);
  FullAdder U12 (IN1[12], IN2[12], w97, Out[12], w99);
  FullAdder U13 (IN1[13], IN2[13], w99, Out[13], w101);
  FullAdder U14 (IN1[14], IN2[14], w101, Out[14], w103);
  FullAdder U15 (IN1[15], IN2[15], w103, Out[15], w105);
  FullAdder U16 (IN1[16], IN2[16], w105, Out[16], w107);
  FullAdder U17 (IN1[17], IN2[17], w107, Out[17], w109);
  FullAdder U18 (IN1[18], IN2[18], w109, Out[18], w111);
  FullAdder U19 (IN1[19], IN2[19], w111, Out[19], w113);
  FullAdder U20 (IN1[20], IN2[20], w113, Out[20], w115);
  FullAdder U21 (IN1[21], IN2[21], w115, Out[21], w117);
  FullAdder U22 (IN1[22], IN2[22], w117, Out[22], w119);
  FullAdder U23 (IN1[23], IN2[23], w119, Out[23], w121);
  FullAdder U24 (IN1[24], IN2[24], w121, Out[24], w123);
  FullAdder U25 (IN1[25], IN2[25], w123, Out[25], w125);
  FullAdder U26 (IN1[26], IN2[26], w125, Out[26], w127);
  FullAdder U27 (IN1[27], IN2[27], w127, Out[27], w129);
  FullAdder U28 (IN1[28], IN2[28], w129, Out[28], w131);
  FullAdder U29 (IN1[29], IN2[29], w131, Out[29], w133);
  FullAdder U30 (IN1[30], IN2[30], w133, Out[30], w135);
  FullAdder U31 (IN1[31], IN2[31], w135, Out[31], w137);
  FullAdder U32 (IN1[32], IN2[32], w137, Out[32], w139);
  FullAdder U33 (IN1[33], IN2[33], w139, Out[33], w141);
  FullAdder U34 (IN1[34], IN2[34], w141, Out[34], w143);
  FullAdder U35 (IN1[35], IN2[35], w143, Out[35], w145);
  FullAdder U36 (IN1[36], IN2[36], w145, Out[36], Out[37]);

endmodule
module NR_17_38(IN1, IN2, Out);
  input [16:0] IN1;
  input [37:0] IN2;
  output [54:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [16:0] P17;
  wire [16:0] P18;
  wire [16:0] P19;
  wire [16:0] P20;
  wire [16:0] P21;
  wire [16:0] P22;
  wire [16:0] P23;
  wire [16:0] P24;
  wire [16:0] P25;
  wire [16:0] P26;
  wire [16:0] P27;
  wire [16:0] P28;
  wire [16:0] P29;
  wire [16:0] P30;
  wire [16:0] P31;
  wire [16:0] P32;
  wire [16:0] P33;
  wire [16:0] P34;
  wire [16:0] P35;
  wire [16:0] P36;
  wire [16:0] P37;
  wire [15:0] P38;
  wire [14:0] P39;
  wire [13:0] P40;
  wire [12:0] P41;
  wire [11:0] P42;
  wire [10:0] P43;
  wire [9:0] P44;
  wire [8:0] P45;
  wire [7:0] P46;
  wire [6:0] P47;
  wire [5:0] P48;
  wire [4:0] P49;
  wire [3:0] P50;
  wire [2:0] P51;
  wire [1:0] P52;
  wire [0:0] P53;
  wire [53:0] R1;
  wire [36:0] R2;
  wire [54:0] aOut;
  U_SP_17_38 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, R1, R2);
  RC_37_37 S2 (R1[53:17], R2, aOut[54:17]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign Out = aOut[54:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
