//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 53
  second input length: 53
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_53_53(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104);
  input [52:0] IN1;
  input [52:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [29:0] P29;
  output [30:0] P30;
  output [31:0] P31;
  output [32:0] P32;
  output [33:0] P33;
  output [34:0] P34;
  output [35:0] P35;
  output [36:0] P36;
  output [37:0] P37;
  output [38:0] P38;
  output [39:0] P39;
  output [40:0] P40;
  output [41:0] P41;
  output [42:0] P42;
  output [43:0] P43;
  output [44:0] P44;
  output [45:0] P45;
  output [46:0] P46;
  output [47:0] P47;
  output [48:0] P48;
  output [49:0] P49;
  output [50:0] P50;
  output [51:0] P51;
  output [52:0] P52;
  output [51:0] P53;
  output [50:0] P54;
  output [49:0] P55;
  output [48:0] P56;
  output [47:0] P57;
  output [46:0] P58;
  output [45:0] P59;
  output [44:0] P60;
  output [43:0] P61;
  output [42:0] P62;
  output [41:0] P63;
  output [40:0] P64;
  output [39:0] P65;
  output [38:0] P66;
  output [37:0] P67;
  output [36:0] P68;
  output [35:0] P69;
  output [34:0] P70;
  output [33:0] P71;
  output [32:0] P72;
  output [31:0] P73;
  output [30:0] P74;
  output [29:0] P75;
  output [28:0] P76;
  output [27:0] P77;
  output [26:0] P78;
  output [25:0] P79;
  output [24:0] P80;
  output [23:0] P81;
  output [22:0] P82;
  output [21:0] P83;
  output [20:0] P84;
  output [19:0] P85;
  output [18:0] P86;
  output [17:0] P87;
  output [16:0] P88;
  output [15:0] P89;
  output [14:0] P90;
  output [13:0] P91;
  output [12:0] P92;
  output [11:0] P93;
  output [10:0] P94;
  output [9:0] P95;
  output [8:0] P96;
  output [7:0] P97;
  output [6:0] P98;
  output [5:0] P99;
  output [4:0] P100;
  output [3:0] P101;
  output [2:0] P102;
  output [1:0] P103;
  output [0:0] P104;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[0] = IN1[1]&IN2[52];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[1] = IN1[2]&IN2[51];
  assign P54[0] = IN1[2]&IN2[52];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[2] = IN1[3]&IN2[50];
  assign P54[1] = IN1[3]&IN2[51];
  assign P55[0] = IN1[3]&IN2[52];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[3] = IN1[4]&IN2[49];
  assign P54[2] = IN1[4]&IN2[50];
  assign P55[1] = IN1[4]&IN2[51];
  assign P56[0] = IN1[4]&IN2[52];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[4] = IN1[5]&IN2[48];
  assign P54[3] = IN1[5]&IN2[49];
  assign P55[2] = IN1[5]&IN2[50];
  assign P56[1] = IN1[5]&IN2[51];
  assign P57[0] = IN1[5]&IN2[52];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[5] = IN1[6]&IN2[47];
  assign P54[4] = IN1[6]&IN2[48];
  assign P55[3] = IN1[6]&IN2[49];
  assign P56[2] = IN1[6]&IN2[50];
  assign P57[1] = IN1[6]&IN2[51];
  assign P58[0] = IN1[6]&IN2[52];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[6] = IN1[7]&IN2[46];
  assign P54[5] = IN1[7]&IN2[47];
  assign P55[4] = IN1[7]&IN2[48];
  assign P56[3] = IN1[7]&IN2[49];
  assign P57[2] = IN1[7]&IN2[50];
  assign P58[1] = IN1[7]&IN2[51];
  assign P59[0] = IN1[7]&IN2[52];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[7] = IN1[8]&IN2[45];
  assign P54[6] = IN1[8]&IN2[46];
  assign P55[5] = IN1[8]&IN2[47];
  assign P56[4] = IN1[8]&IN2[48];
  assign P57[3] = IN1[8]&IN2[49];
  assign P58[2] = IN1[8]&IN2[50];
  assign P59[1] = IN1[8]&IN2[51];
  assign P60[0] = IN1[8]&IN2[52];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[8] = IN1[9]&IN2[44];
  assign P54[7] = IN1[9]&IN2[45];
  assign P55[6] = IN1[9]&IN2[46];
  assign P56[5] = IN1[9]&IN2[47];
  assign P57[4] = IN1[9]&IN2[48];
  assign P58[3] = IN1[9]&IN2[49];
  assign P59[2] = IN1[9]&IN2[50];
  assign P60[1] = IN1[9]&IN2[51];
  assign P61[0] = IN1[9]&IN2[52];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[10] = IN1[10]&IN2[39];
  assign P50[10] = IN1[10]&IN2[40];
  assign P51[10] = IN1[10]&IN2[41];
  assign P52[10] = IN1[10]&IN2[42];
  assign P53[9] = IN1[10]&IN2[43];
  assign P54[8] = IN1[10]&IN2[44];
  assign P55[7] = IN1[10]&IN2[45];
  assign P56[6] = IN1[10]&IN2[46];
  assign P57[5] = IN1[10]&IN2[47];
  assign P58[4] = IN1[10]&IN2[48];
  assign P59[3] = IN1[10]&IN2[49];
  assign P60[2] = IN1[10]&IN2[50];
  assign P61[1] = IN1[10]&IN2[51];
  assign P62[0] = IN1[10]&IN2[52];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[11] = IN1[11]&IN2[38];
  assign P50[11] = IN1[11]&IN2[39];
  assign P51[11] = IN1[11]&IN2[40];
  assign P52[11] = IN1[11]&IN2[41];
  assign P53[10] = IN1[11]&IN2[42];
  assign P54[9] = IN1[11]&IN2[43];
  assign P55[8] = IN1[11]&IN2[44];
  assign P56[7] = IN1[11]&IN2[45];
  assign P57[6] = IN1[11]&IN2[46];
  assign P58[5] = IN1[11]&IN2[47];
  assign P59[4] = IN1[11]&IN2[48];
  assign P60[3] = IN1[11]&IN2[49];
  assign P61[2] = IN1[11]&IN2[50];
  assign P62[1] = IN1[11]&IN2[51];
  assign P63[0] = IN1[11]&IN2[52];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[12] = IN1[12]&IN2[37];
  assign P50[12] = IN1[12]&IN2[38];
  assign P51[12] = IN1[12]&IN2[39];
  assign P52[12] = IN1[12]&IN2[40];
  assign P53[11] = IN1[12]&IN2[41];
  assign P54[10] = IN1[12]&IN2[42];
  assign P55[9] = IN1[12]&IN2[43];
  assign P56[8] = IN1[12]&IN2[44];
  assign P57[7] = IN1[12]&IN2[45];
  assign P58[6] = IN1[12]&IN2[46];
  assign P59[5] = IN1[12]&IN2[47];
  assign P60[4] = IN1[12]&IN2[48];
  assign P61[3] = IN1[12]&IN2[49];
  assign P62[2] = IN1[12]&IN2[50];
  assign P63[1] = IN1[12]&IN2[51];
  assign P64[0] = IN1[12]&IN2[52];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[13] = IN1[13]&IN2[36];
  assign P50[13] = IN1[13]&IN2[37];
  assign P51[13] = IN1[13]&IN2[38];
  assign P52[13] = IN1[13]&IN2[39];
  assign P53[12] = IN1[13]&IN2[40];
  assign P54[11] = IN1[13]&IN2[41];
  assign P55[10] = IN1[13]&IN2[42];
  assign P56[9] = IN1[13]&IN2[43];
  assign P57[8] = IN1[13]&IN2[44];
  assign P58[7] = IN1[13]&IN2[45];
  assign P59[6] = IN1[13]&IN2[46];
  assign P60[5] = IN1[13]&IN2[47];
  assign P61[4] = IN1[13]&IN2[48];
  assign P62[3] = IN1[13]&IN2[49];
  assign P63[2] = IN1[13]&IN2[50];
  assign P64[1] = IN1[13]&IN2[51];
  assign P65[0] = IN1[13]&IN2[52];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[14] = IN1[14]&IN2[24];
  assign P39[14] = IN1[14]&IN2[25];
  assign P40[14] = IN1[14]&IN2[26];
  assign P41[14] = IN1[14]&IN2[27];
  assign P42[14] = IN1[14]&IN2[28];
  assign P43[14] = IN1[14]&IN2[29];
  assign P44[14] = IN1[14]&IN2[30];
  assign P45[14] = IN1[14]&IN2[31];
  assign P46[14] = IN1[14]&IN2[32];
  assign P47[14] = IN1[14]&IN2[33];
  assign P48[14] = IN1[14]&IN2[34];
  assign P49[14] = IN1[14]&IN2[35];
  assign P50[14] = IN1[14]&IN2[36];
  assign P51[14] = IN1[14]&IN2[37];
  assign P52[14] = IN1[14]&IN2[38];
  assign P53[13] = IN1[14]&IN2[39];
  assign P54[12] = IN1[14]&IN2[40];
  assign P55[11] = IN1[14]&IN2[41];
  assign P56[10] = IN1[14]&IN2[42];
  assign P57[9] = IN1[14]&IN2[43];
  assign P58[8] = IN1[14]&IN2[44];
  assign P59[7] = IN1[14]&IN2[45];
  assign P60[6] = IN1[14]&IN2[46];
  assign P61[5] = IN1[14]&IN2[47];
  assign P62[4] = IN1[14]&IN2[48];
  assign P63[3] = IN1[14]&IN2[49];
  assign P64[2] = IN1[14]&IN2[50];
  assign P65[1] = IN1[14]&IN2[51];
  assign P66[0] = IN1[14]&IN2[52];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[15] = IN1[15]&IN2[23];
  assign P39[15] = IN1[15]&IN2[24];
  assign P40[15] = IN1[15]&IN2[25];
  assign P41[15] = IN1[15]&IN2[26];
  assign P42[15] = IN1[15]&IN2[27];
  assign P43[15] = IN1[15]&IN2[28];
  assign P44[15] = IN1[15]&IN2[29];
  assign P45[15] = IN1[15]&IN2[30];
  assign P46[15] = IN1[15]&IN2[31];
  assign P47[15] = IN1[15]&IN2[32];
  assign P48[15] = IN1[15]&IN2[33];
  assign P49[15] = IN1[15]&IN2[34];
  assign P50[15] = IN1[15]&IN2[35];
  assign P51[15] = IN1[15]&IN2[36];
  assign P52[15] = IN1[15]&IN2[37];
  assign P53[14] = IN1[15]&IN2[38];
  assign P54[13] = IN1[15]&IN2[39];
  assign P55[12] = IN1[15]&IN2[40];
  assign P56[11] = IN1[15]&IN2[41];
  assign P57[10] = IN1[15]&IN2[42];
  assign P58[9] = IN1[15]&IN2[43];
  assign P59[8] = IN1[15]&IN2[44];
  assign P60[7] = IN1[15]&IN2[45];
  assign P61[6] = IN1[15]&IN2[46];
  assign P62[5] = IN1[15]&IN2[47];
  assign P63[4] = IN1[15]&IN2[48];
  assign P64[3] = IN1[15]&IN2[49];
  assign P65[2] = IN1[15]&IN2[50];
  assign P66[1] = IN1[15]&IN2[51];
  assign P67[0] = IN1[15]&IN2[52];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[16] = IN1[16]&IN2[22];
  assign P39[16] = IN1[16]&IN2[23];
  assign P40[16] = IN1[16]&IN2[24];
  assign P41[16] = IN1[16]&IN2[25];
  assign P42[16] = IN1[16]&IN2[26];
  assign P43[16] = IN1[16]&IN2[27];
  assign P44[16] = IN1[16]&IN2[28];
  assign P45[16] = IN1[16]&IN2[29];
  assign P46[16] = IN1[16]&IN2[30];
  assign P47[16] = IN1[16]&IN2[31];
  assign P48[16] = IN1[16]&IN2[32];
  assign P49[16] = IN1[16]&IN2[33];
  assign P50[16] = IN1[16]&IN2[34];
  assign P51[16] = IN1[16]&IN2[35];
  assign P52[16] = IN1[16]&IN2[36];
  assign P53[15] = IN1[16]&IN2[37];
  assign P54[14] = IN1[16]&IN2[38];
  assign P55[13] = IN1[16]&IN2[39];
  assign P56[12] = IN1[16]&IN2[40];
  assign P57[11] = IN1[16]&IN2[41];
  assign P58[10] = IN1[16]&IN2[42];
  assign P59[9] = IN1[16]&IN2[43];
  assign P60[8] = IN1[16]&IN2[44];
  assign P61[7] = IN1[16]&IN2[45];
  assign P62[6] = IN1[16]&IN2[46];
  assign P63[5] = IN1[16]&IN2[47];
  assign P64[4] = IN1[16]&IN2[48];
  assign P65[3] = IN1[16]&IN2[49];
  assign P66[2] = IN1[16]&IN2[50];
  assign P67[1] = IN1[16]&IN2[51];
  assign P68[0] = IN1[16]&IN2[52];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[17] = IN1[17]&IN2[21];
  assign P39[17] = IN1[17]&IN2[22];
  assign P40[17] = IN1[17]&IN2[23];
  assign P41[17] = IN1[17]&IN2[24];
  assign P42[17] = IN1[17]&IN2[25];
  assign P43[17] = IN1[17]&IN2[26];
  assign P44[17] = IN1[17]&IN2[27];
  assign P45[17] = IN1[17]&IN2[28];
  assign P46[17] = IN1[17]&IN2[29];
  assign P47[17] = IN1[17]&IN2[30];
  assign P48[17] = IN1[17]&IN2[31];
  assign P49[17] = IN1[17]&IN2[32];
  assign P50[17] = IN1[17]&IN2[33];
  assign P51[17] = IN1[17]&IN2[34];
  assign P52[17] = IN1[17]&IN2[35];
  assign P53[16] = IN1[17]&IN2[36];
  assign P54[15] = IN1[17]&IN2[37];
  assign P55[14] = IN1[17]&IN2[38];
  assign P56[13] = IN1[17]&IN2[39];
  assign P57[12] = IN1[17]&IN2[40];
  assign P58[11] = IN1[17]&IN2[41];
  assign P59[10] = IN1[17]&IN2[42];
  assign P60[9] = IN1[17]&IN2[43];
  assign P61[8] = IN1[17]&IN2[44];
  assign P62[7] = IN1[17]&IN2[45];
  assign P63[6] = IN1[17]&IN2[46];
  assign P64[5] = IN1[17]&IN2[47];
  assign P65[4] = IN1[17]&IN2[48];
  assign P66[3] = IN1[17]&IN2[49];
  assign P67[2] = IN1[17]&IN2[50];
  assign P68[1] = IN1[17]&IN2[51];
  assign P69[0] = IN1[17]&IN2[52];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[18] = IN1[18]&IN2[20];
  assign P39[18] = IN1[18]&IN2[21];
  assign P40[18] = IN1[18]&IN2[22];
  assign P41[18] = IN1[18]&IN2[23];
  assign P42[18] = IN1[18]&IN2[24];
  assign P43[18] = IN1[18]&IN2[25];
  assign P44[18] = IN1[18]&IN2[26];
  assign P45[18] = IN1[18]&IN2[27];
  assign P46[18] = IN1[18]&IN2[28];
  assign P47[18] = IN1[18]&IN2[29];
  assign P48[18] = IN1[18]&IN2[30];
  assign P49[18] = IN1[18]&IN2[31];
  assign P50[18] = IN1[18]&IN2[32];
  assign P51[18] = IN1[18]&IN2[33];
  assign P52[18] = IN1[18]&IN2[34];
  assign P53[17] = IN1[18]&IN2[35];
  assign P54[16] = IN1[18]&IN2[36];
  assign P55[15] = IN1[18]&IN2[37];
  assign P56[14] = IN1[18]&IN2[38];
  assign P57[13] = IN1[18]&IN2[39];
  assign P58[12] = IN1[18]&IN2[40];
  assign P59[11] = IN1[18]&IN2[41];
  assign P60[10] = IN1[18]&IN2[42];
  assign P61[9] = IN1[18]&IN2[43];
  assign P62[8] = IN1[18]&IN2[44];
  assign P63[7] = IN1[18]&IN2[45];
  assign P64[6] = IN1[18]&IN2[46];
  assign P65[5] = IN1[18]&IN2[47];
  assign P66[4] = IN1[18]&IN2[48];
  assign P67[3] = IN1[18]&IN2[49];
  assign P68[2] = IN1[18]&IN2[50];
  assign P69[1] = IN1[18]&IN2[51];
  assign P70[0] = IN1[18]&IN2[52];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[19] = IN1[19]&IN2[19];
  assign P39[19] = IN1[19]&IN2[20];
  assign P40[19] = IN1[19]&IN2[21];
  assign P41[19] = IN1[19]&IN2[22];
  assign P42[19] = IN1[19]&IN2[23];
  assign P43[19] = IN1[19]&IN2[24];
  assign P44[19] = IN1[19]&IN2[25];
  assign P45[19] = IN1[19]&IN2[26];
  assign P46[19] = IN1[19]&IN2[27];
  assign P47[19] = IN1[19]&IN2[28];
  assign P48[19] = IN1[19]&IN2[29];
  assign P49[19] = IN1[19]&IN2[30];
  assign P50[19] = IN1[19]&IN2[31];
  assign P51[19] = IN1[19]&IN2[32];
  assign P52[19] = IN1[19]&IN2[33];
  assign P53[18] = IN1[19]&IN2[34];
  assign P54[17] = IN1[19]&IN2[35];
  assign P55[16] = IN1[19]&IN2[36];
  assign P56[15] = IN1[19]&IN2[37];
  assign P57[14] = IN1[19]&IN2[38];
  assign P58[13] = IN1[19]&IN2[39];
  assign P59[12] = IN1[19]&IN2[40];
  assign P60[11] = IN1[19]&IN2[41];
  assign P61[10] = IN1[19]&IN2[42];
  assign P62[9] = IN1[19]&IN2[43];
  assign P63[8] = IN1[19]&IN2[44];
  assign P64[7] = IN1[19]&IN2[45];
  assign P65[6] = IN1[19]&IN2[46];
  assign P66[5] = IN1[19]&IN2[47];
  assign P67[4] = IN1[19]&IN2[48];
  assign P68[3] = IN1[19]&IN2[49];
  assign P69[2] = IN1[19]&IN2[50];
  assign P70[1] = IN1[19]&IN2[51];
  assign P71[0] = IN1[19]&IN2[52];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[20] = IN1[20]&IN2[18];
  assign P39[20] = IN1[20]&IN2[19];
  assign P40[20] = IN1[20]&IN2[20];
  assign P41[20] = IN1[20]&IN2[21];
  assign P42[20] = IN1[20]&IN2[22];
  assign P43[20] = IN1[20]&IN2[23];
  assign P44[20] = IN1[20]&IN2[24];
  assign P45[20] = IN1[20]&IN2[25];
  assign P46[20] = IN1[20]&IN2[26];
  assign P47[20] = IN1[20]&IN2[27];
  assign P48[20] = IN1[20]&IN2[28];
  assign P49[20] = IN1[20]&IN2[29];
  assign P50[20] = IN1[20]&IN2[30];
  assign P51[20] = IN1[20]&IN2[31];
  assign P52[20] = IN1[20]&IN2[32];
  assign P53[19] = IN1[20]&IN2[33];
  assign P54[18] = IN1[20]&IN2[34];
  assign P55[17] = IN1[20]&IN2[35];
  assign P56[16] = IN1[20]&IN2[36];
  assign P57[15] = IN1[20]&IN2[37];
  assign P58[14] = IN1[20]&IN2[38];
  assign P59[13] = IN1[20]&IN2[39];
  assign P60[12] = IN1[20]&IN2[40];
  assign P61[11] = IN1[20]&IN2[41];
  assign P62[10] = IN1[20]&IN2[42];
  assign P63[9] = IN1[20]&IN2[43];
  assign P64[8] = IN1[20]&IN2[44];
  assign P65[7] = IN1[20]&IN2[45];
  assign P66[6] = IN1[20]&IN2[46];
  assign P67[5] = IN1[20]&IN2[47];
  assign P68[4] = IN1[20]&IN2[48];
  assign P69[3] = IN1[20]&IN2[49];
  assign P70[2] = IN1[20]&IN2[50];
  assign P71[1] = IN1[20]&IN2[51];
  assign P72[0] = IN1[20]&IN2[52];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[21] = IN1[21]&IN2[14];
  assign P36[21] = IN1[21]&IN2[15];
  assign P37[21] = IN1[21]&IN2[16];
  assign P38[21] = IN1[21]&IN2[17];
  assign P39[21] = IN1[21]&IN2[18];
  assign P40[21] = IN1[21]&IN2[19];
  assign P41[21] = IN1[21]&IN2[20];
  assign P42[21] = IN1[21]&IN2[21];
  assign P43[21] = IN1[21]&IN2[22];
  assign P44[21] = IN1[21]&IN2[23];
  assign P45[21] = IN1[21]&IN2[24];
  assign P46[21] = IN1[21]&IN2[25];
  assign P47[21] = IN1[21]&IN2[26];
  assign P48[21] = IN1[21]&IN2[27];
  assign P49[21] = IN1[21]&IN2[28];
  assign P50[21] = IN1[21]&IN2[29];
  assign P51[21] = IN1[21]&IN2[30];
  assign P52[21] = IN1[21]&IN2[31];
  assign P53[20] = IN1[21]&IN2[32];
  assign P54[19] = IN1[21]&IN2[33];
  assign P55[18] = IN1[21]&IN2[34];
  assign P56[17] = IN1[21]&IN2[35];
  assign P57[16] = IN1[21]&IN2[36];
  assign P58[15] = IN1[21]&IN2[37];
  assign P59[14] = IN1[21]&IN2[38];
  assign P60[13] = IN1[21]&IN2[39];
  assign P61[12] = IN1[21]&IN2[40];
  assign P62[11] = IN1[21]&IN2[41];
  assign P63[10] = IN1[21]&IN2[42];
  assign P64[9] = IN1[21]&IN2[43];
  assign P65[8] = IN1[21]&IN2[44];
  assign P66[7] = IN1[21]&IN2[45];
  assign P67[6] = IN1[21]&IN2[46];
  assign P68[5] = IN1[21]&IN2[47];
  assign P69[4] = IN1[21]&IN2[48];
  assign P70[3] = IN1[21]&IN2[49];
  assign P71[2] = IN1[21]&IN2[50];
  assign P72[1] = IN1[21]&IN2[51];
  assign P73[0] = IN1[21]&IN2[52];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[22] = IN1[22]&IN2[13];
  assign P36[22] = IN1[22]&IN2[14];
  assign P37[22] = IN1[22]&IN2[15];
  assign P38[22] = IN1[22]&IN2[16];
  assign P39[22] = IN1[22]&IN2[17];
  assign P40[22] = IN1[22]&IN2[18];
  assign P41[22] = IN1[22]&IN2[19];
  assign P42[22] = IN1[22]&IN2[20];
  assign P43[22] = IN1[22]&IN2[21];
  assign P44[22] = IN1[22]&IN2[22];
  assign P45[22] = IN1[22]&IN2[23];
  assign P46[22] = IN1[22]&IN2[24];
  assign P47[22] = IN1[22]&IN2[25];
  assign P48[22] = IN1[22]&IN2[26];
  assign P49[22] = IN1[22]&IN2[27];
  assign P50[22] = IN1[22]&IN2[28];
  assign P51[22] = IN1[22]&IN2[29];
  assign P52[22] = IN1[22]&IN2[30];
  assign P53[21] = IN1[22]&IN2[31];
  assign P54[20] = IN1[22]&IN2[32];
  assign P55[19] = IN1[22]&IN2[33];
  assign P56[18] = IN1[22]&IN2[34];
  assign P57[17] = IN1[22]&IN2[35];
  assign P58[16] = IN1[22]&IN2[36];
  assign P59[15] = IN1[22]&IN2[37];
  assign P60[14] = IN1[22]&IN2[38];
  assign P61[13] = IN1[22]&IN2[39];
  assign P62[12] = IN1[22]&IN2[40];
  assign P63[11] = IN1[22]&IN2[41];
  assign P64[10] = IN1[22]&IN2[42];
  assign P65[9] = IN1[22]&IN2[43];
  assign P66[8] = IN1[22]&IN2[44];
  assign P67[7] = IN1[22]&IN2[45];
  assign P68[6] = IN1[22]&IN2[46];
  assign P69[5] = IN1[22]&IN2[47];
  assign P70[4] = IN1[22]&IN2[48];
  assign P71[3] = IN1[22]&IN2[49];
  assign P72[2] = IN1[22]&IN2[50];
  assign P73[1] = IN1[22]&IN2[51];
  assign P74[0] = IN1[22]&IN2[52];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[23] = IN1[23]&IN2[12];
  assign P36[23] = IN1[23]&IN2[13];
  assign P37[23] = IN1[23]&IN2[14];
  assign P38[23] = IN1[23]&IN2[15];
  assign P39[23] = IN1[23]&IN2[16];
  assign P40[23] = IN1[23]&IN2[17];
  assign P41[23] = IN1[23]&IN2[18];
  assign P42[23] = IN1[23]&IN2[19];
  assign P43[23] = IN1[23]&IN2[20];
  assign P44[23] = IN1[23]&IN2[21];
  assign P45[23] = IN1[23]&IN2[22];
  assign P46[23] = IN1[23]&IN2[23];
  assign P47[23] = IN1[23]&IN2[24];
  assign P48[23] = IN1[23]&IN2[25];
  assign P49[23] = IN1[23]&IN2[26];
  assign P50[23] = IN1[23]&IN2[27];
  assign P51[23] = IN1[23]&IN2[28];
  assign P52[23] = IN1[23]&IN2[29];
  assign P53[22] = IN1[23]&IN2[30];
  assign P54[21] = IN1[23]&IN2[31];
  assign P55[20] = IN1[23]&IN2[32];
  assign P56[19] = IN1[23]&IN2[33];
  assign P57[18] = IN1[23]&IN2[34];
  assign P58[17] = IN1[23]&IN2[35];
  assign P59[16] = IN1[23]&IN2[36];
  assign P60[15] = IN1[23]&IN2[37];
  assign P61[14] = IN1[23]&IN2[38];
  assign P62[13] = IN1[23]&IN2[39];
  assign P63[12] = IN1[23]&IN2[40];
  assign P64[11] = IN1[23]&IN2[41];
  assign P65[10] = IN1[23]&IN2[42];
  assign P66[9] = IN1[23]&IN2[43];
  assign P67[8] = IN1[23]&IN2[44];
  assign P68[7] = IN1[23]&IN2[45];
  assign P69[6] = IN1[23]&IN2[46];
  assign P70[5] = IN1[23]&IN2[47];
  assign P71[4] = IN1[23]&IN2[48];
  assign P72[3] = IN1[23]&IN2[49];
  assign P73[2] = IN1[23]&IN2[50];
  assign P74[1] = IN1[23]&IN2[51];
  assign P75[0] = IN1[23]&IN2[52];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[24] = IN1[24]&IN2[11];
  assign P36[24] = IN1[24]&IN2[12];
  assign P37[24] = IN1[24]&IN2[13];
  assign P38[24] = IN1[24]&IN2[14];
  assign P39[24] = IN1[24]&IN2[15];
  assign P40[24] = IN1[24]&IN2[16];
  assign P41[24] = IN1[24]&IN2[17];
  assign P42[24] = IN1[24]&IN2[18];
  assign P43[24] = IN1[24]&IN2[19];
  assign P44[24] = IN1[24]&IN2[20];
  assign P45[24] = IN1[24]&IN2[21];
  assign P46[24] = IN1[24]&IN2[22];
  assign P47[24] = IN1[24]&IN2[23];
  assign P48[24] = IN1[24]&IN2[24];
  assign P49[24] = IN1[24]&IN2[25];
  assign P50[24] = IN1[24]&IN2[26];
  assign P51[24] = IN1[24]&IN2[27];
  assign P52[24] = IN1[24]&IN2[28];
  assign P53[23] = IN1[24]&IN2[29];
  assign P54[22] = IN1[24]&IN2[30];
  assign P55[21] = IN1[24]&IN2[31];
  assign P56[20] = IN1[24]&IN2[32];
  assign P57[19] = IN1[24]&IN2[33];
  assign P58[18] = IN1[24]&IN2[34];
  assign P59[17] = IN1[24]&IN2[35];
  assign P60[16] = IN1[24]&IN2[36];
  assign P61[15] = IN1[24]&IN2[37];
  assign P62[14] = IN1[24]&IN2[38];
  assign P63[13] = IN1[24]&IN2[39];
  assign P64[12] = IN1[24]&IN2[40];
  assign P65[11] = IN1[24]&IN2[41];
  assign P66[10] = IN1[24]&IN2[42];
  assign P67[9] = IN1[24]&IN2[43];
  assign P68[8] = IN1[24]&IN2[44];
  assign P69[7] = IN1[24]&IN2[45];
  assign P70[6] = IN1[24]&IN2[46];
  assign P71[5] = IN1[24]&IN2[47];
  assign P72[4] = IN1[24]&IN2[48];
  assign P73[3] = IN1[24]&IN2[49];
  assign P74[2] = IN1[24]&IN2[50];
  assign P75[1] = IN1[24]&IN2[51];
  assign P76[0] = IN1[24]&IN2[52];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[25] = IN1[25]&IN2[10];
  assign P36[25] = IN1[25]&IN2[11];
  assign P37[25] = IN1[25]&IN2[12];
  assign P38[25] = IN1[25]&IN2[13];
  assign P39[25] = IN1[25]&IN2[14];
  assign P40[25] = IN1[25]&IN2[15];
  assign P41[25] = IN1[25]&IN2[16];
  assign P42[25] = IN1[25]&IN2[17];
  assign P43[25] = IN1[25]&IN2[18];
  assign P44[25] = IN1[25]&IN2[19];
  assign P45[25] = IN1[25]&IN2[20];
  assign P46[25] = IN1[25]&IN2[21];
  assign P47[25] = IN1[25]&IN2[22];
  assign P48[25] = IN1[25]&IN2[23];
  assign P49[25] = IN1[25]&IN2[24];
  assign P50[25] = IN1[25]&IN2[25];
  assign P51[25] = IN1[25]&IN2[26];
  assign P52[25] = IN1[25]&IN2[27];
  assign P53[24] = IN1[25]&IN2[28];
  assign P54[23] = IN1[25]&IN2[29];
  assign P55[22] = IN1[25]&IN2[30];
  assign P56[21] = IN1[25]&IN2[31];
  assign P57[20] = IN1[25]&IN2[32];
  assign P58[19] = IN1[25]&IN2[33];
  assign P59[18] = IN1[25]&IN2[34];
  assign P60[17] = IN1[25]&IN2[35];
  assign P61[16] = IN1[25]&IN2[36];
  assign P62[15] = IN1[25]&IN2[37];
  assign P63[14] = IN1[25]&IN2[38];
  assign P64[13] = IN1[25]&IN2[39];
  assign P65[12] = IN1[25]&IN2[40];
  assign P66[11] = IN1[25]&IN2[41];
  assign P67[10] = IN1[25]&IN2[42];
  assign P68[9] = IN1[25]&IN2[43];
  assign P69[8] = IN1[25]&IN2[44];
  assign P70[7] = IN1[25]&IN2[45];
  assign P71[6] = IN1[25]&IN2[46];
  assign P72[5] = IN1[25]&IN2[47];
  assign P73[4] = IN1[25]&IN2[48];
  assign P74[3] = IN1[25]&IN2[49];
  assign P75[2] = IN1[25]&IN2[50];
  assign P76[1] = IN1[25]&IN2[51];
  assign P77[0] = IN1[25]&IN2[52];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[26] = IN1[26]&IN2[3];
  assign P30[26] = IN1[26]&IN2[4];
  assign P31[26] = IN1[26]&IN2[5];
  assign P32[26] = IN1[26]&IN2[6];
  assign P33[26] = IN1[26]&IN2[7];
  assign P34[26] = IN1[26]&IN2[8];
  assign P35[26] = IN1[26]&IN2[9];
  assign P36[26] = IN1[26]&IN2[10];
  assign P37[26] = IN1[26]&IN2[11];
  assign P38[26] = IN1[26]&IN2[12];
  assign P39[26] = IN1[26]&IN2[13];
  assign P40[26] = IN1[26]&IN2[14];
  assign P41[26] = IN1[26]&IN2[15];
  assign P42[26] = IN1[26]&IN2[16];
  assign P43[26] = IN1[26]&IN2[17];
  assign P44[26] = IN1[26]&IN2[18];
  assign P45[26] = IN1[26]&IN2[19];
  assign P46[26] = IN1[26]&IN2[20];
  assign P47[26] = IN1[26]&IN2[21];
  assign P48[26] = IN1[26]&IN2[22];
  assign P49[26] = IN1[26]&IN2[23];
  assign P50[26] = IN1[26]&IN2[24];
  assign P51[26] = IN1[26]&IN2[25];
  assign P52[26] = IN1[26]&IN2[26];
  assign P53[25] = IN1[26]&IN2[27];
  assign P54[24] = IN1[26]&IN2[28];
  assign P55[23] = IN1[26]&IN2[29];
  assign P56[22] = IN1[26]&IN2[30];
  assign P57[21] = IN1[26]&IN2[31];
  assign P58[20] = IN1[26]&IN2[32];
  assign P59[19] = IN1[26]&IN2[33];
  assign P60[18] = IN1[26]&IN2[34];
  assign P61[17] = IN1[26]&IN2[35];
  assign P62[16] = IN1[26]&IN2[36];
  assign P63[15] = IN1[26]&IN2[37];
  assign P64[14] = IN1[26]&IN2[38];
  assign P65[13] = IN1[26]&IN2[39];
  assign P66[12] = IN1[26]&IN2[40];
  assign P67[11] = IN1[26]&IN2[41];
  assign P68[10] = IN1[26]&IN2[42];
  assign P69[9] = IN1[26]&IN2[43];
  assign P70[8] = IN1[26]&IN2[44];
  assign P71[7] = IN1[26]&IN2[45];
  assign P72[6] = IN1[26]&IN2[46];
  assign P73[5] = IN1[26]&IN2[47];
  assign P74[4] = IN1[26]&IN2[48];
  assign P75[3] = IN1[26]&IN2[49];
  assign P76[2] = IN1[26]&IN2[50];
  assign P77[1] = IN1[26]&IN2[51];
  assign P78[0] = IN1[26]&IN2[52];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[27] = IN1[27]&IN2[2];
  assign P30[27] = IN1[27]&IN2[3];
  assign P31[27] = IN1[27]&IN2[4];
  assign P32[27] = IN1[27]&IN2[5];
  assign P33[27] = IN1[27]&IN2[6];
  assign P34[27] = IN1[27]&IN2[7];
  assign P35[27] = IN1[27]&IN2[8];
  assign P36[27] = IN1[27]&IN2[9];
  assign P37[27] = IN1[27]&IN2[10];
  assign P38[27] = IN1[27]&IN2[11];
  assign P39[27] = IN1[27]&IN2[12];
  assign P40[27] = IN1[27]&IN2[13];
  assign P41[27] = IN1[27]&IN2[14];
  assign P42[27] = IN1[27]&IN2[15];
  assign P43[27] = IN1[27]&IN2[16];
  assign P44[27] = IN1[27]&IN2[17];
  assign P45[27] = IN1[27]&IN2[18];
  assign P46[27] = IN1[27]&IN2[19];
  assign P47[27] = IN1[27]&IN2[20];
  assign P48[27] = IN1[27]&IN2[21];
  assign P49[27] = IN1[27]&IN2[22];
  assign P50[27] = IN1[27]&IN2[23];
  assign P51[27] = IN1[27]&IN2[24];
  assign P52[27] = IN1[27]&IN2[25];
  assign P53[26] = IN1[27]&IN2[26];
  assign P54[25] = IN1[27]&IN2[27];
  assign P55[24] = IN1[27]&IN2[28];
  assign P56[23] = IN1[27]&IN2[29];
  assign P57[22] = IN1[27]&IN2[30];
  assign P58[21] = IN1[27]&IN2[31];
  assign P59[20] = IN1[27]&IN2[32];
  assign P60[19] = IN1[27]&IN2[33];
  assign P61[18] = IN1[27]&IN2[34];
  assign P62[17] = IN1[27]&IN2[35];
  assign P63[16] = IN1[27]&IN2[36];
  assign P64[15] = IN1[27]&IN2[37];
  assign P65[14] = IN1[27]&IN2[38];
  assign P66[13] = IN1[27]&IN2[39];
  assign P67[12] = IN1[27]&IN2[40];
  assign P68[11] = IN1[27]&IN2[41];
  assign P69[10] = IN1[27]&IN2[42];
  assign P70[9] = IN1[27]&IN2[43];
  assign P71[8] = IN1[27]&IN2[44];
  assign P72[7] = IN1[27]&IN2[45];
  assign P73[6] = IN1[27]&IN2[46];
  assign P74[5] = IN1[27]&IN2[47];
  assign P75[4] = IN1[27]&IN2[48];
  assign P76[3] = IN1[27]&IN2[49];
  assign P77[2] = IN1[27]&IN2[50];
  assign P78[1] = IN1[27]&IN2[51];
  assign P79[0] = IN1[27]&IN2[52];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[28] = IN1[28]&IN2[1];
  assign P30[28] = IN1[28]&IN2[2];
  assign P31[28] = IN1[28]&IN2[3];
  assign P32[28] = IN1[28]&IN2[4];
  assign P33[28] = IN1[28]&IN2[5];
  assign P34[28] = IN1[28]&IN2[6];
  assign P35[28] = IN1[28]&IN2[7];
  assign P36[28] = IN1[28]&IN2[8];
  assign P37[28] = IN1[28]&IN2[9];
  assign P38[28] = IN1[28]&IN2[10];
  assign P39[28] = IN1[28]&IN2[11];
  assign P40[28] = IN1[28]&IN2[12];
  assign P41[28] = IN1[28]&IN2[13];
  assign P42[28] = IN1[28]&IN2[14];
  assign P43[28] = IN1[28]&IN2[15];
  assign P44[28] = IN1[28]&IN2[16];
  assign P45[28] = IN1[28]&IN2[17];
  assign P46[28] = IN1[28]&IN2[18];
  assign P47[28] = IN1[28]&IN2[19];
  assign P48[28] = IN1[28]&IN2[20];
  assign P49[28] = IN1[28]&IN2[21];
  assign P50[28] = IN1[28]&IN2[22];
  assign P51[28] = IN1[28]&IN2[23];
  assign P52[28] = IN1[28]&IN2[24];
  assign P53[27] = IN1[28]&IN2[25];
  assign P54[26] = IN1[28]&IN2[26];
  assign P55[25] = IN1[28]&IN2[27];
  assign P56[24] = IN1[28]&IN2[28];
  assign P57[23] = IN1[28]&IN2[29];
  assign P58[22] = IN1[28]&IN2[30];
  assign P59[21] = IN1[28]&IN2[31];
  assign P60[20] = IN1[28]&IN2[32];
  assign P61[19] = IN1[28]&IN2[33];
  assign P62[18] = IN1[28]&IN2[34];
  assign P63[17] = IN1[28]&IN2[35];
  assign P64[16] = IN1[28]&IN2[36];
  assign P65[15] = IN1[28]&IN2[37];
  assign P66[14] = IN1[28]&IN2[38];
  assign P67[13] = IN1[28]&IN2[39];
  assign P68[12] = IN1[28]&IN2[40];
  assign P69[11] = IN1[28]&IN2[41];
  assign P70[10] = IN1[28]&IN2[42];
  assign P71[9] = IN1[28]&IN2[43];
  assign P72[8] = IN1[28]&IN2[44];
  assign P73[7] = IN1[28]&IN2[45];
  assign P74[6] = IN1[28]&IN2[46];
  assign P75[5] = IN1[28]&IN2[47];
  assign P76[4] = IN1[28]&IN2[48];
  assign P77[3] = IN1[28]&IN2[49];
  assign P78[2] = IN1[28]&IN2[50];
  assign P79[1] = IN1[28]&IN2[51];
  assign P80[0] = IN1[28]&IN2[52];
  assign P29[29] = IN1[29]&IN2[0];
  assign P30[29] = IN1[29]&IN2[1];
  assign P31[29] = IN1[29]&IN2[2];
  assign P32[29] = IN1[29]&IN2[3];
  assign P33[29] = IN1[29]&IN2[4];
  assign P34[29] = IN1[29]&IN2[5];
  assign P35[29] = IN1[29]&IN2[6];
  assign P36[29] = IN1[29]&IN2[7];
  assign P37[29] = IN1[29]&IN2[8];
  assign P38[29] = IN1[29]&IN2[9];
  assign P39[29] = IN1[29]&IN2[10];
  assign P40[29] = IN1[29]&IN2[11];
  assign P41[29] = IN1[29]&IN2[12];
  assign P42[29] = IN1[29]&IN2[13];
  assign P43[29] = IN1[29]&IN2[14];
  assign P44[29] = IN1[29]&IN2[15];
  assign P45[29] = IN1[29]&IN2[16];
  assign P46[29] = IN1[29]&IN2[17];
  assign P47[29] = IN1[29]&IN2[18];
  assign P48[29] = IN1[29]&IN2[19];
  assign P49[29] = IN1[29]&IN2[20];
  assign P50[29] = IN1[29]&IN2[21];
  assign P51[29] = IN1[29]&IN2[22];
  assign P52[29] = IN1[29]&IN2[23];
  assign P53[28] = IN1[29]&IN2[24];
  assign P54[27] = IN1[29]&IN2[25];
  assign P55[26] = IN1[29]&IN2[26];
  assign P56[25] = IN1[29]&IN2[27];
  assign P57[24] = IN1[29]&IN2[28];
  assign P58[23] = IN1[29]&IN2[29];
  assign P59[22] = IN1[29]&IN2[30];
  assign P60[21] = IN1[29]&IN2[31];
  assign P61[20] = IN1[29]&IN2[32];
  assign P62[19] = IN1[29]&IN2[33];
  assign P63[18] = IN1[29]&IN2[34];
  assign P64[17] = IN1[29]&IN2[35];
  assign P65[16] = IN1[29]&IN2[36];
  assign P66[15] = IN1[29]&IN2[37];
  assign P67[14] = IN1[29]&IN2[38];
  assign P68[13] = IN1[29]&IN2[39];
  assign P69[12] = IN1[29]&IN2[40];
  assign P70[11] = IN1[29]&IN2[41];
  assign P71[10] = IN1[29]&IN2[42];
  assign P72[9] = IN1[29]&IN2[43];
  assign P73[8] = IN1[29]&IN2[44];
  assign P74[7] = IN1[29]&IN2[45];
  assign P75[6] = IN1[29]&IN2[46];
  assign P76[5] = IN1[29]&IN2[47];
  assign P77[4] = IN1[29]&IN2[48];
  assign P78[3] = IN1[29]&IN2[49];
  assign P79[2] = IN1[29]&IN2[50];
  assign P80[1] = IN1[29]&IN2[51];
  assign P81[0] = IN1[29]&IN2[52];
  assign P30[30] = IN1[30]&IN2[0];
  assign P31[30] = IN1[30]&IN2[1];
  assign P32[30] = IN1[30]&IN2[2];
  assign P33[30] = IN1[30]&IN2[3];
  assign P34[30] = IN1[30]&IN2[4];
  assign P35[30] = IN1[30]&IN2[5];
  assign P36[30] = IN1[30]&IN2[6];
  assign P37[30] = IN1[30]&IN2[7];
  assign P38[30] = IN1[30]&IN2[8];
  assign P39[30] = IN1[30]&IN2[9];
  assign P40[30] = IN1[30]&IN2[10];
  assign P41[30] = IN1[30]&IN2[11];
  assign P42[30] = IN1[30]&IN2[12];
  assign P43[30] = IN1[30]&IN2[13];
  assign P44[30] = IN1[30]&IN2[14];
  assign P45[30] = IN1[30]&IN2[15];
  assign P46[30] = IN1[30]&IN2[16];
  assign P47[30] = IN1[30]&IN2[17];
  assign P48[30] = IN1[30]&IN2[18];
  assign P49[30] = IN1[30]&IN2[19];
  assign P50[30] = IN1[30]&IN2[20];
  assign P51[30] = IN1[30]&IN2[21];
  assign P52[30] = IN1[30]&IN2[22];
  assign P53[29] = IN1[30]&IN2[23];
  assign P54[28] = IN1[30]&IN2[24];
  assign P55[27] = IN1[30]&IN2[25];
  assign P56[26] = IN1[30]&IN2[26];
  assign P57[25] = IN1[30]&IN2[27];
  assign P58[24] = IN1[30]&IN2[28];
  assign P59[23] = IN1[30]&IN2[29];
  assign P60[22] = IN1[30]&IN2[30];
  assign P61[21] = IN1[30]&IN2[31];
  assign P62[20] = IN1[30]&IN2[32];
  assign P63[19] = IN1[30]&IN2[33];
  assign P64[18] = IN1[30]&IN2[34];
  assign P65[17] = IN1[30]&IN2[35];
  assign P66[16] = IN1[30]&IN2[36];
  assign P67[15] = IN1[30]&IN2[37];
  assign P68[14] = IN1[30]&IN2[38];
  assign P69[13] = IN1[30]&IN2[39];
  assign P70[12] = IN1[30]&IN2[40];
  assign P71[11] = IN1[30]&IN2[41];
  assign P72[10] = IN1[30]&IN2[42];
  assign P73[9] = IN1[30]&IN2[43];
  assign P74[8] = IN1[30]&IN2[44];
  assign P75[7] = IN1[30]&IN2[45];
  assign P76[6] = IN1[30]&IN2[46];
  assign P77[5] = IN1[30]&IN2[47];
  assign P78[4] = IN1[30]&IN2[48];
  assign P79[3] = IN1[30]&IN2[49];
  assign P80[2] = IN1[30]&IN2[50];
  assign P81[1] = IN1[30]&IN2[51];
  assign P82[0] = IN1[30]&IN2[52];
  assign P31[31] = IN1[31]&IN2[0];
  assign P32[31] = IN1[31]&IN2[1];
  assign P33[31] = IN1[31]&IN2[2];
  assign P34[31] = IN1[31]&IN2[3];
  assign P35[31] = IN1[31]&IN2[4];
  assign P36[31] = IN1[31]&IN2[5];
  assign P37[31] = IN1[31]&IN2[6];
  assign P38[31] = IN1[31]&IN2[7];
  assign P39[31] = IN1[31]&IN2[8];
  assign P40[31] = IN1[31]&IN2[9];
  assign P41[31] = IN1[31]&IN2[10];
  assign P42[31] = IN1[31]&IN2[11];
  assign P43[31] = IN1[31]&IN2[12];
  assign P44[31] = IN1[31]&IN2[13];
  assign P45[31] = IN1[31]&IN2[14];
  assign P46[31] = IN1[31]&IN2[15];
  assign P47[31] = IN1[31]&IN2[16];
  assign P48[31] = IN1[31]&IN2[17];
  assign P49[31] = IN1[31]&IN2[18];
  assign P50[31] = IN1[31]&IN2[19];
  assign P51[31] = IN1[31]&IN2[20];
  assign P52[31] = IN1[31]&IN2[21];
  assign P53[30] = IN1[31]&IN2[22];
  assign P54[29] = IN1[31]&IN2[23];
  assign P55[28] = IN1[31]&IN2[24];
  assign P56[27] = IN1[31]&IN2[25];
  assign P57[26] = IN1[31]&IN2[26];
  assign P58[25] = IN1[31]&IN2[27];
  assign P59[24] = IN1[31]&IN2[28];
  assign P60[23] = IN1[31]&IN2[29];
  assign P61[22] = IN1[31]&IN2[30];
  assign P62[21] = IN1[31]&IN2[31];
  assign P63[20] = IN1[31]&IN2[32];
  assign P64[19] = IN1[31]&IN2[33];
  assign P65[18] = IN1[31]&IN2[34];
  assign P66[17] = IN1[31]&IN2[35];
  assign P67[16] = IN1[31]&IN2[36];
  assign P68[15] = IN1[31]&IN2[37];
  assign P69[14] = IN1[31]&IN2[38];
  assign P70[13] = IN1[31]&IN2[39];
  assign P71[12] = IN1[31]&IN2[40];
  assign P72[11] = IN1[31]&IN2[41];
  assign P73[10] = IN1[31]&IN2[42];
  assign P74[9] = IN1[31]&IN2[43];
  assign P75[8] = IN1[31]&IN2[44];
  assign P76[7] = IN1[31]&IN2[45];
  assign P77[6] = IN1[31]&IN2[46];
  assign P78[5] = IN1[31]&IN2[47];
  assign P79[4] = IN1[31]&IN2[48];
  assign P80[3] = IN1[31]&IN2[49];
  assign P81[2] = IN1[31]&IN2[50];
  assign P82[1] = IN1[31]&IN2[51];
  assign P83[0] = IN1[31]&IN2[52];
  assign P32[32] = IN1[32]&IN2[0];
  assign P33[32] = IN1[32]&IN2[1];
  assign P34[32] = IN1[32]&IN2[2];
  assign P35[32] = IN1[32]&IN2[3];
  assign P36[32] = IN1[32]&IN2[4];
  assign P37[32] = IN1[32]&IN2[5];
  assign P38[32] = IN1[32]&IN2[6];
  assign P39[32] = IN1[32]&IN2[7];
  assign P40[32] = IN1[32]&IN2[8];
  assign P41[32] = IN1[32]&IN2[9];
  assign P42[32] = IN1[32]&IN2[10];
  assign P43[32] = IN1[32]&IN2[11];
  assign P44[32] = IN1[32]&IN2[12];
  assign P45[32] = IN1[32]&IN2[13];
  assign P46[32] = IN1[32]&IN2[14];
  assign P47[32] = IN1[32]&IN2[15];
  assign P48[32] = IN1[32]&IN2[16];
  assign P49[32] = IN1[32]&IN2[17];
  assign P50[32] = IN1[32]&IN2[18];
  assign P51[32] = IN1[32]&IN2[19];
  assign P52[32] = IN1[32]&IN2[20];
  assign P53[31] = IN1[32]&IN2[21];
  assign P54[30] = IN1[32]&IN2[22];
  assign P55[29] = IN1[32]&IN2[23];
  assign P56[28] = IN1[32]&IN2[24];
  assign P57[27] = IN1[32]&IN2[25];
  assign P58[26] = IN1[32]&IN2[26];
  assign P59[25] = IN1[32]&IN2[27];
  assign P60[24] = IN1[32]&IN2[28];
  assign P61[23] = IN1[32]&IN2[29];
  assign P62[22] = IN1[32]&IN2[30];
  assign P63[21] = IN1[32]&IN2[31];
  assign P64[20] = IN1[32]&IN2[32];
  assign P65[19] = IN1[32]&IN2[33];
  assign P66[18] = IN1[32]&IN2[34];
  assign P67[17] = IN1[32]&IN2[35];
  assign P68[16] = IN1[32]&IN2[36];
  assign P69[15] = IN1[32]&IN2[37];
  assign P70[14] = IN1[32]&IN2[38];
  assign P71[13] = IN1[32]&IN2[39];
  assign P72[12] = IN1[32]&IN2[40];
  assign P73[11] = IN1[32]&IN2[41];
  assign P74[10] = IN1[32]&IN2[42];
  assign P75[9] = IN1[32]&IN2[43];
  assign P76[8] = IN1[32]&IN2[44];
  assign P77[7] = IN1[32]&IN2[45];
  assign P78[6] = IN1[32]&IN2[46];
  assign P79[5] = IN1[32]&IN2[47];
  assign P80[4] = IN1[32]&IN2[48];
  assign P81[3] = IN1[32]&IN2[49];
  assign P82[2] = IN1[32]&IN2[50];
  assign P83[1] = IN1[32]&IN2[51];
  assign P84[0] = IN1[32]&IN2[52];
  assign P33[33] = IN1[33]&IN2[0];
  assign P34[33] = IN1[33]&IN2[1];
  assign P35[33] = IN1[33]&IN2[2];
  assign P36[33] = IN1[33]&IN2[3];
  assign P37[33] = IN1[33]&IN2[4];
  assign P38[33] = IN1[33]&IN2[5];
  assign P39[33] = IN1[33]&IN2[6];
  assign P40[33] = IN1[33]&IN2[7];
  assign P41[33] = IN1[33]&IN2[8];
  assign P42[33] = IN1[33]&IN2[9];
  assign P43[33] = IN1[33]&IN2[10];
  assign P44[33] = IN1[33]&IN2[11];
  assign P45[33] = IN1[33]&IN2[12];
  assign P46[33] = IN1[33]&IN2[13];
  assign P47[33] = IN1[33]&IN2[14];
  assign P48[33] = IN1[33]&IN2[15];
  assign P49[33] = IN1[33]&IN2[16];
  assign P50[33] = IN1[33]&IN2[17];
  assign P51[33] = IN1[33]&IN2[18];
  assign P52[33] = IN1[33]&IN2[19];
  assign P53[32] = IN1[33]&IN2[20];
  assign P54[31] = IN1[33]&IN2[21];
  assign P55[30] = IN1[33]&IN2[22];
  assign P56[29] = IN1[33]&IN2[23];
  assign P57[28] = IN1[33]&IN2[24];
  assign P58[27] = IN1[33]&IN2[25];
  assign P59[26] = IN1[33]&IN2[26];
  assign P60[25] = IN1[33]&IN2[27];
  assign P61[24] = IN1[33]&IN2[28];
  assign P62[23] = IN1[33]&IN2[29];
  assign P63[22] = IN1[33]&IN2[30];
  assign P64[21] = IN1[33]&IN2[31];
  assign P65[20] = IN1[33]&IN2[32];
  assign P66[19] = IN1[33]&IN2[33];
  assign P67[18] = IN1[33]&IN2[34];
  assign P68[17] = IN1[33]&IN2[35];
  assign P69[16] = IN1[33]&IN2[36];
  assign P70[15] = IN1[33]&IN2[37];
  assign P71[14] = IN1[33]&IN2[38];
  assign P72[13] = IN1[33]&IN2[39];
  assign P73[12] = IN1[33]&IN2[40];
  assign P74[11] = IN1[33]&IN2[41];
  assign P75[10] = IN1[33]&IN2[42];
  assign P76[9] = IN1[33]&IN2[43];
  assign P77[8] = IN1[33]&IN2[44];
  assign P78[7] = IN1[33]&IN2[45];
  assign P79[6] = IN1[33]&IN2[46];
  assign P80[5] = IN1[33]&IN2[47];
  assign P81[4] = IN1[33]&IN2[48];
  assign P82[3] = IN1[33]&IN2[49];
  assign P83[2] = IN1[33]&IN2[50];
  assign P84[1] = IN1[33]&IN2[51];
  assign P85[0] = IN1[33]&IN2[52];
  assign P34[34] = IN1[34]&IN2[0];
  assign P35[34] = IN1[34]&IN2[1];
  assign P36[34] = IN1[34]&IN2[2];
  assign P37[34] = IN1[34]&IN2[3];
  assign P38[34] = IN1[34]&IN2[4];
  assign P39[34] = IN1[34]&IN2[5];
  assign P40[34] = IN1[34]&IN2[6];
  assign P41[34] = IN1[34]&IN2[7];
  assign P42[34] = IN1[34]&IN2[8];
  assign P43[34] = IN1[34]&IN2[9];
  assign P44[34] = IN1[34]&IN2[10];
  assign P45[34] = IN1[34]&IN2[11];
  assign P46[34] = IN1[34]&IN2[12];
  assign P47[34] = IN1[34]&IN2[13];
  assign P48[34] = IN1[34]&IN2[14];
  assign P49[34] = IN1[34]&IN2[15];
  assign P50[34] = IN1[34]&IN2[16];
  assign P51[34] = IN1[34]&IN2[17];
  assign P52[34] = IN1[34]&IN2[18];
  assign P53[33] = IN1[34]&IN2[19];
  assign P54[32] = IN1[34]&IN2[20];
  assign P55[31] = IN1[34]&IN2[21];
  assign P56[30] = IN1[34]&IN2[22];
  assign P57[29] = IN1[34]&IN2[23];
  assign P58[28] = IN1[34]&IN2[24];
  assign P59[27] = IN1[34]&IN2[25];
  assign P60[26] = IN1[34]&IN2[26];
  assign P61[25] = IN1[34]&IN2[27];
  assign P62[24] = IN1[34]&IN2[28];
  assign P63[23] = IN1[34]&IN2[29];
  assign P64[22] = IN1[34]&IN2[30];
  assign P65[21] = IN1[34]&IN2[31];
  assign P66[20] = IN1[34]&IN2[32];
  assign P67[19] = IN1[34]&IN2[33];
  assign P68[18] = IN1[34]&IN2[34];
  assign P69[17] = IN1[34]&IN2[35];
  assign P70[16] = IN1[34]&IN2[36];
  assign P71[15] = IN1[34]&IN2[37];
  assign P72[14] = IN1[34]&IN2[38];
  assign P73[13] = IN1[34]&IN2[39];
  assign P74[12] = IN1[34]&IN2[40];
  assign P75[11] = IN1[34]&IN2[41];
  assign P76[10] = IN1[34]&IN2[42];
  assign P77[9] = IN1[34]&IN2[43];
  assign P78[8] = IN1[34]&IN2[44];
  assign P79[7] = IN1[34]&IN2[45];
  assign P80[6] = IN1[34]&IN2[46];
  assign P81[5] = IN1[34]&IN2[47];
  assign P82[4] = IN1[34]&IN2[48];
  assign P83[3] = IN1[34]&IN2[49];
  assign P84[2] = IN1[34]&IN2[50];
  assign P85[1] = IN1[34]&IN2[51];
  assign P86[0] = IN1[34]&IN2[52];
  assign P35[35] = IN1[35]&IN2[0];
  assign P36[35] = IN1[35]&IN2[1];
  assign P37[35] = IN1[35]&IN2[2];
  assign P38[35] = IN1[35]&IN2[3];
  assign P39[35] = IN1[35]&IN2[4];
  assign P40[35] = IN1[35]&IN2[5];
  assign P41[35] = IN1[35]&IN2[6];
  assign P42[35] = IN1[35]&IN2[7];
  assign P43[35] = IN1[35]&IN2[8];
  assign P44[35] = IN1[35]&IN2[9];
  assign P45[35] = IN1[35]&IN2[10];
  assign P46[35] = IN1[35]&IN2[11];
  assign P47[35] = IN1[35]&IN2[12];
  assign P48[35] = IN1[35]&IN2[13];
  assign P49[35] = IN1[35]&IN2[14];
  assign P50[35] = IN1[35]&IN2[15];
  assign P51[35] = IN1[35]&IN2[16];
  assign P52[35] = IN1[35]&IN2[17];
  assign P53[34] = IN1[35]&IN2[18];
  assign P54[33] = IN1[35]&IN2[19];
  assign P55[32] = IN1[35]&IN2[20];
  assign P56[31] = IN1[35]&IN2[21];
  assign P57[30] = IN1[35]&IN2[22];
  assign P58[29] = IN1[35]&IN2[23];
  assign P59[28] = IN1[35]&IN2[24];
  assign P60[27] = IN1[35]&IN2[25];
  assign P61[26] = IN1[35]&IN2[26];
  assign P62[25] = IN1[35]&IN2[27];
  assign P63[24] = IN1[35]&IN2[28];
  assign P64[23] = IN1[35]&IN2[29];
  assign P65[22] = IN1[35]&IN2[30];
  assign P66[21] = IN1[35]&IN2[31];
  assign P67[20] = IN1[35]&IN2[32];
  assign P68[19] = IN1[35]&IN2[33];
  assign P69[18] = IN1[35]&IN2[34];
  assign P70[17] = IN1[35]&IN2[35];
  assign P71[16] = IN1[35]&IN2[36];
  assign P72[15] = IN1[35]&IN2[37];
  assign P73[14] = IN1[35]&IN2[38];
  assign P74[13] = IN1[35]&IN2[39];
  assign P75[12] = IN1[35]&IN2[40];
  assign P76[11] = IN1[35]&IN2[41];
  assign P77[10] = IN1[35]&IN2[42];
  assign P78[9] = IN1[35]&IN2[43];
  assign P79[8] = IN1[35]&IN2[44];
  assign P80[7] = IN1[35]&IN2[45];
  assign P81[6] = IN1[35]&IN2[46];
  assign P82[5] = IN1[35]&IN2[47];
  assign P83[4] = IN1[35]&IN2[48];
  assign P84[3] = IN1[35]&IN2[49];
  assign P85[2] = IN1[35]&IN2[50];
  assign P86[1] = IN1[35]&IN2[51];
  assign P87[0] = IN1[35]&IN2[52];
  assign P36[36] = IN1[36]&IN2[0];
  assign P37[36] = IN1[36]&IN2[1];
  assign P38[36] = IN1[36]&IN2[2];
  assign P39[36] = IN1[36]&IN2[3];
  assign P40[36] = IN1[36]&IN2[4];
  assign P41[36] = IN1[36]&IN2[5];
  assign P42[36] = IN1[36]&IN2[6];
  assign P43[36] = IN1[36]&IN2[7];
  assign P44[36] = IN1[36]&IN2[8];
  assign P45[36] = IN1[36]&IN2[9];
  assign P46[36] = IN1[36]&IN2[10];
  assign P47[36] = IN1[36]&IN2[11];
  assign P48[36] = IN1[36]&IN2[12];
  assign P49[36] = IN1[36]&IN2[13];
  assign P50[36] = IN1[36]&IN2[14];
  assign P51[36] = IN1[36]&IN2[15];
  assign P52[36] = IN1[36]&IN2[16];
  assign P53[35] = IN1[36]&IN2[17];
  assign P54[34] = IN1[36]&IN2[18];
  assign P55[33] = IN1[36]&IN2[19];
  assign P56[32] = IN1[36]&IN2[20];
  assign P57[31] = IN1[36]&IN2[21];
  assign P58[30] = IN1[36]&IN2[22];
  assign P59[29] = IN1[36]&IN2[23];
  assign P60[28] = IN1[36]&IN2[24];
  assign P61[27] = IN1[36]&IN2[25];
  assign P62[26] = IN1[36]&IN2[26];
  assign P63[25] = IN1[36]&IN2[27];
  assign P64[24] = IN1[36]&IN2[28];
  assign P65[23] = IN1[36]&IN2[29];
  assign P66[22] = IN1[36]&IN2[30];
  assign P67[21] = IN1[36]&IN2[31];
  assign P68[20] = IN1[36]&IN2[32];
  assign P69[19] = IN1[36]&IN2[33];
  assign P70[18] = IN1[36]&IN2[34];
  assign P71[17] = IN1[36]&IN2[35];
  assign P72[16] = IN1[36]&IN2[36];
  assign P73[15] = IN1[36]&IN2[37];
  assign P74[14] = IN1[36]&IN2[38];
  assign P75[13] = IN1[36]&IN2[39];
  assign P76[12] = IN1[36]&IN2[40];
  assign P77[11] = IN1[36]&IN2[41];
  assign P78[10] = IN1[36]&IN2[42];
  assign P79[9] = IN1[36]&IN2[43];
  assign P80[8] = IN1[36]&IN2[44];
  assign P81[7] = IN1[36]&IN2[45];
  assign P82[6] = IN1[36]&IN2[46];
  assign P83[5] = IN1[36]&IN2[47];
  assign P84[4] = IN1[36]&IN2[48];
  assign P85[3] = IN1[36]&IN2[49];
  assign P86[2] = IN1[36]&IN2[50];
  assign P87[1] = IN1[36]&IN2[51];
  assign P88[0] = IN1[36]&IN2[52];
  assign P37[37] = IN1[37]&IN2[0];
  assign P38[37] = IN1[37]&IN2[1];
  assign P39[37] = IN1[37]&IN2[2];
  assign P40[37] = IN1[37]&IN2[3];
  assign P41[37] = IN1[37]&IN2[4];
  assign P42[37] = IN1[37]&IN2[5];
  assign P43[37] = IN1[37]&IN2[6];
  assign P44[37] = IN1[37]&IN2[7];
  assign P45[37] = IN1[37]&IN2[8];
  assign P46[37] = IN1[37]&IN2[9];
  assign P47[37] = IN1[37]&IN2[10];
  assign P48[37] = IN1[37]&IN2[11];
  assign P49[37] = IN1[37]&IN2[12];
  assign P50[37] = IN1[37]&IN2[13];
  assign P51[37] = IN1[37]&IN2[14];
  assign P52[37] = IN1[37]&IN2[15];
  assign P53[36] = IN1[37]&IN2[16];
  assign P54[35] = IN1[37]&IN2[17];
  assign P55[34] = IN1[37]&IN2[18];
  assign P56[33] = IN1[37]&IN2[19];
  assign P57[32] = IN1[37]&IN2[20];
  assign P58[31] = IN1[37]&IN2[21];
  assign P59[30] = IN1[37]&IN2[22];
  assign P60[29] = IN1[37]&IN2[23];
  assign P61[28] = IN1[37]&IN2[24];
  assign P62[27] = IN1[37]&IN2[25];
  assign P63[26] = IN1[37]&IN2[26];
  assign P64[25] = IN1[37]&IN2[27];
  assign P65[24] = IN1[37]&IN2[28];
  assign P66[23] = IN1[37]&IN2[29];
  assign P67[22] = IN1[37]&IN2[30];
  assign P68[21] = IN1[37]&IN2[31];
  assign P69[20] = IN1[37]&IN2[32];
  assign P70[19] = IN1[37]&IN2[33];
  assign P71[18] = IN1[37]&IN2[34];
  assign P72[17] = IN1[37]&IN2[35];
  assign P73[16] = IN1[37]&IN2[36];
  assign P74[15] = IN1[37]&IN2[37];
  assign P75[14] = IN1[37]&IN2[38];
  assign P76[13] = IN1[37]&IN2[39];
  assign P77[12] = IN1[37]&IN2[40];
  assign P78[11] = IN1[37]&IN2[41];
  assign P79[10] = IN1[37]&IN2[42];
  assign P80[9] = IN1[37]&IN2[43];
  assign P81[8] = IN1[37]&IN2[44];
  assign P82[7] = IN1[37]&IN2[45];
  assign P83[6] = IN1[37]&IN2[46];
  assign P84[5] = IN1[37]&IN2[47];
  assign P85[4] = IN1[37]&IN2[48];
  assign P86[3] = IN1[37]&IN2[49];
  assign P87[2] = IN1[37]&IN2[50];
  assign P88[1] = IN1[37]&IN2[51];
  assign P89[0] = IN1[37]&IN2[52];
  assign P38[38] = IN1[38]&IN2[0];
  assign P39[38] = IN1[38]&IN2[1];
  assign P40[38] = IN1[38]&IN2[2];
  assign P41[38] = IN1[38]&IN2[3];
  assign P42[38] = IN1[38]&IN2[4];
  assign P43[38] = IN1[38]&IN2[5];
  assign P44[38] = IN1[38]&IN2[6];
  assign P45[38] = IN1[38]&IN2[7];
  assign P46[38] = IN1[38]&IN2[8];
  assign P47[38] = IN1[38]&IN2[9];
  assign P48[38] = IN1[38]&IN2[10];
  assign P49[38] = IN1[38]&IN2[11];
  assign P50[38] = IN1[38]&IN2[12];
  assign P51[38] = IN1[38]&IN2[13];
  assign P52[38] = IN1[38]&IN2[14];
  assign P53[37] = IN1[38]&IN2[15];
  assign P54[36] = IN1[38]&IN2[16];
  assign P55[35] = IN1[38]&IN2[17];
  assign P56[34] = IN1[38]&IN2[18];
  assign P57[33] = IN1[38]&IN2[19];
  assign P58[32] = IN1[38]&IN2[20];
  assign P59[31] = IN1[38]&IN2[21];
  assign P60[30] = IN1[38]&IN2[22];
  assign P61[29] = IN1[38]&IN2[23];
  assign P62[28] = IN1[38]&IN2[24];
  assign P63[27] = IN1[38]&IN2[25];
  assign P64[26] = IN1[38]&IN2[26];
  assign P65[25] = IN1[38]&IN2[27];
  assign P66[24] = IN1[38]&IN2[28];
  assign P67[23] = IN1[38]&IN2[29];
  assign P68[22] = IN1[38]&IN2[30];
  assign P69[21] = IN1[38]&IN2[31];
  assign P70[20] = IN1[38]&IN2[32];
  assign P71[19] = IN1[38]&IN2[33];
  assign P72[18] = IN1[38]&IN2[34];
  assign P73[17] = IN1[38]&IN2[35];
  assign P74[16] = IN1[38]&IN2[36];
  assign P75[15] = IN1[38]&IN2[37];
  assign P76[14] = IN1[38]&IN2[38];
  assign P77[13] = IN1[38]&IN2[39];
  assign P78[12] = IN1[38]&IN2[40];
  assign P79[11] = IN1[38]&IN2[41];
  assign P80[10] = IN1[38]&IN2[42];
  assign P81[9] = IN1[38]&IN2[43];
  assign P82[8] = IN1[38]&IN2[44];
  assign P83[7] = IN1[38]&IN2[45];
  assign P84[6] = IN1[38]&IN2[46];
  assign P85[5] = IN1[38]&IN2[47];
  assign P86[4] = IN1[38]&IN2[48];
  assign P87[3] = IN1[38]&IN2[49];
  assign P88[2] = IN1[38]&IN2[50];
  assign P89[1] = IN1[38]&IN2[51];
  assign P90[0] = IN1[38]&IN2[52];
  assign P39[39] = IN1[39]&IN2[0];
  assign P40[39] = IN1[39]&IN2[1];
  assign P41[39] = IN1[39]&IN2[2];
  assign P42[39] = IN1[39]&IN2[3];
  assign P43[39] = IN1[39]&IN2[4];
  assign P44[39] = IN1[39]&IN2[5];
  assign P45[39] = IN1[39]&IN2[6];
  assign P46[39] = IN1[39]&IN2[7];
  assign P47[39] = IN1[39]&IN2[8];
  assign P48[39] = IN1[39]&IN2[9];
  assign P49[39] = IN1[39]&IN2[10];
  assign P50[39] = IN1[39]&IN2[11];
  assign P51[39] = IN1[39]&IN2[12];
  assign P52[39] = IN1[39]&IN2[13];
  assign P53[38] = IN1[39]&IN2[14];
  assign P54[37] = IN1[39]&IN2[15];
  assign P55[36] = IN1[39]&IN2[16];
  assign P56[35] = IN1[39]&IN2[17];
  assign P57[34] = IN1[39]&IN2[18];
  assign P58[33] = IN1[39]&IN2[19];
  assign P59[32] = IN1[39]&IN2[20];
  assign P60[31] = IN1[39]&IN2[21];
  assign P61[30] = IN1[39]&IN2[22];
  assign P62[29] = IN1[39]&IN2[23];
  assign P63[28] = IN1[39]&IN2[24];
  assign P64[27] = IN1[39]&IN2[25];
  assign P65[26] = IN1[39]&IN2[26];
  assign P66[25] = IN1[39]&IN2[27];
  assign P67[24] = IN1[39]&IN2[28];
  assign P68[23] = IN1[39]&IN2[29];
  assign P69[22] = IN1[39]&IN2[30];
  assign P70[21] = IN1[39]&IN2[31];
  assign P71[20] = IN1[39]&IN2[32];
  assign P72[19] = IN1[39]&IN2[33];
  assign P73[18] = IN1[39]&IN2[34];
  assign P74[17] = IN1[39]&IN2[35];
  assign P75[16] = IN1[39]&IN2[36];
  assign P76[15] = IN1[39]&IN2[37];
  assign P77[14] = IN1[39]&IN2[38];
  assign P78[13] = IN1[39]&IN2[39];
  assign P79[12] = IN1[39]&IN2[40];
  assign P80[11] = IN1[39]&IN2[41];
  assign P81[10] = IN1[39]&IN2[42];
  assign P82[9] = IN1[39]&IN2[43];
  assign P83[8] = IN1[39]&IN2[44];
  assign P84[7] = IN1[39]&IN2[45];
  assign P85[6] = IN1[39]&IN2[46];
  assign P86[5] = IN1[39]&IN2[47];
  assign P87[4] = IN1[39]&IN2[48];
  assign P88[3] = IN1[39]&IN2[49];
  assign P89[2] = IN1[39]&IN2[50];
  assign P90[1] = IN1[39]&IN2[51];
  assign P91[0] = IN1[39]&IN2[52];
  assign P40[40] = IN1[40]&IN2[0];
  assign P41[40] = IN1[40]&IN2[1];
  assign P42[40] = IN1[40]&IN2[2];
  assign P43[40] = IN1[40]&IN2[3];
  assign P44[40] = IN1[40]&IN2[4];
  assign P45[40] = IN1[40]&IN2[5];
  assign P46[40] = IN1[40]&IN2[6];
  assign P47[40] = IN1[40]&IN2[7];
  assign P48[40] = IN1[40]&IN2[8];
  assign P49[40] = IN1[40]&IN2[9];
  assign P50[40] = IN1[40]&IN2[10];
  assign P51[40] = IN1[40]&IN2[11];
  assign P52[40] = IN1[40]&IN2[12];
  assign P53[39] = IN1[40]&IN2[13];
  assign P54[38] = IN1[40]&IN2[14];
  assign P55[37] = IN1[40]&IN2[15];
  assign P56[36] = IN1[40]&IN2[16];
  assign P57[35] = IN1[40]&IN2[17];
  assign P58[34] = IN1[40]&IN2[18];
  assign P59[33] = IN1[40]&IN2[19];
  assign P60[32] = IN1[40]&IN2[20];
  assign P61[31] = IN1[40]&IN2[21];
  assign P62[30] = IN1[40]&IN2[22];
  assign P63[29] = IN1[40]&IN2[23];
  assign P64[28] = IN1[40]&IN2[24];
  assign P65[27] = IN1[40]&IN2[25];
  assign P66[26] = IN1[40]&IN2[26];
  assign P67[25] = IN1[40]&IN2[27];
  assign P68[24] = IN1[40]&IN2[28];
  assign P69[23] = IN1[40]&IN2[29];
  assign P70[22] = IN1[40]&IN2[30];
  assign P71[21] = IN1[40]&IN2[31];
  assign P72[20] = IN1[40]&IN2[32];
  assign P73[19] = IN1[40]&IN2[33];
  assign P74[18] = IN1[40]&IN2[34];
  assign P75[17] = IN1[40]&IN2[35];
  assign P76[16] = IN1[40]&IN2[36];
  assign P77[15] = IN1[40]&IN2[37];
  assign P78[14] = IN1[40]&IN2[38];
  assign P79[13] = IN1[40]&IN2[39];
  assign P80[12] = IN1[40]&IN2[40];
  assign P81[11] = IN1[40]&IN2[41];
  assign P82[10] = IN1[40]&IN2[42];
  assign P83[9] = IN1[40]&IN2[43];
  assign P84[8] = IN1[40]&IN2[44];
  assign P85[7] = IN1[40]&IN2[45];
  assign P86[6] = IN1[40]&IN2[46];
  assign P87[5] = IN1[40]&IN2[47];
  assign P88[4] = IN1[40]&IN2[48];
  assign P89[3] = IN1[40]&IN2[49];
  assign P90[2] = IN1[40]&IN2[50];
  assign P91[1] = IN1[40]&IN2[51];
  assign P92[0] = IN1[40]&IN2[52];
  assign P41[41] = IN1[41]&IN2[0];
  assign P42[41] = IN1[41]&IN2[1];
  assign P43[41] = IN1[41]&IN2[2];
  assign P44[41] = IN1[41]&IN2[3];
  assign P45[41] = IN1[41]&IN2[4];
  assign P46[41] = IN1[41]&IN2[5];
  assign P47[41] = IN1[41]&IN2[6];
  assign P48[41] = IN1[41]&IN2[7];
  assign P49[41] = IN1[41]&IN2[8];
  assign P50[41] = IN1[41]&IN2[9];
  assign P51[41] = IN1[41]&IN2[10];
  assign P52[41] = IN1[41]&IN2[11];
  assign P53[40] = IN1[41]&IN2[12];
  assign P54[39] = IN1[41]&IN2[13];
  assign P55[38] = IN1[41]&IN2[14];
  assign P56[37] = IN1[41]&IN2[15];
  assign P57[36] = IN1[41]&IN2[16];
  assign P58[35] = IN1[41]&IN2[17];
  assign P59[34] = IN1[41]&IN2[18];
  assign P60[33] = IN1[41]&IN2[19];
  assign P61[32] = IN1[41]&IN2[20];
  assign P62[31] = IN1[41]&IN2[21];
  assign P63[30] = IN1[41]&IN2[22];
  assign P64[29] = IN1[41]&IN2[23];
  assign P65[28] = IN1[41]&IN2[24];
  assign P66[27] = IN1[41]&IN2[25];
  assign P67[26] = IN1[41]&IN2[26];
  assign P68[25] = IN1[41]&IN2[27];
  assign P69[24] = IN1[41]&IN2[28];
  assign P70[23] = IN1[41]&IN2[29];
  assign P71[22] = IN1[41]&IN2[30];
  assign P72[21] = IN1[41]&IN2[31];
  assign P73[20] = IN1[41]&IN2[32];
  assign P74[19] = IN1[41]&IN2[33];
  assign P75[18] = IN1[41]&IN2[34];
  assign P76[17] = IN1[41]&IN2[35];
  assign P77[16] = IN1[41]&IN2[36];
  assign P78[15] = IN1[41]&IN2[37];
  assign P79[14] = IN1[41]&IN2[38];
  assign P80[13] = IN1[41]&IN2[39];
  assign P81[12] = IN1[41]&IN2[40];
  assign P82[11] = IN1[41]&IN2[41];
  assign P83[10] = IN1[41]&IN2[42];
  assign P84[9] = IN1[41]&IN2[43];
  assign P85[8] = IN1[41]&IN2[44];
  assign P86[7] = IN1[41]&IN2[45];
  assign P87[6] = IN1[41]&IN2[46];
  assign P88[5] = IN1[41]&IN2[47];
  assign P89[4] = IN1[41]&IN2[48];
  assign P90[3] = IN1[41]&IN2[49];
  assign P91[2] = IN1[41]&IN2[50];
  assign P92[1] = IN1[41]&IN2[51];
  assign P93[0] = IN1[41]&IN2[52];
  assign P42[42] = IN1[42]&IN2[0];
  assign P43[42] = IN1[42]&IN2[1];
  assign P44[42] = IN1[42]&IN2[2];
  assign P45[42] = IN1[42]&IN2[3];
  assign P46[42] = IN1[42]&IN2[4];
  assign P47[42] = IN1[42]&IN2[5];
  assign P48[42] = IN1[42]&IN2[6];
  assign P49[42] = IN1[42]&IN2[7];
  assign P50[42] = IN1[42]&IN2[8];
  assign P51[42] = IN1[42]&IN2[9];
  assign P52[42] = IN1[42]&IN2[10];
  assign P53[41] = IN1[42]&IN2[11];
  assign P54[40] = IN1[42]&IN2[12];
  assign P55[39] = IN1[42]&IN2[13];
  assign P56[38] = IN1[42]&IN2[14];
  assign P57[37] = IN1[42]&IN2[15];
  assign P58[36] = IN1[42]&IN2[16];
  assign P59[35] = IN1[42]&IN2[17];
  assign P60[34] = IN1[42]&IN2[18];
  assign P61[33] = IN1[42]&IN2[19];
  assign P62[32] = IN1[42]&IN2[20];
  assign P63[31] = IN1[42]&IN2[21];
  assign P64[30] = IN1[42]&IN2[22];
  assign P65[29] = IN1[42]&IN2[23];
  assign P66[28] = IN1[42]&IN2[24];
  assign P67[27] = IN1[42]&IN2[25];
  assign P68[26] = IN1[42]&IN2[26];
  assign P69[25] = IN1[42]&IN2[27];
  assign P70[24] = IN1[42]&IN2[28];
  assign P71[23] = IN1[42]&IN2[29];
  assign P72[22] = IN1[42]&IN2[30];
  assign P73[21] = IN1[42]&IN2[31];
  assign P74[20] = IN1[42]&IN2[32];
  assign P75[19] = IN1[42]&IN2[33];
  assign P76[18] = IN1[42]&IN2[34];
  assign P77[17] = IN1[42]&IN2[35];
  assign P78[16] = IN1[42]&IN2[36];
  assign P79[15] = IN1[42]&IN2[37];
  assign P80[14] = IN1[42]&IN2[38];
  assign P81[13] = IN1[42]&IN2[39];
  assign P82[12] = IN1[42]&IN2[40];
  assign P83[11] = IN1[42]&IN2[41];
  assign P84[10] = IN1[42]&IN2[42];
  assign P85[9] = IN1[42]&IN2[43];
  assign P86[8] = IN1[42]&IN2[44];
  assign P87[7] = IN1[42]&IN2[45];
  assign P88[6] = IN1[42]&IN2[46];
  assign P89[5] = IN1[42]&IN2[47];
  assign P90[4] = IN1[42]&IN2[48];
  assign P91[3] = IN1[42]&IN2[49];
  assign P92[2] = IN1[42]&IN2[50];
  assign P93[1] = IN1[42]&IN2[51];
  assign P94[0] = IN1[42]&IN2[52];
  assign P43[43] = IN1[43]&IN2[0];
  assign P44[43] = IN1[43]&IN2[1];
  assign P45[43] = IN1[43]&IN2[2];
  assign P46[43] = IN1[43]&IN2[3];
  assign P47[43] = IN1[43]&IN2[4];
  assign P48[43] = IN1[43]&IN2[5];
  assign P49[43] = IN1[43]&IN2[6];
  assign P50[43] = IN1[43]&IN2[7];
  assign P51[43] = IN1[43]&IN2[8];
  assign P52[43] = IN1[43]&IN2[9];
  assign P53[42] = IN1[43]&IN2[10];
  assign P54[41] = IN1[43]&IN2[11];
  assign P55[40] = IN1[43]&IN2[12];
  assign P56[39] = IN1[43]&IN2[13];
  assign P57[38] = IN1[43]&IN2[14];
  assign P58[37] = IN1[43]&IN2[15];
  assign P59[36] = IN1[43]&IN2[16];
  assign P60[35] = IN1[43]&IN2[17];
  assign P61[34] = IN1[43]&IN2[18];
  assign P62[33] = IN1[43]&IN2[19];
  assign P63[32] = IN1[43]&IN2[20];
  assign P64[31] = IN1[43]&IN2[21];
  assign P65[30] = IN1[43]&IN2[22];
  assign P66[29] = IN1[43]&IN2[23];
  assign P67[28] = IN1[43]&IN2[24];
  assign P68[27] = IN1[43]&IN2[25];
  assign P69[26] = IN1[43]&IN2[26];
  assign P70[25] = IN1[43]&IN2[27];
  assign P71[24] = IN1[43]&IN2[28];
  assign P72[23] = IN1[43]&IN2[29];
  assign P73[22] = IN1[43]&IN2[30];
  assign P74[21] = IN1[43]&IN2[31];
  assign P75[20] = IN1[43]&IN2[32];
  assign P76[19] = IN1[43]&IN2[33];
  assign P77[18] = IN1[43]&IN2[34];
  assign P78[17] = IN1[43]&IN2[35];
  assign P79[16] = IN1[43]&IN2[36];
  assign P80[15] = IN1[43]&IN2[37];
  assign P81[14] = IN1[43]&IN2[38];
  assign P82[13] = IN1[43]&IN2[39];
  assign P83[12] = IN1[43]&IN2[40];
  assign P84[11] = IN1[43]&IN2[41];
  assign P85[10] = IN1[43]&IN2[42];
  assign P86[9] = IN1[43]&IN2[43];
  assign P87[8] = IN1[43]&IN2[44];
  assign P88[7] = IN1[43]&IN2[45];
  assign P89[6] = IN1[43]&IN2[46];
  assign P90[5] = IN1[43]&IN2[47];
  assign P91[4] = IN1[43]&IN2[48];
  assign P92[3] = IN1[43]&IN2[49];
  assign P93[2] = IN1[43]&IN2[50];
  assign P94[1] = IN1[43]&IN2[51];
  assign P95[0] = IN1[43]&IN2[52];
  assign P44[44] = IN1[44]&IN2[0];
  assign P45[44] = IN1[44]&IN2[1];
  assign P46[44] = IN1[44]&IN2[2];
  assign P47[44] = IN1[44]&IN2[3];
  assign P48[44] = IN1[44]&IN2[4];
  assign P49[44] = IN1[44]&IN2[5];
  assign P50[44] = IN1[44]&IN2[6];
  assign P51[44] = IN1[44]&IN2[7];
  assign P52[44] = IN1[44]&IN2[8];
  assign P53[43] = IN1[44]&IN2[9];
  assign P54[42] = IN1[44]&IN2[10];
  assign P55[41] = IN1[44]&IN2[11];
  assign P56[40] = IN1[44]&IN2[12];
  assign P57[39] = IN1[44]&IN2[13];
  assign P58[38] = IN1[44]&IN2[14];
  assign P59[37] = IN1[44]&IN2[15];
  assign P60[36] = IN1[44]&IN2[16];
  assign P61[35] = IN1[44]&IN2[17];
  assign P62[34] = IN1[44]&IN2[18];
  assign P63[33] = IN1[44]&IN2[19];
  assign P64[32] = IN1[44]&IN2[20];
  assign P65[31] = IN1[44]&IN2[21];
  assign P66[30] = IN1[44]&IN2[22];
  assign P67[29] = IN1[44]&IN2[23];
  assign P68[28] = IN1[44]&IN2[24];
  assign P69[27] = IN1[44]&IN2[25];
  assign P70[26] = IN1[44]&IN2[26];
  assign P71[25] = IN1[44]&IN2[27];
  assign P72[24] = IN1[44]&IN2[28];
  assign P73[23] = IN1[44]&IN2[29];
  assign P74[22] = IN1[44]&IN2[30];
  assign P75[21] = IN1[44]&IN2[31];
  assign P76[20] = IN1[44]&IN2[32];
  assign P77[19] = IN1[44]&IN2[33];
  assign P78[18] = IN1[44]&IN2[34];
  assign P79[17] = IN1[44]&IN2[35];
  assign P80[16] = IN1[44]&IN2[36];
  assign P81[15] = IN1[44]&IN2[37];
  assign P82[14] = IN1[44]&IN2[38];
  assign P83[13] = IN1[44]&IN2[39];
  assign P84[12] = IN1[44]&IN2[40];
  assign P85[11] = IN1[44]&IN2[41];
  assign P86[10] = IN1[44]&IN2[42];
  assign P87[9] = IN1[44]&IN2[43];
  assign P88[8] = IN1[44]&IN2[44];
  assign P89[7] = IN1[44]&IN2[45];
  assign P90[6] = IN1[44]&IN2[46];
  assign P91[5] = IN1[44]&IN2[47];
  assign P92[4] = IN1[44]&IN2[48];
  assign P93[3] = IN1[44]&IN2[49];
  assign P94[2] = IN1[44]&IN2[50];
  assign P95[1] = IN1[44]&IN2[51];
  assign P96[0] = IN1[44]&IN2[52];
  assign P45[45] = IN1[45]&IN2[0];
  assign P46[45] = IN1[45]&IN2[1];
  assign P47[45] = IN1[45]&IN2[2];
  assign P48[45] = IN1[45]&IN2[3];
  assign P49[45] = IN1[45]&IN2[4];
  assign P50[45] = IN1[45]&IN2[5];
  assign P51[45] = IN1[45]&IN2[6];
  assign P52[45] = IN1[45]&IN2[7];
  assign P53[44] = IN1[45]&IN2[8];
  assign P54[43] = IN1[45]&IN2[9];
  assign P55[42] = IN1[45]&IN2[10];
  assign P56[41] = IN1[45]&IN2[11];
  assign P57[40] = IN1[45]&IN2[12];
  assign P58[39] = IN1[45]&IN2[13];
  assign P59[38] = IN1[45]&IN2[14];
  assign P60[37] = IN1[45]&IN2[15];
  assign P61[36] = IN1[45]&IN2[16];
  assign P62[35] = IN1[45]&IN2[17];
  assign P63[34] = IN1[45]&IN2[18];
  assign P64[33] = IN1[45]&IN2[19];
  assign P65[32] = IN1[45]&IN2[20];
  assign P66[31] = IN1[45]&IN2[21];
  assign P67[30] = IN1[45]&IN2[22];
  assign P68[29] = IN1[45]&IN2[23];
  assign P69[28] = IN1[45]&IN2[24];
  assign P70[27] = IN1[45]&IN2[25];
  assign P71[26] = IN1[45]&IN2[26];
  assign P72[25] = IN1[45]&IN2[27];
  assign P73[24] = IN1[45]&IN2[28];
  assign P74[23] = IN1[45]&IN2[29];
  assign P75[22] = IN1[45]&IN2[30];
  assign P76[21] = IN1[45]&IN2[31];
  assign P77[20] = IN1[45]&IN2[32];
  assign P78[19] = IN1[45]&IN2[33];
  assign P79[18] = IN1[45]&IN2[34];
  assign P80[17] = IN1[45]&IN2[35];
  assign P81[16] = IN1[45]&IN2[36];
  assign P82[15] = IN1[45]&IN2[37];
  assign P83[14] = IN1[45]&IN2[38];
  assign P84[13] = IN1[45]&IN2[39];
  assign P85[12] = IN1[45]&IN2[40];
  assign P86[11] = IN1[45]&IN2[41];
  assign P87[10] = IN1[45]&IN2[42];
  assign P88[9] = IN1[45]&IN2[43];
  assign P89[8] = IN1[45]&IN2[44];
  assign P90[7] = IN1[45]&IN2[45];
  assign P91[6] = IN1[45]&IN2[46];
  assign P92[5] = IN1[45]&IN2[47];
  assign P93[4] = IN1[45]&IN2[48];
  assign P94[3] = IN1[45]&IN2[49];
  assign P95[2] = IN1[45]&IN2[50];
  assign P96[1] = IN1[45]&IN2[51];
  assign P97[0] = IN1[45]&IN2[52];
  assign P46[46] = IN1[46]&IN2[0];
  assign P47[46] = IN1[46]&IN2[1];
  assign P48[46] = IN1[46]&IN2[2];
  assign P49[46] = IN1[46]&IN2[3];
  assign P50[46] = IN1[46]&IN2[4];
  assign P51[46] = IN1[46]&IN2[5];
  assign P52[46] = IN1[46]&IN2[6];
  assign P53[45] = IN1[46]&IN2[7];
  assign P54[44] = IN1[46]&IN2[8];
  assign P55[43] = IN1[46]&IN2[9];
  assign P56[42] = IN1[46]&IN2[10];
  assign P57[41] = IN1[46]&IN2[11];
  assign P58[40] = IN1[46]&IN2[12];
  assign P59[39] = IN1[46]&IN2[13];
  assign P60[38] = IN1[46]&IN2[14];
  assign P61[37] = IN1[46]&IN2[15];
  assign P62[36] = IN1[46]&IN2[16];
  assign P63[35] = IN1[46]&IN2[17];
  assign P64[34] = IN1[46]&IN2[18];
  assign P65[33] = IN1[46]&IN2[19];
  assign P66[32] = IN1[46]&IN2[20];
  assign P67[31] = IN1[46]&IN2[21];
  assign P68[30] = IN1[46]&IN2[22];
  assign P69[29] = IN1[46]&IN2[23];
  assign P70[28] = IN1[46]&IN2[24];
  assign P71[27] = IN1[46]&IN2[25];
  assign P72[26] = IN1[46]&IN2[26];
  assign P73[25] = IN1[46]&IN2[27];
  assign P74[24] = IN1[46]&IN2[28];
  assign P75[23] = IN1[46]&IN2[29];
  assign P76[22] = IN1[46]&IN2[30];
  assign P77[21] = IN1[46]&IN2[31];
  assign P78[20] = IN1[46]&IN2[32];
  assign P79[19] = IN1[46]&IN2[33];
  assign P80[18] = IN1[46]&IN2[34];
  assign P81[17] = IN1[46]&IN2[35];
  assign P82[16] = IN1[46]&IN2[36];
  assign P83[15] = IN1[46]&IN2[37];
  assign P84[14] = IN1[46]&IN2[38];
  assign P85[13] = IN1[46]&IN2[39];
  assign P86[12] = IN1[46]&IN2[40];
  assign P87[11] = IN1[46]&IN2[41];
  assign P88[10] = IN1[46]&IN2[42];
  assign P89[9] = IN1[46]&IN2[43];
  assign P90[8] = IN1[46]&IN2[44];
  assign P91[7] = IN1[46]&IN2[45];
  assign P92[6] = IN1[46]&IN2[46];
  assign P93[5] = IN1[46]&IN2[47];
  assign P94[4] = IN1[46]&IN2[48];
  assign P95[3] = IN1[46]&IN2[49];
  assign P96[2] = IN1[46]&IN2[50];
  assign P97[1] = IN1[46]&IN2[51];
  assign P98[0] = IN1[46]&IN2[52];
  assign P47[47] = IN1[47]&IN2[0];
  assign P48[47] = IN1[47]&IN2[1];
  assign P49[47] = IN1[47]&IN2[2];
  assign P50[47] = IN1[47]&IN2[3];
  assign P51[47] = IN1[47]&IN2[4];
  assign P52[47] = IN1[47]&IN2[5];
  assign P53[46] = IN1[47]&IN2[6];
  assign P54[45] = IN1[47]&IN2[7];
  assign P55[44] = IN1[47]&IN2[8];
  assign P56[43] = IN1[47]&IN2[9];
  assign P57[42] = IN1[47]&IN2[10];
  assign P58[41] = IN1[47]&IN2[11];
  assign P59[40] = IN1[47]&IN2[12];
  assign P60[39] = IN1[47]&IN2[13];
  assign P61[38] = IN1[47]&IN2[14];
  assign P62[37] = IN1[47]&IN2[15];
  assign P63[36] = IN1[47]&IN2[16];
  assign P64[35] = IN1[47]&IN2[17];
  assign P65[34] = IN1[47]&IN2[18];
  assign P66[33] = IN1[47]&IN2[19];
  assign P67[32] = IN1[47]&IN2[20];
  assign P68[31] = IN1[47]&IN2[21];
  assign P69[30] = IN1[47]&IN2[22];
  assign P70[29] = IN1[47]&IN2[23];
  assign P71[28] = IN1[47]&IN2[24];
  assign P72[27] = IN1[47]&IN2[25];
  assign P73[26] = IN1[47]&IN2[26];
  assign P74[25] = IN1[47]&IN2[27];
  assign P75[24] = IN1[47]&IN2[28];
  assign P76[23] = IN1[47]&IN2[29];
  assign P77[22] = IN1[47]&IN2[30];
  assign P78[21] = IN1[47]&IN2[31];
  assign P79[20] = IN1[47]&IN2[32];
  assign P80[19] = IN1[47]&IN2[33];
  assign P81[18] = IN1[47]&IN2[34];
  assign P82[17] = IN1[47]&IN2[35];
  assign P83[16] = IN1[47]&IN2[36];
  assign P84[15] = IN1[47]&IN2[37];
  assign P85[14] = IN1[47]&IN2[38];
  assign P86[13] = IN1[47]&IN2[39];
  assign P87[12] = IN1[47]&IN2[40];
  assign P88[11] = IN1[47]&IN2[41];
  assign P89[10] = IN1[47]&IN2[42];
  assign P90[9] = IN1[47]&IN2[43];
  assign P91[8] = IN1[47]&IN2[44];
  assign P92[7] = IN1[47]&IN2[45];
  assign P93[6] = IN1[47]&IN2[46];
  assign P94[5] = IN1[47]&IN2[47];
  assign P95[4] = IN1[47]&IN2[48];
  assign P96[3] = IN1[47]&IN2[49];
  assign P97[2] = IN1[47]&IN2[50];
  assign P98[1] = IN1[47]&IN2[51];
  assign P99[0] = IN1[47]&IN2[52];
  assign P48[48] = IN1[48]&IN2[0];
  assign P49[48] = IN1[48]&IN2[1];
  assign P50[48] = IN1[48]&IN2[2];
  assign P51[48] = IN1[48]&IN2[3];
  assign P52[48] = IN1[48]&IN2[4];
  assign P53[47] = IN1[48]&IN2[5];
  assign P54[46] = IN1[48]&IN2[6];
  assign P55[45] = IN1[48]&IN2[7];
  assign P56[44] = IN1[48]&IN2[8];
  assign P57[43] = IN1[48]&IN2[9];
  assign P58[42] = IN1[48]&IN2[10];
  assign P59[41] = IN1[48]&IN2[11];
  assign P60[40] = IN1[48]&IN2[12];
  assign P61[39] = IN1[48]&IN2[13];
  assign P62[38] = IN1[48]&IN2[14];
  assign P63[37] = IN1[48]&IN2[15];
  assign P64[36] = IN1[48]&IN2[16];
  assign P65[35] = IN1[48]&IN2[17];
  assign P66[34] = IN1[48]&IN2[18];
  assign P67[33] = IN1[48]&IN2[19];
  assign P68[32] = IN1[48]&IN2[20];
  assign P69[31] = IN1[48]&IN2[21];
  assign P70[30] = IN1[48]&IN2[22];
  assign P71[29] = IN1[48]&IN2[23];
  assign P72[28] = IN1[48]&IN2[24];
  assign P73[27] = IN1[48]&IN2[25];
  assign P74[26] = IN1[48]&IN2[26];
  assign P75[25] = IN1[48]&IN2[27];
  assign P76[24] = IN1[48]&IN2[28];
  assign P77[23] = IN1[48]&IN2[29];
  assign P78[22] = IN1[48]&IN2[30];
  assign P79[21] = IN1[48]&IN2[31];
  assign P80[20] = IN1[48]&IN2[32];
  assign P81[19] = IN1[48]&IN2[33];
  assign P82[18] = IN1[48]&IN2[34];
  assign P83[17] = IN1[48]&IN2[35];
  assign P84[16] = IN1[48]&IN2[36];
  assign P85[15] = IN1[48]&IN2[37];
  assign P86[14] = IN1[48]&IN2[38];
  assign P87[13] = IN1[48]&IN2[39];
  assign P88[12] = IN1[48]&IN2[40];
  assign P89[11] = IN1[48]&IN2[41];
  assign P90[10] = IN1[48]&IN2[42];
  assign P91[9] = IN1[48]&IN2[43];
  assign P92[8] = IN1[48]&IN2[44];
  assign P93[7] = IN1[48]&IN2[45];
  assign P94[6] = IN1[48]&IN2[46];
  assign P95[5] = IN1[48]&IN2[47];
  assign P96[4] = IN1[48]&IN2[48];
  assign P97[3] = IN1[48]&IN2[49];
  assign P98[2] = IN1[48]&IN2[50];
  assign P99[1] = IN1[48]&IN2[51];
  assign P100[0] = IN1[48]&IN2[52];
  assign P49[49] = IN1[49]&IN2[0];
  assign P50[49] = IN1[49]&IN2[1];
  assign P51[49] = IN1[49]&IN2[2];
  assign P52[49] = IN1[49]&IN2[3];
  assign P53[48] = IN1[49]&IN2[4];
  assign P54[47] = IN1[49]&IN2[5];
  assign P55[46] = IN1[49]&IN2[6];
  assign P56[45] = IN1[49]&IN2[7];
  assign P57[44] = IN1[49]&IN2[8];
  assign P58[43] = IN1[49]&IN2[9];
  assign P59[42] = IN1[49]&IN2[10];
  assign P60[41] = IN1[49]&IN2[11];
  assign P61[40] = IN1[49]&IN2[12];
  assign P62[39] = IN1[49]&IN2[13];
  assign P63[38] = IN1[49]&IN2[14];
  assign P64[37] = IN1[49]&IN2[15];
  assign P65[36] = IN1[49]&IN2[16];
  assign P66[35] = IN1[49]&IN2[17];
  assign P67[34] = IN1[49]&IN2[18];
  assign P68[33] = IN1[49]&IN2[19];
  assign P69[32] = IN1[49]&IN2[20];
  assign P70[31] = IN1[49]&IN2[21];
  assign P71[30] = IN1[49]&IN2[22];
  assign P72[29] = IN1[49]&IN2[23];
  assign P73[28] = IN1[49]&IN2[24];
  assign P74[27] = IN1[49]&IN2[25];
  assign P75[26] = IN1[49]&IN2[26];
  assign P76[25] = IN1[49]&IN2[27];
  assign P77[24] = IN1[49]&IN2[28];
  assign P78[23] = IN1[49]&IN2[29];
  assign P79[22] = IN1[49]&IN2[30];
  assign P80[21] = IN1[49]&IN2[31];
  assign P81[20] = IN1[49]&IN2[32];
  assign P82[19] = IN1[49]&IN2[33];
  assign P83[18] = IN1[49]&IN2[34];
  assign P84[17] = IN1[49]&IN2[35];
  assign P85[16] = IN1[49]&IN2[36];
  assign P86[15] = IN1[49]&IN2[37];
  assign P87[14] = IN1[49]&IN2[38];
  assign P88[13] = IN1[49]&IN2[39];
  assign P89[12] = IN1[49]&IN2[40];
  assign P90[11] = IN1[49]&IN2[41];
  assign P91[10] = IN1[49]&IN2[42];
  assign P92[9] = IN1[49]&IN2[43];
  assign P93[8] = IN1[49]&IN2[44];
  assign P94[7] = IN1[49]&IN2[45];
  assign P95[6] = IN1[49]&IN2[46];
  assign P96[5] = IN1[49]&IN2[47];
  assign P97[4] = IN1[49]&IN2[48];
  assign P98[3] = IN1[49]&IN2[49];
  assign P99[2] = IN1[49]&IN2[50];
  assign P100[1] = IN1[49]&IN2[51];
  assign P101[0] = IN1[49]&IN2[52];
  assign P50[50] = IN1[50]&IN2[0];
  assign P51[50] = IN1[50]&IN2[1];
  assign P52[50] = IN1[50]&IN2[2];
  assign P53[49] = IN1[50]&IN2[3];
  assign P54[48] = IN1[50]&IN2[4];
  assign P55[47] = IN1[50]&IN2[5];
  assign P56[46] = IN1[50]&IN2[6];
  assign P57[45] = IN1[50]&IN2[7];
  assign P58[44] = IN1[50]&IN2[8];
  assign P59[43] = IN1[50]&IN2[9];
  assign P60[42] = IN1[50]&IN2[10];
  assign P61[41] = IN1[50]&IN2[11];
  assign P62[40] = IN1[50]&IN2[12];
  assign P63[39] = IN1[50]&IN2[13];
  assign P64[38] = IN1[50]&IN2[14];
  assign P65[37] = IN1[50]&IN2[15];
  assign P66[36] = IN1[50]&IN2[16];
  assign P67[35] = IN1[50]&IN2[17];
  assign P68[34] = IN1[50]&IN2[18];
  assign P69[33] = IN1[50]&IN2[19];
  assign P70[32] = IN1[50]&IN2[20];
  assign P71[31] = IN1[50]&IN2[21];
  assign P72[30] = IN1[50]&IN2[22];
  assign P73[29] = IN1[50]&IN2[23];
  assign P74[28] = IN1[50]&IN2[24];
  assign P75[27] = IN1[50]&IN2[25];
  assign P76[26] = IN1[50]&IN2[26];
  assign P77[25] = IN1[50]&IN2[27];
  assign P78[24] = IN1[50]&IN2[28];
  assign P79[23] = IN1[50]&IN2[29];
  assign P80[22] = IN1[50]&IN2[30];
  assign P81[21] = IN1[50]&IN2[31];
  assign P82[20] = IN1[50]&IN2[32];
  assign P83[19] = IN1[50]&IN2[33];
  assign P84[18] = IN1[50]&IN2[34];
  assign P85[17] = IN1[50]&IN2[35];
  assign P86[16] = IN1[50]&IN2[36];
  assign P87[15] = IN1[50]&IN2[37];
  assign P88[14] = IN1[50]&IN2[38];
  assign P89[13] = IN1[50]&IN2[39];
  assign P90[12] = IN1[50]&IN2[40];
  assign P91[11] = IN1[50]&IN2[41];
  assign P92[10] = IN1[50]&IN2[42];
  assign P93[9] = IN1[50]&IN2[43];
  assign P94[8] = IN1[50]&IN2[44];
  assign P95[7] = IN1[50]&IN2[45];
  assign P96[6] = IN1[50]&IN2[46];
  assign P97[5] = IN1[50]&IN2[47];
  assign P98[4] = IN1[50]&IN2[48];
  assign P99[3] = IN1[50]&IN2[49];
  assign P100[2] = IN1[50]&IN2[50];
  assign P101[1] = IN1[50]&IN2[51];
  assign P102[0] = IN1[50]&IN2[52];
  assign P51[51] = IN1[51]&IN2[0];
  assign P52[51] = IN1[51]&IN2[1];
  assign P53[50] = IN1[51]&IN2[2];
  assign P54[49] = IN1[51]&IN2[3];
  assign P55[48] = IN1[51]&IN2[4];
  assign P56[47] = IN1[51]&IN2[5];
  assign P57[46] = IN1[51]&IN2[6];
  assign P58[45] = IN1[51]&IN2[7];
  assign P59[44] = IN1[51]&IN2[8];
  assign P60[43] = IN1[51]&IN2[9];
  assign P61[42] = IN1[51]&IN2[10];
  assign P62[41] = IN1[51]&IN2[11];
  assign P63[40] = IN1[51]&IN2[12];
  assign P64[39] = IN1[51]&IN2[13];
  assign P65[38] = IN1[51]&IN2[14];
  assign P66[37] = IN1[51]&IN2[15];
  assign P67[36] = IN1[51]&IN2[16];
  assign P68[35] = IN1[51]&IN2[17];
  assign P69[34] = IN1[51]&IN2[18];
  assign P70[33] = IN1[51]&IN2[19];
  assign P71[32] = IN1[51]&IN2[20];
  assign P72[31] = IN1[51]&IN2[21];
  assign P73[30] = IN1[51]&IN2[22];
  assign P74[29] = IN1[51]&IN2[23];
  assign P75[28] = IN1[51]&IN2[24];
  assign P76[27] = IN1[51]&IN2[25];
  assign P77[26] = IN1[51]&IN2[26];
  assign P78[25] = IN1[51]&IN2[27];
  assign P79[24] = IN1[51]&IN2[28];
  assign P80[23] = IN1[51]&IN2[29];
  assign P81[22] = IN1[51]&IN2[30];
  assign P82[21] = IN1[51]&IN2[31];
  assign P83[20] = IN1[51]&IN2[32];
  assign P84[19] = IN1[51]&IN2[33];
  assign P85[18] = IN1[51]&IN2[34];
  assign P86[17] = IN1[51]&IN2[35];
  assign P87[16] = IN1[51]&IN2[36];
  assign P88[15] = IN1[51]&IN2[37];
  assign P89[14] = IN1[51]&IN2[38];
  assign P90[13] = IN1[51]&IN2[39];
  assign P91[12] = IN1[51]&IN2[40];
  assign P92[11] = IN1[51]&IN2[41];
  assign P93[10] = IN1[51]&IN2[42];
  assign P94[9] = IN1[51]&IN2[43];
  assign P95[8] = IN1[51]&IN2[44];
  assign P96[7] = IN1[51]&IN2[45];
  assign P97[6] = IN1[51]&IN2[46];
  assign P98[5] = IN1[51]&IN2[47];
  assign P99[4] = IN1[51]&IN2[48];
  assign P100[3] = IN1[51]&IN2[49];
  assign P101[2] = IN1[51]&IN2[50];
  assign P102[1] = IN1[51]&IN2[51];
  assign P103[0] = IN1[51]&IN2[52];
  assign P52[52] = IN1[52]&IN2[0];
  assign P53[51] = IN1[52]&IN2[1];
  assign P54[50] = IN1[52]&IN2[2];
  assign P55[49] = IN1[52]&IN2[3];
  assign P56[48] = IN1[52]&IN2[4];
  assign P57[47] = IN1[52]&IN2[5];
  assign P58[46] = IN1[52]&IN2[6];
  assign P59[45] = IN1[52]&IN2[7];
  assign P60[44] = IN1[52]&IN2[8];
  assign P61[43] = IN1[52]&IN2[9];
  assign P62[42] = IN1[52]&IN2[10];
  assign P63[41] = IN1[52]&IN2[11];
  assign P64[40] = IN1[52]&IN2[12];
  assign P65[39] = IN1[52]&IN2[13];
  assign P66[38] = IN1[52]&IN2[14];
  assign P67[37] = IN1[52]&IN2[15];
  assign P68[36] = IN1[52]&IN2[16];
  assign P69[35] = IN1[52]&IN2[17];
  assign P70[34] = IN1[52]&IN2[18];
  assign P71[33] = IN1[52]&IN2[19];
  assign P72[32] = IN1[52]&IN2[20];
  assign P73[31] = IN1[52]&IN2[21];
  assign P74[30] = IN1[52]&IN2[22];
  assign P75[29] = IN1[52]&IN2[23];
  assign P76[28] = IN1[52]&IN2[24];
  assign P77[27] = IN1[52]&IN2[25];
  assign P78[26] = IN1[52]&IN2[26];
  assign P79[25] = IN1[52]&IN2[27];
  assign P80[24] = IN1[52]&IN2[28];
  assign P81[23] = IN1[52]&IN2[29];
  assign P82[22] = IN1[52]&IN2[30];
  assign P83[21] = IN1[52]&IN2[31];
  assign P84[20] = IN1[52]&IN2[32];
  assign P85[19] = IN1[52]&IN2[33];
  assign P86[18] = IN1[52]&IN2[34];
  assign P87[17] = IN1[52]&IN2[35];
  assign P88[16] = IN1[52]&IN2[36];
  assign P89[15] = IN1[52]&IN2[37];
  assign P90[14] = IN1[52]&IN2[38];
  assign P91[13] = IN1[52]&IN2[39];
  assign P92[12] = IN1[52]&IN2[40];
  assign P93[11] = IN1[52]&IN2[41];
  assign P94[10] = IN1[52]&IN2[42];
  assign P95[9] = IN1[52]&IN2[43];
  assign P96[8] = IN1[52]&IN2[44];
  assign P97[7] = IN1[52]&IN2[45];
  assign P98[6] = IN1[52]&IN2[46];
  assign P99[5] = IN1[52]&IN2[47];
  assign P100[4] = IN1[52]&IN2[48];
  assign P101[3] = IN1[52]&IN2[49];
  assign P102[2] = IN1[52]&IN2[50];
  assign P103[1] = IN1[52]&IN2[51];
  assign P104[0] = IN1[52]&IN2[52];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, IN79, IN80, IN81, IN82, IN83, IN84, IN85, IN86, IN87, IN88, IN89, IN90, IN91, IN92, IN93, IN94, IN95, IN96, IN97, IN98, IN99, IN100, IN101, IN102, IN103, IN104, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [29:0] IN29;
  input [30:0] IN30;
  input [31:0] IN31;
  input [32:0] IN32;
  input [33:0] IN33;
  input [34:0] IN34;
  input [35:0] IN35;
  input [36:0] IN36;
  input [37:0] IN37;
  input [38:0] IN38;
  input [39:0] IN39;
  input [40:0] IN40;
  input [41:0] IN41;
  input [42:0] IN42;
  input [43:0] IN43;
  input [44:0] IN44;
  input [45:0] IN45;
  input [46:0] IN46;
  input [47:0] IN47;
  input [48:0] IN48;
  input [49:0] IN49;
  input [50:0] IN50;
  input [51:0] IN51;
  input [52:0] IN52;
  input [51:0] IN53;
  input [50:0] IN54;
  input [49:0] IN55;
  input [48:0] IN56;
  input [47:0] IN57;
  input [46:0] IN58;
  input [45:0] IN59;
  input [44:0] IN60;
  input [43:0] IN61;
  input [42:0] IN62;
  input [41:0] IN63;
  input [40:0] IN64;
  input [39:0] IN65;
  input [38:0] IN66;
  input [37:0] IN67;
  input [36:0] IN68;
  input [35:0] IN69;
  input [34:0] IN70;
  input [33:0] IN71;
  input [32:0] IN72;
  input [31:0] IN73;
  input [30:0] IN74;
  input [29:0] IN75;
  input [28:0] IN76;
  input [27:0] IN77;
  input [26:0] IN78;
  input [25:0] IN79;
  input [24:0] IN80;
  input [23:0] IN81;
  input [22:0] IN82;
  input [21:0] IN83;
  input [20:0] IN84;
  input [19:0] IN85;
  input [18:0] IN86;
  input [17:0] IN87;
  input [16:0] IN88;
  input [15:0] IN89;
  input [14:0] IN90;
  input [13:0] IN91;
  input [12:0] IN92;
  input [11:0] IN93;
  input [10:0] IN94;
  input [9:0] IN95;
  input [8:0] IN96;
  input [7:0] IN97;
  input [6:0] IN98;
  input [5:0] IN99;
  input [4:0] IN100;
  input [3:0] IN101;
  input [2:0] IN102;
  input [1:0] IN103;
  input [0:0] IN104;
  output [104:0] Out1;
  output [51:0] Out2;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2854;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2860;
  wire w2861;
  wire w2862;
  wire w2863;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2885;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2896;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2934;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2950;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2979;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2985;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2990;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3014;
  wire w3015;
  wire w3016;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3040;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3084;
  wire w3085;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3094;
  wire w3095;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3130;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3254;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3262;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3272;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3285;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3327;
  wire w3328;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3334;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3362;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3366;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3385;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3414;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3443;
  wire w3444;
  wire w3445;
  wire w3446;
  wire w3447;
  wire w3448;
  wire w3449;
  wire w3450;
  wire w3451;
  wire w3452;
  wire w3453;
  wire w3454;
  wire w3455;
  wire w3456;
  wire w3457;
  wire w3458;
  wire w3459;
  wire w3460;
  wire w3461;
  wire w3462;
  wire w3463;
  wire w3464;
  wire w3465;
  wire w3466;
  wire w3467;
  wire w3468;
  wire w3469;
  wire w3470;
  wire w3471;
  wire w3472;
  wire w3473;
  wire w3474;
  wire w3475;
  wire w3476;
  wire w3477;
  wire w3478;
  wire w3479;
  wire w3480;
  wire w3481;
  wire w3482;
  wire w3483;
  wire w3484;
  wire w3485;
  wire w3486;
  wire w3487;
  wire w3488;
  wire w3489;
  wire w3490;
  wire w3491;
  wire w3492;
  wire w3493;
  wire w3494;
  wire w3495;
  wire w3496;
  wire w3497;
  wire w3498;
  wire w3499;
  wire w3500;
  wire w3501;
  wire w3502;
  wire w3503;
  wire w3504;
  wire w3505;
  wire w3506;
  wire w3507;
  wire w3508;
  wire w3509;
  wire w3510;
  wire w3511;
  wire w3512;
  wire w3513;
  wire w3514;
  wire w3515;
  wire w3516;
  wire w3517;
  wire w3518;
  wire w3519;
  wire w3520;
  wire w3521;
  wire w3522;
  wire w3523;
  wire w3524;
  wire w3525;
  wire w3526;
  wire w3527;
  wire w3528;
  wire w3529;
  wire w3530;
  wire w3531;
  wire w3532;
  wire w3533;
  wire w3534;
  wire w3535;
  wire w3536;
  wire w3538;
  wire w3539;
  wire w3540;
  wire w3541;
  wire w3542;
  wire w3543;
  wire w3544;
  wire w3545;
  wire w3546;
  wire w3547;
  wire w3548;
  wire w3549;
  wire w3550;
  wire w3551;
  wire w3552;
  wire w3553;
  wire w3554;
  wire w3555;
  wire w3556;
  wire w3557;
  wire w3558;
  wire w3559;
  wire w3560;
  wire w3561;
  wire w3562;
  wire w3563;
  wire w3564;
  wire w3565;
  wire w3566;
  wire w3567;
  wire w3568;
  wire w3569;
  wire w3570;
  wire w3571;
  wire w3572;
  wire w3573;
  wire w3574;
  wire w3575;
  wire w3576;
  wire w3577;
  wire w3578;
  wire w3579;
  wire w3580;
  wire w3581;
  wire w3582;
  wire w3583;
  wire w3584;
  wire w3585;
  wire w3586;
  wire w3587;
  wire w3588;
  wire w3589;
  wire w3590;
  wire w3591;
  wire w3592;
  wire w3593;
  wire w3594;
  wire w3595;
  wire w3596;
  wire w3597;
  wire w3598;
  wire w3599;
  wire w3600;
  wire w3601;
  wire w3602;
  wire w3603;
  wire w3604;
  wire w3605;
  wire w3606;
  wire w3607;
  wire w3608;
  wire w3609;
  wire w3610;
  wire w3611;
  wire w3612;
  wire w3613;
  wire w3614;
  wire w3615;
  wire w3616;
  wire w3617;
  wire w3618;
  wire w3619;
  wire w3620;
  wire w3621;
  wire w3622;
  wire w3623;
  wire w3624;
  wire w3625;
  wire w3626;
  wire w3627;
  wire w3628;
  wire w3629;
  wire w3630;
  wire w3631;
  wire w3632;
  wire w3633;
  wire w3634;
  wire w3635;
  wire w3636;
  wire w3637;
  wire w3638;
  wire w3639;
  wire w3640;
  wire w3642;
  wire w3643;
  wire w3644;
  wire w3645;
  wire w3646;
  wire w3647;
  wire w3648;
  wire w3649;
  wire w3650;
  wire w3651;
  wire w3652;
  wire w3653;
  wire w3654;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3662;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3685;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3734;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3742;
  wire w3743;
  wire w3744;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3762;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3768;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3785;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3814;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3836;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3862;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3882;
  wire w3883;
  wire w3884;
  wire w3885;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3894;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3930;
  wire w3931;
  wire w3932;
  wire w3933;
  wire w3934;
  wire w3935;
  wire w3936;
  wire w3937;
  wire w3938;
  wire w3939;
  wire w3940;
  wire w3941;
  wire w3942;
  wire w3943;
  wire w3944;
  wire w3945;
  wire w3946;
  wire w3947;
  wire w3948;
  wire w3949;
  wire w3950;
  wire w3951;
  wire w3952;
  wire w3954;
  wire w3955;
  wire w3956;
  wire w3957;
  wire w3958;
  wire w3959;
  wire w3960;
  wire w3961;
  wire w3962;
  wire w3963;
  wire w3964;
  wire w3965;
  wire w3966;
  wire w3967;
  wire w3968;
  wire w3969;
  wire w3970;
  wire w3971;
  wire w3972;
  wire w3973;
  wire w3974;
  wire w3975;
  wire w3976;
  wire w3977;
  wire w3978;
  wire w3979;
  wire w3980;
  wire w3981;
  wire w3982;
  wire w3983;
  wire w3984;
  wire w3985;
  wire w3986;
  wire w3987;
  wire w3988;
  wire w3989;
  wire w3990;
  wire w3991;
  wire w3992;
  wire w3993;
  wire w3994;
  wire w3995;
  wire w3996;
  wire w3997;
  wire w3998;
  wire w3999;
  wire w4000;
  wire w4001;
  wire w4002;
  wire w4003;
  wire w4004;
  wire w4005;
  wire w4006;
  wire w4007;
  wire w4008;
  wire w4009;
  wire w4010;
  wire w4011;
  wire w4012;
  wire w4013;
  wire w4014;
  wire w4015;
  wire w4016;
  wire w4017;
  wire w4018;
  wire w4019;
  wire w4020;
  wire w4021;
  wire w4022;
  wire w4023;
  wire w4024;
  wire w4025;
  wire w4026;
  wire w4027;
  wire w4028;
  wire w4029;
  wire w4030;
  wire w4031;
  wire w4032;
  wire w4033;
  wire w4034;
  wire w4035;
  wire w4036;
  wire w4037;
  wire w4038;
  wire w4039;
  wire w4040;
  wire w4041;
  wire w4042;
  wire w4043;
  wire w4044;
  wire w4045;
  wire w4046;
  wire w4047;
  wire w4048;
  wire w4049;
  wire w4050;
  wire w4051;
  wire w4052;
  wire w4053;
  wire w4054;
  wire w4055;
  wire w4056;
  wire w4058;
  wire w4059;
  wire w4060;
  wire w4061;
  wire w4062;
  wire w4063;
  wire w4064;
  wire w4065;
  wire w4066;
  wire w4067;
  wire w4068;
  wire w4069;
  wire w4070;
  wire w4071;
  wire w4072;
  wire w4073;
  wire w4074;
  wire w4075;
  wire w4076;
  wire w4077;
  wire w4078;
  wire w4079;
  wire w4080;
  wire w4081;
  wire w4082;
  wire w4083;
  wire w4084;
  wire w4085;
  wire w4086;
  wire w4087;
  wire w4088;
  wire w4089;
  wire w4090;
  wire w4091;
  wire w4092;
  wire w4093;
  wire w4094;
  wire w4095;
  wire w4096;
  wire w4097;
  wire w4098;
  wire w4099;
  wire w4100;
  wire w4101;
  wire w4102;
  wire w4103;
  wire w4104;
  wire w4105;
  wire w4106;
  wire w4107;
  wire w4108;
  wire w4109;
  wire w4110;
  wire w4111;
  wire w4112;
  wire w4113;
  wire w4114;
  wire w4115;
  wire w4116;
  wire w4117;
  wire w4118;
  wire w4119;
  wire w4120;
  wire w4121;
  wire w4122;
  wire w4123;
  wire w4124;
  wire w4125;
  wire w4126;
  wire w4127;
  wire w4128;
  wire w4129;
  wire w4130;
  wire w4131;
  wire w4132;
  wire w4133;
  wire w4134;
  wire w4135;
  wire w4136;
  wire w4137;
  wire w4138;
  wire w4139;
  wire w4140;
  wire w4141;
  wire w4142;
  wire w4143;
  wire w4144;
  wire w4145;
  wire w4146;
  wire w4147;
  wire w4148;
  wire w4149;
  wire w4150;
  wire w4151;
  wire w4152;
  wire w4153;
  wire w4154;
  wire w4155;
  wire w4156;
  wire w4157;
  wire w4158;
  wire w4159;
  wire w4160;
  wire w4162;
  wire w4163;
  wire w4164;
  wire w4165;
  wire w4166;
  wire w4167;
  wire w4168;
  wire w4169;
  wire w4170;
  wire w4171;
  wire w4172;
  wire w4173;
  wire w4174;
  wire w4175;
  wire w4176;
  wire w4177;
  wire w4178;
  wire w4179;
  wire w4180;
  wire w4181;
  wire w4182;
  wire w4183;
  wire w4184;
  wire w4185;
  wire w4186;
  wire w4187;
  wire w4188;
  wire w4189;
  wire w4190;
  wire w4191;
  wire w4192;
  wire w4193;
  wire w4194;
  wire w4195;
  wire w4196;
  wire w4197;
  wire w4198;
  wire w4199;
  wire w4200;
  wire w4201;
  wire w4202;
  wire w4203;
  wire w4204;
  wire w4205;
  wire w4206;
  wire w4207;
  wire w4208;
  wire w4209;
  wire w4210;
  wire w4211;
  wire w4212;
  wire w4213;
  wire w4214;
  wire w4215;
  wire w4216;
  wire w4217;
  wire w4218;
  wire w4219;
  wire w4220;
  wire w4221;
  wire w4222;
  wire w4223;
  wire w4224;
  wire w4225;
  wire w4226;
  wire w4227;
  wire w4228;
  wire w4229;
  wire w4230;
  wire w4231;
  wire w4232;
  wire w4233;
  wire w4234;
  wire w4235;
  wire w4236;
  wire w4237;
  wire w4238;
  wire w4239;
  wire w4240;
  wire w4241;
  wire w4242;
  wire w4243;
  wire w4244;
  wire w4245;
  wire w4246;
  wire w4247;
  wire w4248;
  wire w4249;
  wire w4250;
  wire w4251;
  wire w4252;
  wire w4253;
  wire w4254;
  wire w4255;
  wire w4256;
  wire w4257;
  wire w4258;
  wire w4259;
  wire w4260;
  wire w4261;
  wire w4262;
  wire w4263;
  wire w4264;
  wire w4266;
  wire w4267;
  wire w4268;
  wire w4269;
  wire w4270;
  wire w4271;
  wire w4272;
  wire w4273;
  wire w4274;
  wire w4275;
  wire w4276;
  wire w4277;
  wire w4278;
  wire w4279;
  wire w4280;
  wire w4281;
  wire w4282;
  wire w4283;
  wire w4284;
  wire w4285;
  wire w4286;
  wire w4287;
  wire w4288;
  wire w4289;
  wire w4290;
  wire w4291;
  wire w4292;
  wire w4293;
  wire w4294;
  wire w4295;
  wire w4296;
  wire w4297;
  wire w4298;
  wire w4299;
  wire w4300;
  wire w4301;
  wire w4302;
  wire w4303;
  wire w4304;
  wire w4305;
  wire w4306;
  wire w4307;
  wire w4308;
  wire w4309;
  wire w4310;
  wire w4311;
  wire w4312;
  wire w4313;
  wire w4314;
  wire w4315;
  wire w4316;
  wire w4317;
  wire w4318;
  wire w4319;
  wire w4320;
  wire w4321;
  wire w4322;
  wire w4323;
  wire w4324;
  wire w4325;
  wire w4326;
  wire w4327;
  wire w4328;
  wire w4329;
  wire w4330;
  wire w4331;
  wire w4332;
  wire w4333;
  wire w4334;
  wire w4335;
  wire w4336;
  wire w4337;
  wire w4338;
  wire w4339;
  wire w4340;
  wire w4341;
  wire w4342;
  wire w4343;
  wire w4344;
  wire w4345;
  wire w4346;
  wire w4347;
  wire w4348;
  wire w4349;
  wire w4350;
  wire w4351;
  wire w4352;
  wire w4353;
  wire w4354;
  wire w4355;
  wire w4356;
  wire w4357;
  wire w4358;
  wire w4359;
  wire w4360;
  wire w4361;
  wire w4362;
  wire w4363;
  wire w4364;
  wire w4365;
  wire w4366;
  wire w4367;
  wire w4368;
  wire w4370;
  wire w4371;
  wire w4372;
  wire w4373;
  wire w4374;
  wire w4375;
  wire w4376;
  wire w4377;
  wire w4378;
  wire w4379;
  wire w4380;
  wire w4381;
  wire w4382;
  wire w4383;
  wire w4384;
  wire w4385;
  wire w4386;
  wire w4387;
  wire w4388;
  wire w4389;
  wire w4390;
  wire w4391;
  wire w4392;
  wire w4393;
  wire w4394;
  wire w4395;
  wire w4396;
  wire w4397;
  wire w4398;
  wire w4399;
  wire w4400;
  wire w4401;
  wire w4402;
  wire w4403;
  wire w4404;
  wire w4405;
  wire w4406;
  wire w4407;
  wire w4408;
  wire w4409;
  wire w4410;
  wire w4411;
  wire w4412;
  wire w4413;
  wire w4414;
  wire w4415;
  wire w4416;
  wire w4417;
  wire w4418;
  wire w4419;
  wire w4420;
  wire w4421;
  wire w4422;
  wire w4423;
  wire w4424;
  wire w4425;
  wire w4426;
  wire w4427;
  wire w4428;
  wire w4429;
  wire w4430;
  wire w4431;
  wire w4432;
  wire w4433;
  wire w4434;
  wire w4435;
  wire w4436;
  wire w4437;
  wire w4438;
  wire w4439;
  wire w4440;
  wire w4441;
  wire w4442;
  wire w4443;
  wire w4444;
  wire w4445;
  wire w4446;
  wire w4447;
  wire w4448;
  wire w4449;
  wire w4450;
  wire w4451;
  wire w4452;
  wire w4453;
  wire w4454;
  wire w4455;
  wire w4456;
  wire w4457;
  wire w4458;
  wire w4459;
  wire w4460;
  wire w4461;
  wire w4462;
  wire w4463;
  wire w4464;
  wire w4465;
  wire w4466;
  wire w4467;
  wire w4468;
  wire w4469;
  wire w4470;
  wire w4471;
  wire w4472;
  wire w4474;
  wire w4475;
  wire w4476;
  wire w4477;
  wire w4478;
  wire w4479;
  wire w4480;
  wire w4481;
  wire w4482;
  wire w4483;
  wire w4484;
  wire w4485;
  wire w4486;
  wire w4487;
  wire w4488;
  wire w4489;
  wire w4490;
  wire w4491;
  wire w4492;
  wire w4493;
  wire w4494;
  wire w4495;
  wire w4496;
  wire w4497;
  wire w4498;
  wire w4499;
  wire w4500;
  wire w4501;
  wire w4502;
  wire w4503;
  wire w4504;
  wire w4505;
  wire w4506;
  wire w4507;
  wire w4508;
  wire w4509;
  wire w4510;
  wire w4511;
  wire w4512;
  wire w4513;
  wire w4514;
  wire w4515;
  wire w4516;
  wire w4517;
  wire w4518;
  wire w4519;
  wire w4520;
  wire w4521;
  wire w4522;
  wire w4523;
  wire w4524;
  wire w4525;
  wire w4526;
  wire w4527;
  wire w4528;
  wire w4529;
  wire w4530;
  wire w4531;
  wire w4532;
  wire w4533;
  wire w4534;
  wire w4535;
  wire w4536;
  wire w4537;
  wire w4538;
  wire w4539;
  wire w4540;
  wire w4541;
  wire w4542;
  wire w4543;
  wire w4544;
  wire w4545;
  wire w4546;
  wire w4547;
  wire w4548;
  wire w4549;
  wire w4550;
  wire w4551;
  wire w4552;
  wire w4553;
  wire w4554;
  wire w4555;
  wire w4556;
  wire w4557;
  wire w4558;
  wire w4559;
  wire w4560;
  wire w4561;
  wire w4562;
  wire w4563;
  wire w4564;
  wire w4565;
  wire w4566;
  wire w4567;
  wire w4568;
  wire w4569;
  wire w4570;
  wire w4571;
  wire w4572;
  wire w4573;
  wire w4574;
  wire w4575;
  wire w4576;
  wire w4578;
  wire w4579;
  wire w4580;
  wire w4581;
  wire w4582;
  wire w4583;
  wire w4584;
  wire w4585;
  wire w4586;
  wire w4587;
  wire w4588;
  wire w4589;
  wire w4590;
  wire w4591;
  wire w4592;
  wire w4593;
  wire w4594;
  wire w4595;
  wire w4596;
  wire w4597;
  wire w4598;
  wire w4599;
  wire w4600;
  wire w4601;
  wire w4602;
  wire w4603;
  wire w4604;
  wire w4605;
  wire w4606;
  wire w4607;
  wire w4608;
  wire w4609;
  wire w4610;
  wire w4611;
  wire w4612;
  wire w4613;
  wire w4614;
  wire w4615;
  wire w4616;
  wire w4617;
  wire w4618;
  wire w4619;
  wire w4620;
  wire w4621;
  wire w4622;
  wire w4623;
  wire w4624;
  wire w4625;
  wire w4626;
  wire w4627;
  wire w4628;
  wire w4629;
  wire w4630;
  wire w4631;
  wire w4632;
  wire w4633;
  wire w4634;
  wire w4635;
  wire w4636;
  wire w4637;
  wire w4638;
  wire w4639;
  wire w4640;
  wire w4641;
  wire w4642;
  wire w4643;
  wire w4644;
  wire w4645;
  wire w4646;
  wire w4647;
  wire w4648;
  wire w4649;
  wire w4650;
  wire w4651;
  wire w4652;
  wire w4653;
  wire w4654;
  wire w4655;
  wire w4656;
  wire w4657;
  wire w4658;
  wire w4659;
  wire w4660;
  wire w4661;
  wire w4662;
  wire w4663;
  wire w4664;
  wire w4665;
  wire w4666;
  wire w4667;
  wire w4668;
  wire w4669;
  wire w4670;
  wire w4671;
  wire w4672;
  wire w4673;
  wire w4674;
  wire w4675;
  wire w4676;
  wire w4677;
  wire w4678;
  wire w4679;
  wire w4680;
  wire w4682;
  wire w4683;
  wire w4684;
  wire w4685;
  wire w4686;
  wire w4687;
  wire w4688;
  wire w4689;
  wire w4690;
  wire w4691;
  wire w4692;
  wire w4693;
  wire w4694;
  wire w4695;
  wire w4696;
  wire w4697;
  wire w4698;
  wire w4699;
  wire w4700;
  wire w4701;
  wire w4702;
  wire w4703;
  wire w4704;
  wire w4705;
  wire w4706;
  wire w4707;
  wire w4708;
  wire w4709;
  wire w4710;
  wire w4711;
  wire w4712;
  wire w4713;
  wire w4714;
  wire w4715;
  wire w4716;
  wire w4717;
  wire w4718;
  wire w4719;
  wire w4720;
  wire w4721;
  wire w4722;
  wire w4723;
  wire w4724;
  wire w4725;
  wire w4726;
  wire w4727;
  wire w4728;
  wire w4729;
  wire w4730;
  wire w4731;
  wire w4732;
  wire w4733;
  wire w4734;
  wire w4735;
  wire w4736;
  wire w4737;
  wire w4738;
  wire w4739;
  wire w4740;
  wire w4741;
  wire w4742;
  wire w4743;
  wire w4744;
  wire w4745;
  wire w4746;
  wire w4747;
  wire w4748;
  wire w4749;
  wire w4750;
  wire w4751;
  wire w4752;
  wire w4753;
  wire w4754;
  wire w4755;
  wire w4756;
  wire w4757;
  wire w4758;
  wire w4759;
  wire w4760;
  wire w4761;
  wire w4762;
  wire w4763;
  wire w4764;
  wire w4765;
  wire w4766;
  wire w4767;
  wire w4768;
  wire w4769;
  wire w4770;
  wire w4771;
  wire w4772;
  wire w4773;
  wire w4774;
  wire w4775;
  wire w4776;
  wire w4777;
  wire w4778;
  wire w4779;
  wire w4780;
  wire w4781;
  wire w4782;
  wire w4783;
  wire w4784;
  wire w4786;
  wire w4787;
  wire w4788;
  wire w4789;
  wire w4790;
  wire w4791;
  wire w4792;
  wire w4793;
  wire w4794;
  wire w4795;
  wire w4796;
  wire w4797;
  wire w4798;
  wire w4799;
  wire w4800;
  wire w4801;
  wire w4802;
  wire w4803;
  wire w4804;
  wire w4805;
  wire w4806;
  wire w4807;
  wire w4808;
  wire w4809;
  wire w4810;
  wire w4811;
  wire w4812;
  wire w4813;
  wire w4814;
  wire w4815;
  wire w4816;
  wire w4817;
  wire w4818;
  wire w4819;
  wire w4820;
  wire w4821;
  wire w4822;
  wire w4823;
  wire w4824;
  wire w4825;
  wire w4826;
  wire w4827;
  wire w4828;
  wire w4829;
  wire w4830;
  wire w4831;
  wire w4832;
  wire w4833;
  wire w4834;
  wire w4835;
  wire w4836;
  wire w4837;
  wire w4838;
  wire w4839;
  wire w4840;
  wire w4841;
  wire w4842;
  wire w4843;
  wire w4844;
  wire w4845;
  wire w4846;
  wire w4847;
  wire w4848;
  wire w4849;
  wire w4850;
  wire w4851;
  wire w4852;
  wire w4853;
  wire w4854;
  wire w4855;
  wire w4856;
  wire w4857;
  wire w4858;
  wire w4859;
  wire w4860;
  wire w4861;
  wire w4862;
  wire w4863;
  wire w4864;
  wire w4865;
  wire w4866;
  wire w4867;
  wire w4868;
  wire w4869;
  wire w4870;
  wire w4871;
  wire w4872;
  wire w4873;
  wire w4874;
  wire w4875;
  wire w4876;
  wire w4877;
  wire w4878;
  wire w4879;
  wire w4880;
  wire w4881;
  wire w4882;
  wire w4883;
  wire w4884;
  wire w4885;
  wire w4886;
  wire w4887;
  wire w4888;
  wire w4890;
  wire w4891;
  wire w4892;
  wire w4893;
  wire w4894;
  wire w4895;
  wire w4896;
  wire w4897;
  wire w4898;
  wire w4899;
  wire w4900;
  wire w4901;
  wire w4902;
  wire w4903;
  wire w4904;
  wire w4905;
  wire w4906;
  wire w4907;
  wire w4908;
  wire w4909;
  wire w4910;
  wire w4911;
  wire w4912;
  wire w4913;
  wire w4914;
  wire w4915;
  wire w4916;
  wire w4917;
  wire w4918;
  wire w4919;
  wire w4920;
  wire w4921;
  wire w4922;
  wire w4923;
  wire w4924;
  wire w4925;
  wire w4926;
  wire w4927;
  wire w4928;
  wire w4929;
  wire w4930;
  wire w4931;
  wire w4932;
  wire w4933;
  wire w4934;
  wire w4935;
  wire w4936;
  wire w4937;
  wire w4938;
  wire w4939;
  wire w4940;
  wire w4941;
  wire w4942;
  wire w4943;
  wire w4944;
  wire w4945;
  wire w4946;
  wire w4947;
  wire w4948;
  wire w4949;
  wire w4950;
  wire w4951;
  wire w4952;
  wire w4953;
  wire w4954;
  wire w4955;
  wire w4956;
  wire w4957;
  wire w4958;
  wire w4959;
  wire w4960;
  wire w4961;
  wire w4962;
  wire w4963;
  wire w4964;
  wire w4965;
  wire w4966;
  wire w4967;
  wire w4968;
  wire w4969;
  wire w4970;
  wire w4971;
  wire w4972;
  wire w4973;
  wire w4974;
  wire w4975;
  wire w4976;
  wire w4977;
  wire w4978;
  wire w4979;
  wire w4980;
  wire w4981;
  wire w4982;
  wire w4983;
  wire w4984;
  wire w4985;
  wire w4986;
  wire w4987;
  wire w4988;
  wire w4989;
  wire w4990;
  wire w4991;
  wire w4992;
  wire w4994;
  wire w4995;
  wire w4996;
  wire w4997;
  wire w4998;
  wire w4999;
  wire w5000;
  wire w5001;
  wire w5002;
  wire w5003;
  wire w5004;
  wire w5005;
  wire w5006;
  wire w5007;
  wire w5008;
  wire w5009;
  wire w5010;
  wire w5011;
  wire w5012;
  wire w5013;
  wire w5014;
  wire w5015;
  wire w5016;
  wire w5017;
  wire w5018;
  wire w5019;
  wire w5020;
  wire w5021;
  wire w5022;
  wire w5023;
  wire w5024;
  wire w5025;
  wire w5026;
  wire w5027;
  wire w5028;
  wire w5029;
  wire w5030;
  wire w5031;
  wire w5032;
  wire w5033;
  wire w5034;
  wire w5035;
  wire w5036;
  wire w5037;
  wire w5038;
  wire w5039;
  wire w5040;
  wire w5041;
  wire w5042;
  wire w5043;
  wire w5044;
  wire w5045;
  wire w5046;
  wire w5047;
  wire w5048;
  wire w5049;
  wire w5050;
  wire w5051;
  wire w5052;
  wire w5053;
  wire w5054;
  wire w5055;
  wire w5056;
  wire w5057;
  wire w5058;
  wire w5059;
  wire w5060;
  wire w5061;
  wire w5062;
  wire w5063;
  wire w5064;
  wire w5065;
  wire w5066;
  wire w5067;
  wire w5068;
  wire w5069;
  wire w5070;
  wire w5071;
  wire w5072;
  wire w5073;
  wire w5074;
  wire w5075;
  wire w5076;
  wire w5077;
  wire w5078;
  wire w5079;
  wire w5080;
  wire w5081;
  wire w5082;
  wire w5083;
  wire w5084;
  wire w5085;
  wire w5086;
  wire w5087;
  wire w5088;
  wire w5089;
  wire w5090;
  wire w5091;
  wire w5092;
  wire w5093;
  wire w5094;
  wire w5095;
  wire w5096;
  wire w5098;
  wire w5099;
  wire w5100;
  wire w5101;
  wire w5102;
  wire w5103;
  wire w5104;
  wire w5105;
  wire w5106;
  wire w5107;
  wire w5108;
  wire w5109;
  wire w5110;
  wire w5111;
  wire w5112;
  wire w5113;
  wire w5114;
  wire w5115;
  wire w5116;
  wire w5117;
  wire w5118;
  wire w5119;
  wire w5120;
  wire w5121;
  wire w5122;
  wire w5123;
  wire w5124;
  wire w5125;
  wire w5126;
  wire w5127;
  wire w5128;
  wire w5129;
  wire w5130;
  wire w5131;
  wire w5132;
  wire w5133;
  wire w5134;
  wire w5135;
  wire w5136;
  wire w5137;
  wire w5138;
  wire w5139;
  wire w5140;
  wire w5141;
  wire w5142;
  wire w5143;
  wire w5144;
  wire w5145;
  wire w5146;
  wire w5147;
  wire w5148;
  wire w5149;
  wire w5150;
  wire w5151;
  wire w5152;
  wire w5153;
  wire w5154;
  wire w5155;
  wire w5156;
  wire w5157;
  wire w5158;
  wire w5159;
  wire w5160;
  wire w5161;
  wire w5162;
  wire w5163;
  wire w5164;
  wire w5165;
  wire w5166;
  wire w5167;
  wire w5168;
  wire w5169;
  wire w5170;
  wire w5171;
  wire w5172;
  wire w5173;
  wire w5174;
  wire w5175;
  wire w5176;
  wire w5177;
  wire w5178;
  wire w5179;
  wire w5180;
  wire w5181;
  wire w5182;
  wire w5183;
  wire w5184;
  wire w5185;
  wire w5186;
  wire w5187;
  wire w5188;
  wire w5189;
  wire w5190;
  wire w5191;
  wire w5192;
  wire w5193;
  wire w5194;
  wire w5195;
  wire w5196;
  wire w5197;
  wire w5198;
  wire w5199;
  wire w5200;
  wire w5202;
  wire w5203;
  wire w5204;
  wire w5205;
  wire w5206;
  wire w5207;
  wire w5208;
  wire w5209;
  wire w5210;
  wire w5211;
  wire w5212;
  wire w5213;
  wire w5214;
  wire w5215;
  wire w5216;
  wire w5217;
  wire w5218;
  wire w5219;
  wire w5220;
  wire w5221;
  wire w5222;
  wire w5223;
  wire w5224;
  wire w5225;
  wire w5226;
  wire w5227;
  wire w5228;
  wire w5229;
  wire w5230;
  wire w5231;
  wire w5232;
  wire w5233;
  wire w5234;
  wire w5235;
  wire w5236;
  wire w5237;
  wire w5238;
  wire w5239;
  wire w5240;
  wire w5241;
  wire w5242;
  wire w5243;
  wire w5244;
  wire w5245;
  wire w5246;
  wire w5247;
  wire w5248;
  wire w5249;
  wire w5250;
  wire w5251;
  wire w5252;
  wire w5253;
  wire w5254;
  wire w5255;
  wire w5256;
  wire w5257;
  wire w5258;
  wire w5259;
  wire w5260;
  wire w5261;
  wire w5262;
  wire w5263;
  wire w5264;
  wire w5265;
  wire w5266;
  wire w5267;
  wire w5268;
  wire w5269;
  wire w5270;
  wire w5271;
  wire w5272;
  wire w5273;
  wire w5274;
  wire w5275;
  wire w5276;
  wire w5277;
  wire w5278;
  wire w5279;
  wire w5280;
  wire w5281;
  wire w5282;
  wire w5283;
  wire w5284;
  wire w5285;
  wire w5286;
  wire w5287;
  wire w5288;
  wire w5289;
  wire w5290;
  wire w5291;
  wire w5292;
  wire w5293;
  wire w5294;
  wire w5295;
  wire w5296;
  wire w5297;
  wire w5298;
  wire w5299;
  wire w5300;
  wire w5301;
  wire w5302;
  wire w5303;
  wire w5304;
  wire w5306;
  wire w5307;
  wire w5308;
  wire w5309;
  wire w5310;
  wire w5311;
  wire w5312;
  wire w5313;
  wire w5314;
  wire w5315;
  wire w5316;
  wire w5317;
  wire w5318;
  wire w5319;
  wire w5320;
  wire w5321;
  wire w5322;
  wire w5323;
  wire w5324;
  wire w5325;
  wire w5326;
  wire w5327;
  wire w5328;
  wire w5329;
  wire w5330;
  wire w5331;
  wire w5332;
  wire w5333;
  wire w5334;
  wire w5335;
  wire w5336;
  wire w5337;
  wire w5338;
  wire w5339;
  wire w5340;
  wire w5341;
  wire w5342;
  wire w5343;
  wire w5344;
  wire w5345;
  wire w5346;
  wire w5347;
  wire w5348;
  wire w5349;
  wire w5350;
  wire w5351;
  wire w5352;
  wire w5353;
  wire w5354;
  wire w5355;
  wire w5356;
  wire w5357;
  wire w5358;
  wire w5359;
  wire w5360;
  wire w5361;
  wire w5362;
  wire w5363;
  wire w5364;
  wire w5365;
  wire w5366;
  wire w5367;
  wire w5368;
  wire w5369;
  wire w5370;
  wire w5371;
  wire w5372;
  wire w5373;
  wire w5374;
  wire w5375;
  wire w5376;
  wire w5377;
  wire w5378;
  wire w5379;
  wire w5380;
  wire w5381;
  wire w5382;
  wire w5383;
  wire w5384;
  wire w5385;
  wire w5386;
  wire w5387;
  wire w5388;
  wire w5389;
  wire w5390;
  wire w5391;
  wire w5392;
  wire w5393;
  wire w5394;
  wire w5395;
  wire w5396;
  wire w5397;
  wire w5398;
  wire w5399;
  wire w5400;
  wire w5401;
  wire w5402;
  wire w5403;
  wire w5404;
  wire w5405;
  wire w5406;
  wire w5407;
  wire w5408;
  wire w5410;
  wire w5411;
  wire w5412;
  wire w5413;
  wire w5414;
  wire w5415;
  wire w5416;
  wire w5417;
  wire w5418;
  wire w5419;
  wire w5420;
  wire w5421;
  wire w5422;
  wire w5423;
  wire w5424;
  wire w5425;
  wire w5426;
  wire w5427;
  wire w5428;
  wire w5429;
  wire w5430;
  wire w5431;
  wire w5432;
  wire w5433;
  wire w5434;
  wire w5435;
  wire w5436;
  wire w5437;
  wire w5438;
  wire w5439;
  wire w5440;
  wire w5441;
  wire w5442;
  wire w5443;
  wire w5444;
  wire w5445;
  wire w5446;
  wire w5447;
  wire w5448;
  wire w5449;
  wire w5450;
  wire w5451;
  wire w5452;
  wire w5453;
  wire w5454;
  wire w5455;
  wire w5456;
  wire w5457;
  wire w5458;
  wire w5459;
  wire w5460;
  wire w5461;
  wire w5462;
  wire w5463;
  wire w5464;
  wire w5465;
  wire w5466;
  wire w5467;
  wire w5468;
  wire w5469;
  wire w5470;
  wire w5471;
  wire w5472;
  wire w5473;
  wire w5474;
  wire w5475;
  wire w5476;
  wire w5477;
  wire w5478;
  wire w5479;
  wire w5480;
  wire w5481;
  wire w5482;
  wire w5483;
  wire w5484;
  wire w5485;
  wire w5486;
  wire w5487;
  wire w5488;
  wire w5489;
  wire w5490;
  wire w5491;
  wire w5492;
  wire w5493;
  wire w5494;
  wire w5495;
  wire w5496;
  wire w5497;
  wire w5498;
  wire w5499;
  wire w5500;
  wire w5501;
  wire w5502;
  wire w5503;
  wire w5504;
  wire w5505;
  wire w5506;
  wire w5507;
  wire w5508;
  wire w5509;
  wire w5510;
  wire w5511;
  wire w5512;
  wire w5514;
  wire w5515;
  wire w5516;
  wire w5517;
  wire w5518;
  wire w5519;
  wire w5520;
  wire w5521;
  wire w5522;
  wire w5523;
  wire w5524;
  wire w5525;
  wire w5526;
  wire w5527;
  wire w5528;
  wire w5529;
  wire w5530;
  wire w5531;
  wire w5532;
  wire w5533;
  wire w5534;
  wire w5535;
  wire w5536;
  wire w5537;
  wire w5538;
  wire w5539;
  wire w5540;
  wire w5541;
  wire w5542;
  wire w5543;
  wire w5544;
  wire w5545;
  wire w5546;
  wire w5547;
  wire w5548;
  wire w5549;
  wire w5550;
  wire w5551;
  wire w5552;
  wire w5553;
  wire w5554;
  wire w5555;
  wire w5556;
  wire w5557;
  wire w5558;
  wire w5559;
  wire w5560;
  wire w5561;
  wire w5562;
  wire w5563;
  wire w5564;
  wire w5565;
  wire w5566;
  wire w5567;
  wire w5568;
  wire w5569;
  wire w5570;
  wire w5571;
  wire w5572;
  wire w5573;
  wire w5574;
  wire w5575;
  wire w5576;
  wire w5577;
  wire w5578;
  wire w5579;
  wire w5580;
  wire w5581;
  wire w5582;
  wire w5583;
  wire w5584;
  wire w5585;
  wire w5586;
  wire w5587;
  wire w5588;
  wire w5589;
  wire w5590;
  wire w5591;
  wire w5592;
  wire w5593;
  wire w5594;
  wire w5595;
  wire w5596;
  wire w5597;
  wire w5598;
  wire w5599;
  wire w5600;
  wire w5601;
  wire w5602;
  wire w5603;
  wire w5604;
  wire w5605;
  wire w5606;
  wire w5607;
  wire w5608;
  wire w5609;
  wire w5610;
  wire w5611;
  wire w5612;
  wire w5613;
  wire w5614;
  wire w5615;
  wire w5616;
  wire w5618;
  wire w5619;
  wire w5620;
  wire w5621;
  wire w5622;
  wire w5623;
  wire w5624;
  wire w5625;
  wire w5626;
  wire w5627;
  wire w5628;
  wire w5629;
  wire w5630;
  wire w5631;
  wire w5632;
  wire w5633;
  wire w5634;
  wire w5635;
  wire w5636;
  wire w5637;
  wire w5638;
  wire w5639;
  wire w5640;
  wire w5641;
  wire w5642;
  wire w5643;
  wire w5644;
  wire w5645;
  wire w5646;
  wire w5647;
  wire w5648;
  wire w5649;
  wire w5650;
  wire w5651;
  wire w5652;
  wire w5653;
  wire w5654;
  wire w5655;
  wire w5656;
  wire w5657;
  wire w5658;
  wire w5659;
  wire w5660;
  wire w5661;
  wire w5662;
  wire w5663;
  wire w5664;
  wire w5665;
  wire w5666;
  wire w5667;
  wire w5668;
  wire w5669;
  wire w5670;
  wire w5671;
  wire w5672;
  wire w5673;
  wire w5674;
  wire w5675;
  wire w5676;
  wire w5677;
  wire w5678;
  wire w5679;
  wire w5680;
  wire w5681;
  wire w5682;
  wire w5683;
  wire w5684;
  wire w5685;
  wire w5686;
  wire w5687;
  wire w5688;
  wire w5689;
  wire w5690;
  wire w5691;
  wire w5692;
  wire w5693;
  wire w5694;
  wire w5695;
  wire w5696;
  wire w5697;
  wire w5698;
  wire w5699;
  wire w5700;
  wire w5701;
  wire w5702;
  wire w5703;
  wire w5704;
  wire w5705;
  wire w5706;
  wire w5707;
  wire w5708;
  wire w5709;
  wire w5710;
  wire w5711;
  wire w5712;
  wire w5713;
  wire w5714;
  wire w5715;
  wire w5716;
  wire w5717;
  wire w5718;
  wire w5719;
  wire w5720;
  wire w5722;
  wire w5723;
  wire w5724;
  wire w5725;
  wire w5726;
  wire w5727;
  wire w5728;
  wire w5729;
  wire w5730;
  wire w5731;
  wire w5732;
  wire w5733;
  wire w5734;
  wire w5735;
  wire w5736;
  wire w5737;
  wire w5738;
  wire w5739;
  wire w5740;
  wire w5741;
  wire w5742;
  wire w5743;
  wire w5744;
  wire w5745;
  wire w5746;
  wire w5747;
  wire w5748;
  wire w5749;
  wire w5750;
  wire w5751;
  wire w5752;
  wire w5753;
  wire w5754;
  wire w5755;
  wire w5756;
  wire w5757;
  wire w5758;
  wire w5759;
  wire w5760;
  wire w5761;
  wire w5762;
  wire w5763;
  wire w5764;
  wire w5765;
  wire w5766;
  wire w5767;
  wire w5768;
  wire w5769;
  wire w5770;
  wire w5771;
  wire w5772;
  wire w5773;
  wire w5774;
  wire w5775;
  wire w5776;
  wire w5777;
  wire w5778;
  wire w5779;
  wire w5780;
  wire w5781;
  wire w5782;
  wire w5783;
  wire w5784;
  wire w5785;
  wire w5786;
  wire w5787;
  wire w5788;
  wire w5789;
  wire w5790;
  wire w5791;
  wire w5792;
  wire w5793;
  wire w5794;
  wire w5795;
  wire w5796;
  wire w5797;
  wire w5798;
  wire w5799;
  wire w5800;
  wire w5801;
  wire w5802;
  wire w5803;
  wire w5804;
  wire w5805;
  wire w5806;
  wire w5807;
  wire w5808;
  wire w5809;
  wire w5810;
  wire w5811;
  wire w5812;
  wire w5813;
  wire w5814;
  wire w5815;
  wire w5816;
  wire w5817;
  wire w5818;
  wire w5819;
  wire w5820;
  wire w5821;
  wire w5822;
  wire w5823;
  wire w5824;
  wire w5826;
  wire w5827;
  wire w5828;
  wire w5829;
  wire w5830;
  wire w5831;
  wire w5832;
  wire w5833;
  wire w5834;
  wire w5835;
  wire w5836;
  wire w5837;
  wire w5838;
  wire w5839;
  wire w5840;
  wire w5841;
  wire w5842;
  wire w5843;
  wire w5844;
  wire w5845;
  wire w5846;
  wire w5847;
  wire w5848;
  wire w5849;
  wire w5850;
  wire w5851;
  wire w5852;
  wire w5853;
  wire w5854;
  wire w5855;
  wire w5856;
  wire w5857;
  wire w5858;
  wire w5859;
  wire w5860;
  wire w5861;
  wire w5862;
  wire w5863;
  wire w5864;
  wire w5865;
  wire w5866;
  wire w5867;
  wire w5868;
  wire w5869;
  wire w5870;
  wire w5871;
  wire w5872;
  wire w5873;
  wire w5874;
  wire w5875;
  wire w5876;
  wire w5877;
  wire w5878;
  wire w5879;
  wire w5880;
  wire w5881;
  wire w5882;
  wire w5883;
  wire w5884;
  wire w5885;
  wire w5886;
  wire w5887;
  wire w5888;
  wire w5889;
  wire w5890;
  wire w5891;
  wire w5892;
  wire w5893;
  wire w5894;
  wire w5895;
  wire w5896;
  wire w5897;
  wire w5898;
  wire w5899;
  wire w5900;
  wire w5901;
  wire w5902;
  wire w5903;
  wire w5904;
  wire w5905;
  wire w5906;
  wire w5907;
  wire w5908;
  wire w5909;
  wire w5910;
  wire w5911;
  wire w5912;
  wire w5913;
  wire w5914;
  wire w5915;
  wire w5916;
  wire w5917;
  wire w5918;
  wire w5919;
  wire w5920;
  wire w5921;
  wire w5922;
  wire w5923;
  wire w5924;
  wire w5925;
  wire w5926;
  wire w5927;
  wire w5928;
  wire w5930;
  wire w5931;
  wire w5932;
  wire w5933;
  wire w5934;
  wire w5935;
  wire w5936;
  wire w5937;
  wire w5938;
  wire w5939;
  wire w5940;
  wire w5941;
  wire w5942;
  wire w5943;
  wire w5944;
  wire w5945;
  wire w5946;
  wire w5947;
  wire w5948;
  wire w5949;
  wire w5950;
  wire w5951;
  wire w5952;
  wire w5953;
  wire w5954;
  wire w5955;
  wire w5956;
  wire w5957;
  wire w5958;
  wire w5959;
  wire w5960;
  wire w5961;
  wire w5962;
  wire w5963;
  wire w5964;
  wire w5965;
  wire w5966;
  wire w5967;
  wire w5968;
  wire w5969;
  wire w5970;
  wire w5971;
  wire w5972;
  wire w5973;
  wire w5974;
  wire w5975;
  wire w5976;
  wire w5977;
  wire w5978;
  wire w5979;
  wire w5980;
  wire w5981;
  wire w5982;
  wire w5983;
  wire w5984;
  wire w5985;
  wire w5986;
  wire w5987;
  wire w5988;
  wire w5989;
  wire w5990;
  wire w5991;
  wire w5992;
  wire w5993;
  wire w5994;
  wire w5995;
  wire w5996;
  wire w5997;
  wire w5998;
  wire w5999;
  wire w6000;
  wire w6001;
  wire w6002;
  wire w6003;
  wire w6004;
  wire w6005;
  wire w6006;
  wire w6007;
  wire w6008;
  wire w6009;
  wire w6010;
  wire w6011;
  wire w6012;
  wire w6013;
  wire w6014;
  wire w6015;
  wire w6016;
  wire w6017;
  wire w6018;
  wire w6019;
  wire w6020;
  wire w6021;
  wire w6022;
  wire w6023;
  wire w6024;
  wire w6025;
  wire w6026;
  wire w6027;
  wire w6028;
  wire w6029;
  wire w6030;
  wire w6031;
  wire w6032;
  wire w6034;
  wire w6035;
  wire w6036;
  wire w6037;
  wire w6038;
  wire w6039;
  wire w6040;
  wire w6041;
  wire w6042;
  wire w6043;
  wire w6044;
  wire w6045;
  wire w6046;
  wire w6047;
  wire w6048;
  wire w6049;
  wire w6050;
  wire w6051;
  wire w6052;
  wire w6053;
  wire w6054;
  wire w6055;
  wire w6056;
  wire w6057;
  wire w6058;
  wire w6059;
  wire w6060;
  wire w6061;
  wire w6062;
  wire w6063;
  wire w6064;
  wire w6065;
  wire w6066;
  wire w6067;
  wire w6068;
  wire w6069;
  wire w6070;
  wire w6071;
  wire w6072;
  wire w6073;
  wire w6074;
  wire w6075;
  wire w6076;
  wire w6077;
  wire w6078;
  wire w6079;
  wire w6080;
  wire w6081;
  wire w6082;
  wire w6083;
  wire w6084;
  wire w6085;
  wire w6086;
  wire w6087;
  wire w6088;
  wire w6089;
  wire w6090;
  wire w6091;
  wire w6092;
  wire w6093;
  wire w6094;
  wire w6095;
  wire w6096;
  wire w6097;
  wire w6098;
  wire w6099;
  wire w6100;
  wire w6101;
  wire w6102;
  wire w6103;
  wire w6104;
  wire w6105;
  wire w6106;
  wire w6107;
  wire w6108;
  wire w6109;
  wire w6110;
  wire w6111;
  wire w6112;
  wire w6113;
  wire w6114;
  wire w6115;
  wire w6116;
  wire w6117;
  wire w6118;
  wire w6119;
  wire w6120;
  wire w6121;
  wire w6122;
  wire w6123;
  wire w6124;
  wire w6125;
  wire w6126;
  wire w6127;
  wire w6128;
  wire w6129;
  wire w6130;
  wire w6131;
  wire w6132;
  wire w6133;
  wire w6134;
  wire w6135;
  wire w6136;
  wire w6138;
  wire w6139;
  wire w6140;
  wire w6141;
  wire w6142;
  wire w6143;
  wire w6144;
  wire w6145;
  wire w6146;
  wire w6147;
  wire w6148;
  wire w6149;
  wire w6150;
  wire w6151;
  wire w6152;
  wire w6153;
  wire w6154;
  wire w6155;
  wire w6156;
  wire w6157;
  wire w6158;
  wire w6159;
  wire w6160;
  wire w6161;
  wire w6162;
  wire w6163;
  wire w6164;
  wire w6165;
  wire w6166;
  wire w6167;
  wire w6168;
  wire w6169;
  wire w6170;
  wire w6171;
  wire w6172;
  wire w6173;
  wire w6174;
  wire w6175;
  wire w6176;
  wire w6177;
  wire w6178;
  wire w6179;
  wire w6180;
  wire w6181;
  wire w6182;
  wire w6183;
  wire w6184;
  wire w6185;
  wire w6186;
  wire w6187;
  wire w6188;
  wire w6189;
  wire w6190;
  wire w6191;
  wire w6192;
  wire w6193;
  wire w6194;
  wire w6195;
  wire w6196;
  wire w6197;
  wire w6198;
  wire w6199;
  wire w6200;
  wire w6201;
  wire w6202;
  wire w6203;
  wire w6204;
  wire w6205;
  wire w6206;
  wire w6207;
  wire w6208;
  wire w6209;
  wire w6210;
  wire w6211;
  wire w6212;
  wire w6213;
  wire w6214;
  wire w6215;
  wire w6216;
  wire w6217;
  wire w6218;
  wire w6219;
  wire w6220;
  wire w6221;
  wire w6222;
  wire w6223;
  wire w6224;
  wire w6225;
  wire w6226;
  wire w6227;
  wire w6228;
  wire w6229;
  wire w6230;
  wire w6231;
  wire w6232;
  wire w6233;
  wire w6234;
  wire w6235;
  wire w6236;
  wire w6237;
  wire w6238;
  wire w6239;
  wire w6240;
  wire w6242;
  wire w6243;
  wire w6244;
  wire w6245;
  wire w6246;
  wire w6247;
  wire w6248;
  wire w6249;
  wire w6250;
  wire w6251;
  wire w6252;
  wire w6253;
  wire w6254;
  wire w6255;
  wire w6256;
  wire w6257;
  wire w6258;
  wire w6259;
  wire w6260;
  wire w6261;
  wire w6262;
  wire w6263;
  wire w6264;
  wire w6265;
  wire w6266;
  wire w6267;
  wire w6268;
  wire w6269;
  wire w6270;
  wire w6271;
  wire w6272;
  wire w6273;
  wire w6274;
  wire w6275;
  wire w6276;
  wire w6277;
  wire w6278;
  wire w6279;
  wire w6280;
  wire w6281;
  wire w6282;
  wire w6283;
  wire w6284;
  wire w6285;
  wire w6286;
  wire w6287;
  wire w6288;
  wire w6289;
  wire w6290;
  wire w6291;
  wire w6292;
  wire w6293;
  wire w6294;
  wire w6295;
  wire w6296;
  wire w6297;
  wire w6298;
  wire w6299;
  wire w6300;
  wire w6301;
  wire w6302;
  wire w6303;
  wire w6304;
  wire w6305;
  wire w6306;
  wire w6307;
  wire w6308;
  wire w6309;
  wire w6310;
  wire w6311;
  wire w6312;
  wire w6313;
  wire w6314;
  wire w6315;
  wire w6316;
  wire w6317;
  wire w6318;
  wire w6319;
  wire w6320;
  wire w6321;
  wire w6322;
  wire w6323;
  wire w6324;
  wire w6325;
  wire w6326;
  wire w6327;
  wire w6328;
  wire w6329;
  wire w6330;
  wire w6331;
  wire w6332;
  wire w6333;
  wire w6334;
  wire w6335;
  wire w6336;
  wire w6337;
  wire w6338;
  wire w6339;
  wire w6340;
  wire w6341;
  wire w6342;
  wire w6343;
  wire w6344;
  wire w6346;
  wire w6347;
  wire w6348;
  wire w6349;
  wire w6350;
  wire w6351;
  wire w6352;
  wire w6353;
  wire w6354;
  wire w6355;
  wire w6356;
  wire w6357;
  wire w6358;
  wire w6359;
  wire w6360;
  wire w6361;
  wire w6362;
  wire w6363;
  wire w6364;
  wire w6365;
  wire w6366;
  wire w6367;
  wire w6368;
  wire w6369;
  wire w6370;
  wire w6371;
  wire w6372;
  wire w6373;
  wire w6374;
  wire w6375;
  wire w6376;
  wire w6377;
  wire w6378;
  wire w6379;
  wire w6380;
  wire w6381;
  wire w6382;
  wire w6383;
  wire w6384;
  wire w6385;
  wire w6386;
  wire w6387;
  wire w6388;
  wire w6389;
  wire w6390;
  wire w6391;
  wire w6392;
  wire w6393;
  wire w6394;
  wire w6395;
  wire w6396;
  wire w6397;
  wire w6398;
  wire w6399;
  wire w6400;
  wire w6401;
  wire w6402;
  wire w6403;
  wire w6404;
  wire w6405;
  wire w6406;
  wire w6407;
  wire w6408;
  wire w6409;
  wire w6410;
  wire w6411;
  wire w6412;
  wire w6413;
  wire w6414;
  wire w6415;
  wire w6416;
  wire w6417;
  wire w6418;
  wire w6419;
  wire w6420;
  wire w6421;
  wire w6422;
  wire w6423;
  wire w6424;
  wire w6425;
  wire w6426;
  wire w6427;
  wire w6428;
  wire w6429;
  wire w6430;
  wire w6431;
  wire w6432;
  wire w6433;
  wire w6434;
  wire w6435;
  wire w6436;
  wire w6437;
  wire w6438;
  wire w6439;
  wire w6440;
  wire w6441;
  wire w6442;
  wire w6443;
  wire w6444;
  wire w6445;
  wire w6446;
  wire w6447;
  wire w6448;
  wire w6450;
  wire w6451;
  wire w6452;
  wire w6453;
  wire w6454;
  wire w6455;
  wire w6456;
  wire w6457;
  wire w6458;
  wire w6459;
  wire w6460;
  wire w6461;
  wire w6462;
  wire w6463;
  wire w6464;
  wire w6465;
  wire w6466;
  wire w6467;
  wire w6468;
  wire w6469;
  wire w6470;
  wire w6471;
  wire w6472;
  wire w6473;
  wire w6474;
  wire w6475;
  wire w6476;
  wire w6477;
  wire w6478;
  wire w6479;
  wire w6480;
  wire w6481;
  wire w6482;
  wire w6483;
  wire w6484;
  wire w6485;
  wire w6486;
  wire w6487;
  wire w6488;
  wire w6489;
  wire w6490;
  wire w6491;
  wire w6492;
  wire w6493;
  wire w6494;
  wire w6495;
  wire w6496;
  wire w6497;
  wire w6498;
  wire w6499;
  wire w6500;
  wire w6501;
  wire w6502;
  wire w6503;
  wire w6504;
  wire w6505;
  wire w6506;
  wire w6507;
  wire w6508;
  wire w6509;
  wire w6510;
  wire w6511;
  wire w6512;
  wire w6513;
  wire w6514;
  wire w6515;
  wire w6516;
  wire w6517;
  wire w6518;
  wire w6519;
  wire w6520;
  wire w6521;
  wire w6522;
  wire w6523;
  wire w6524;
  wire w6525;
  wire w6526;
  wire w6527;
  wire w6528;
  wire w6529;
  wire w6530;
  wire w6531;
  wire w6532;
  wire w6533;
  wire w6534;
  wire w6535;
  wire w6536;
  wire w6537;
  wire w6538;
  wire w6539;
  wire w6540;
  wire w6541;
  wire w6542;
  wire w6543;
  wire w6544;
  wire w6545;
  wire w6546;
  wire w6547;
  wire w6548;
  wire w6549;
  wire w6550;
  wire w6551;
  wire w6552;
  wire w6554;
  wire w6555;
  wire w6556;
  wire w6557;
  wire w6558;
  wire w6559;
  wire w6560;
  wire w6561;
  wire w6562;
  wire w6563;
  wire w6564;
  wire w6565;
  wire w6566;
  wire w6567;
  wire w6568;
  wire w6569;
  wire w6570;
  wire w6571;
  wire w6572;
  wire w6573;
  wire w6574;
  wire w6575;
  wire w6576;
  wire w6577;
  wire w6578;
  wire w6579;
  wire w6580;
  wire w6581;
  wire w6582;
  wire w6583;
  wire w6584;
  wire w6585;
  wire w6586;
  wire w6587;
  wire w6588;
  wire w6589;
  wire w6590;
  wire w6591;
  wire w6592;
  wire w6593;
  wire w6594;
  wire w6595;
  wire w6596;
  wire w6597;
  wire w6598;
  wire w6599;
  wire w6600;
  wire w6601;
  wire w6602;
  wire w6603;
  wire w6604;
  wire w6605;
  wire w6606;
  wire w6607;
  wire w6608;
  wire w6609;
  wire w6610;
  wire w6611;
  wire w6612;
  wire w6613;
  wire w6614;
  wire w6615;
  wire w6616;
  wire w6617;
  wire w6618;
  wire w6619;
  wire w6620;
  wire w6621;
  wire w6622;
  wire w6623;
  wire w6624;
  wire w6625;
  wire w6626;
  wire w6627;
  wire w6628;
  wire w6629;
  wire w6630;
  wire w6631;
  wire w6632;
  wire w6633;
  wire w6634;
  wire w6635;
  wire w6636;
  wire w6637;
  wire w6638;
  wire w6639;
  wire w6640;
  wire w6641;
  wire w6642;
  wire w6643;
  wire w6644;
  wire w6645;
  wire w6646;
  wire w6647;
  wire w6648;
  wire w6649;
  wire w6650;
  wire w6651;
  wire w6652;
  wire w6653;
  wire w6654;
  wire w6655;
  wire w6656;
  wire w6658;
  wire w6659;
  wire w6660;
  wire w6661;
  wire w6662;
  wire w6663;
  wire w6664;
  wire w6665;
  wire w6666;
  wire w6667;
  wire w6668;
  wire w6669;
  wire w6670;
  wire w6671;
  wire w6672;
  wire w6673;
  wire w6674;
  wire w6675;
  wire w6676;
  wire w6677;
  wire w6678;
  wire w6679;
  wire w6680;
  wire w6681;
  wire w6682;
  wire w6683;
  wire w6684;
  wire w6685;
  wire w6686;
  wire w6687;
  wire w6688;
  wire w6689;
  wire w6690;
  wire w6691;
  wire w6692;
  wire w6693;
  wire w6694;
  wire w6695;
  wire w6696;
  wire w6697;
  wire w6698;
  wire w6699;
  wire w6700;
  wire w6701;
  wire w6702;
  wire w6703;
  wire w6704;
  wire w6705;
  wire w6706;
  wire w6707;
  wire w6708;
  wire w6709;
  wire w6710;
  wire w6711;
  wire w6712;
  wire w6713;
  wire w6714;
  wire w6715;
  wire w6716;
  wire w6717;
  wire w6718;
  wire w6719;
  wire w6720;
  wire w6721;
  wire w6722;
  wire w6723;
  wire w6724;
  wire w6725;
  wire w6726;
  wire w6727;
  wire w6728;
  wire w6729;
  wire w6730;
  wire w6731;
  wire w6732;
  wire w6733;
  wire w6734;
  wire w6735;
  wire w6736;
  wire w6737;
  wire w6738;
  wire w6739;
  wire w6740;
  wire w6741;
  wire w6742;
  wire w6743;
  wire w6744;
  wire w6745;
  wire w6746;
  wire w6747;
  wire w6748;
  wire w6749;
  wire w6750;
  wire w6751;
  wire w6752;
  wire w6753;
  wire w6754;
  wire w6755;
  wire w6756;
  wire w6757;
  wire w6758;
  wire w6759;
  wire w6760;
  wire w6762;
  wire w6763;
  wire w6764;
  wire w6765;
  wire w6766;
  wire w6767;
  wire w6768;
  wire w6769;
  wire w6770;
  wire w6771;
  wire w6772;
  wire w6773;
  wire w6774;
  wire w6775;
  wire w6776;
  wire w6777;
  wire w6778;
  wire w6779;
  wire w6780;
  wire w6781;
  wire w6782;
  wire w6783;
  wire w6784;
  wire w6785;
  wire w6786;
  wire w6787;
  wire w6788;
  wire w6789;
  wire w6790;
  wire w6791;
  wire w6792;
  wire w6793;
  wire w6794;
  wire w6795;
  wire w6796;
  wire w6797;
  wire w6798;
  wire w6799;
  wire w6800;
  wire w6801;
  wire w6802;
  wire w6803;
  wire w6804;
  wire w6805;
  wire w6806;
  wire w6807;
  wire w6808;
  wire w6809;
  wire w6810;
  wire w6811;
  wire w6812;
  wire w6813;
  wire w6814;
  wire w6815;
  wire w6816;
  wire w6817;
  wire w6818;
  wire w6819;
  wire w6820;
  wire w6821;
  wire w6822;
  wire w6823;
  wire w6824;
  wire w6825;
  wire w6826;
  wire w6827;
  wire w6828;
  wire w6829;
  wire w6830;
  wire w6831;
  wire w6832;
  wire w6833;
  wire w6834;
  wire w6835;
  wire w6836;
  wire w6837;
  wire w6838;
  wire w6839;
  wire w6840;
  wire w6841;
  wire w6842;
  wire w6843;
  wire w6844;
  wire w6845;
  wire w6846;
  wire w6847;
  wire w6848;
  wire w6849;
  wire w6850;
  wire w6851;
  wire w6852;
  wire w6853;
  wire w6854;
  wire w6855;
  wire w6856;
  wire w6857;
  wire w6858;
  wire w6859;
  wire w6860;
  wire w6861;
  wire w6862;
  wire w6863;
  wire w6864;
  wire w6866;
  wire w6867;
  wire w6868;
  wire w6869;
  wire w6870;
  wire w6871;
  wire w6872;
  wire w6873;
  wire w6874;
  wire w6875;
  wire w6876;
  wire w6877;
  wire w6878;
  wire w6879;
  wire w6880;
  wire w6881;
  wire w6882;
  wire w6883;
  wire w6884;
  wire w6885;
  wire w6886;
  wire w6887;
  wire w6888;
  wire w6889;
  wire w6890;
  wire w6891;
  wire w6892;
  wire w6893;
  wire w6894;
  wire w6895;
  wire w6896;
  wire w6897;
  wire w6898;
  wire w6899;
  wire w6900;
  wire w6901;
  wire w6902;
  wire w6903;
  wire w6904;
  wire w6905;
  wire w6906;
  wire w6907;
  wire w6908;
  wire w6909;
  wire w6910;
  wire w6911;
  wire w6912;
  wire w6913;
  wire w6914;
  wire w6915;
  wire w6916;
  wire w6917;
  wire w6918;
  wire w6919;
  wire w6920;
  wire w6921;
  wire w6922;
  wire w6923;
  wire w6924;
  wire w6925;
  wire w6926;
  wire w6927;
  wire w6928;
  wire w6929;
  wire w6930;
  wire w6931;
  wire w6932;
  wire w6933;
  wire w6934;
  wire w6935;
  wire w6936;
  wire w6937;
  wire w6938;
  wire w6939;
  wire w6940;
  wire w6941;
  wire w6942;
  wire w6943;
  wire w6944;
  wire w6945;
  wire w6946;
  wire w6947;
  wire w6948;
  wire w6949;
  wire w6950;
  wire w6951;
  wire w6952;
  wire w6953;
  wire w6954;
  wire w6955;
  wire w6956;
  wire w6957;
  wire w6958;
  wire w6959;
  wire w6960;
  wire w6961;
  wire w6962;
  wire w6963;
  wire w6964;
  wire w6965;
  wire w6966;
  wire w6967;
  wire w6968;
  wire w6970;
  wire w6971;
  wire w6972;
  wire w6973;
  wire w6974;
  wire w6975;
  wire w6976;
  wire w6977;
  wire w6978;
  wire w6979;
  wire w6980;
  wire w6981;
  wire w6982;
  wire w6983;
  wire w6984;
  wire w6985;
  wire w6986;
  wire w6987;
  wire w6988;
  wire w6989;
  wire w6990;
  wire w6991;
  wire w6992;
  wire w6993;
  wire w6994;
  wire w6995;
  wire w6996;
  wire w6997;
  wire w6998;
  wire w6999;
  wire w7000;
  wire w7001;
  wire w7002;
  wire w7003;
  wire w7004;
  wire w7005;
  wire w7006;
  wire w7007;
  wire w7008;
  wire w7009;
  wire w7010;
  wire w7011;
  wire w7012;
  wire w7013;
  wire w7014;
  wire w7015;
  wire w7016;
  wire w7017;
  wire w7018;
  wire w7019;
  wire w7020;
  wire w7021;
  wire w7022;
  wire w7023;
  wire w7024;
  wire w7025;
  wire w7026;
  wire w7027;
  wire w7028;
  wire w7029;
  wire w7030;
  wire w7031;
  wire w7032;
  wire w7033;
  wire w7034;
  wire w7035;
  wire w7036;
  wire w7037;
  wire w7038;
  wire w7039;
  wire w7040;
  wire w7041;
  wire w7042;
  wire w7043;
  wire w7044;
  wire w7045;
  wire w7046;
  wire w7047;
  wire w7048;
  wire w7049;
  wire w7050;
  wire w7051;
  wire w7052;
  wire w7053;
  wire w7054;
  wire w7055;
  wire w7056;
  wire w7057;
  wire w7058;
  wire w7059;
  wire w7060;
  wire w7061;
  wire w7062;
  wire w7063;
  wire w7064;
  wire w7065;
  wire w7066;
  wire w7067;
  wire w7068;
  wire w7069;
  wire w7070;
  wire w7071;
  wire w7072;
  wire w7074;
  wire w7075;
  wire w7076;
  wire w7077;
  wire w7078;
  wire w7079;
  wire w7080;
  wire w7081;
  wire w7082;
  wire w7083;
  wire w7084;
  wire w7085;
  wire w7086;
  wire w7087;
  wire w7088;
  wire w7089;
  wire w7090;
  wire w7091;
  wire w7092;
  wire w7093;
  wire w7094;
  wire w7095;
  wire w7096;
  wire w7097;
  wire w7098;
  wire w7099;
  wire w7100;
  wire w7101;
  wire w7102;
  wire w7103;
  wire w7104;
  wire w7105;
  wire w7106;
  wire w7107;
  wire w7108;
  wire w7109;
  wire w7110;
  wire w7111;
  wire w7112;
  wire w7113;
  wire w7114;
  wire w7115;
  wire w7116;
  wire w7117;
  wire w7118;
  wire w7119;
  wire w7120;
  wire w7121;
  wire w7122;
  wire w7123;
  wire w7124;
  wire w7125;
  wire w7126;
  wire w7127;
  wire w7128;
  wire w7129;
  wire w7130;
  wire w7131;
  wire w7132;
  wire w7133;
  wire w7134;
  wire w7135;
  wire w7136;
  wire w7137;
  wire w7138;
  wire w7139;
  wire w7140;
  wire w7141;
  wire w7142;
  wire w7143;
  wire w7144;
  wire w7145;
  wire w7146;
  wire w7147;
  wire w7148;
  wire w7149;
  wire w7150;
  wire w7151;
  wire w7152;
  wire w7153;
  wire w7154;
  wire w7155;
  wire w7156;
  wire w7157;
  wire w7158;
  wire w7159;
  wire w7160;
  wire w7161;
  wire w7162;
  wire w7163;
  wire w7164;
  wire w7165;
  wire w7166;
  wire w7167;
  wire w7168;
  wire w7169;
  wire w7170;
  wire w7171;
  wire w7172;
  wire w7173;
  wire w7174;
  wire w7175;
  wire w7176;
  wire w7178;
  wire w7179;
  wire w7180;
  wire w7181;
  wire w7182;
  wire w7183;
  wire w7184;
  wire w7185;
  wire w7186;
  wire w7187;
  wire w7188;
  wire w7189;
  wire w7190;
  wire w7191;
  wire w7192;
  wire w7193;
  wire w7194;
  wire w7195;
  wire w7196;
  wire w7197;
  wire w7198;
  wire w7199;
  wire w7200;
  wire w7201;
  wire w7202;
  wire w7203;
  wire w7204;
  wire w7205;
  wire w7206;
  wire w7207;
  wire w7208;
  wire w7209;
  wire w7210;
  wire w7211;
  wire w7212;
  wire w7213;
  wire w7214;
  wire w7215;
  wire w7216;
  wire w7217;
  wire w7218;
  wire w7219;
  wire w7220;
  wire w7221;
  wire w7222;
  wire w7223;
  wire w7224;
  wire w7225;
  wire w7226;
  wire w7227;
  wire w7228;
  wire w7229;
  wire w7230;
  wire w7231;
  wire w7232;
  wire w7233;
  wire w7234;
  wire w7235;
  wire w7236;
  wire w7237;
  wire w7238;
  wire w7239;
  wire w7240;
  wire w7241;
  wire w7242;
  wire w7243;
  wire w7244;
  wire w7245;
  wire w7246;
  wire w7247;
  wire w7248;
  wire w7249;
  wire w7250;
  wire w7251;
  wire w7252;
  wire w7253;
  wire w7254;
  wire w7255;
  wire w7256;
  wire w7257;
  wire w7258;
  wire w7259;
  wire w7260;
  wire w7261;
  wire w7262;
  wire w7263;
  wire w7264;
  wire w7265;
  wire w7266;
  wire w7267;
  wire w7268;
  wire w7269;
  wire w7270;
  wire w7271;
  wire w7272;
  wire w7273;
  wire w7274;
  wire w7275;
  wire w7276;
  wire w7277;
  wire w7278;
  wire w7279;
  wire w7280;
  wire w7282;
  wire w7283;
  wire w7284;
  wire w7285;
  wire w7286;
  wire w7287;
  wire w7288;
  wire w7289;
  wire w7290;
  wire w7291;
  wire w7292;
  wire w7293;
  wire w7294;
  wire w7295;
  wire w7296;
  wire w7297;
  wire w7298;
  wire w7299;
  wire w7300;
  wire w7301;
  wire w7302;
  wire w7303;
  wire w7304;
  wire w7305;
  wire w7306;
  wire w7307;
  wire w7308;
  wire w7309;
  wire w7310;
  wire w7311;
  wire w7312;
  wire w7313;
  wire w7314;
  wire w7315;
  wire w7316;
  wire w7317;
  wire w7318;
  wire w7319;
  wire w7320;
  wire w7321;
  wire w7322;
  wire w7323;
  wire w7324;
  wire w7325;
  wire w7326;
  wire w7327;
  wire w7328;
  wire w7329;
  wire w7330;
  wire w7331;
  wire w7332;
  wire w7333;
  wire w7334;
  wire w7335;
  wire w7336;
  wire w7337;
  wire w7338;
  wire w7339;
  wire w7340;
  wire w7341;
  wire w7342;
  wire w7343;
  wire w7344;
  wire w7345;
  wire w7346;
  wire w7347;
  wire w7348;
  wire w7349;
  wire w7350;
  wire w7351;
  wire w7352;
  wire w7353;
  wire w7354;
  wire w7355;
  wire w7356;
  wire w7357;
  wire w7358;
  wire w7359;
  wire w7360;
  wire w7361;
  wire w7362;
  wire w7363;
  wire w7364;
  wire w7365;
  wire w7366;
  wire w7367;
  wire w7368;
  wire w7369;
  wire w7370;
  wire w7371;
  wire w7372;
  wire w7373;
  wire w7374;
  wire w7375;
  wire w7376;
  wire w7377;
  wire w7378;
  wire w7379;
  wire w7380;
  wire w7381;
  wire w7382;
  wire w7383;
  wire w7384;
  wire w7386;
  wire w7387;
  wire w7388;
  wire w7389;
  wire w7390;
  wire w7391;
  wire w7392;
  wire w7393;
  wire w7394;
  wire w7395;
  wire w7396;
  wire w7397;
  wire w7398;
  wire w7399;
  wire w7400;
  wire w7401;
  wire w7402;
  wire w7403;
  wire w7404;
  wire w7405;
  wire w7406;
  wire w7407;
  wire w7408;
  wire w7409;
  wire w7410;
  wire w7411;
  wire w7412;
  wire w7413;
  wire w7414;
  wire w7415;
  wire w7416;
  wire w7417;
  wire w7418;
  wire w7419;
  wire w7420;
  wire w7421;
  wire w7422;
  wire w7423;
  wire w7424;
  wire w7425;
  wire w7426;
  wire w7427;
  wire w7428;
  wire w7429;
  wire w7430;
  wire w7431;
  wire w7432;
  wire w7433;
  wire w7434;
  wire w7435;
  wire w7436;
  wire w7437;
  wire w7438;
  wire w7439;
  wire w7440;
  wire w7441;
  wire w7442;
  wire w7443;
  wire w7444;
  wire w7445;
  wire w7446;
  wire w7447;
  wire w7448;
  wire w7449;
  wire w7450;
  wire w7451;
  wire w7452;
  wire w7453;
  wire w7454;
  wire w7455;
  wire w7456;
  wire w7457;
  wire w7458;
  wire w7459;
  wire w7460;
  wire w7461;
  wire w7462;
  wire w7463;
  wire w7464;
  wire w7465;
  wire w7466;
  wire w7467;
  wire w7468;
  wire w7469;
  wire w7470;
  wire w7471;
  wire w7472;
  wire w7473;
  wire w7474;
  wire w7475;
  wire w7476;
  wire w7477;
  wire w7478;
  wire w7479;
  wire w7480;
  wire w7481;
  wire w7482;
  wire w7483;
  wire w7484;
  wire w7485;
  wire w7486;
  wire w7487;
  wire w7488;
  wire w7490;
  wire w7491;
  wire w7492;
  wire w7493;
  wire w7494;
  wire w7495;
  wire w7496;
  wire w7497;
  wire w7498;
  wire w7499;
  wire w7500;
  wire w7501;
  wire w7502;
  wire w7503;
  wire w7504;
  wire w7505;
  wire w7506;
  wire w7507;
  wire w7508;
  wire w7509;
  wire w7510;
  wire w7511;
  wire w7512;
  wire w7513;
  wire w7514;
  wire w7515;
  wire w7516;
  wire w7517;
  wire w7518;
  wire w7519;
  wire w7520;
  wire w7521;
  wire w7522;
  wire w7523;
  wire w7524;
  wire w7525;
  wire w7526;
  wire w7527;
  wire w7528;
  wire w7529;
  wire w7530;
  wire w7531;
  wire w7532;
  wire w7533;
  wire w7534;
  wire w7535;
  wire w7536;
  wire w7537;
  wire w7538;
  wire w7539;
  wire w7540;
  wire w7541;
  wire w7542;
  wire w7543;
  wire w7544;
  wire w7545;
  wire w7546;
  wire w7547;
  wire w7548;
  wire w7549;
  wire w7550;
  wire w7551;
  wire w7552;
  wire w7553;
  wire w7554;
  wire w7555;
  wire w7556;
  wire w7557;
  wire w7558;
  wire w7559;
  wire w7560;
  wire w7561;
  wire w7562;
  wire w7563;
  wire w7564;
  wire w7565;
  wire w7566;
  wire w7567;
  wire w7568;
  wire w7569;
  wire w7570;
  wire w7571;
  wire w7572;
  wire w7573;
  wire w7574;
  wire w7575;
  wire w7576;
  wire w7577;
  wire w7578;
  wire w7579;
  wire w7580;
  wire w7581;
  wire w7582;
  wire w7583;
  wire w7584;
  wire w7585;
  wire w7586;
  wire w7587;
  wire w7588;
  wire w7589;
  wire w7590;
  wire w7591;
  wire w7592;
  wire w7594;
  wire w7595;
  wire w7596;
  wire w7597;
  wire w7598;
  wire w7599;
  wire w7600;
  wire w7601;
  wire w7602;
  wire w7603;
  wire w7604;
  wire w7605;
  wire w7606;
  wire w7607;
  wire w7608;
  wire w7609;
  wire w7610;
  wire w7611;
  wire w7612;
  wire w7613;
  wire w7614;
  wire w7615;
  wire w7616;
  wire w7617;
  wire w7618;
  wire w7619;
  wire w7620;
  wire w7621;
  wire w7622;
  wire w7623;
  wire w7624;
  wire w7625;
  wire w7626;
  wire w7627;
  wire w7628;
  wire w7629;
  wire w7630;
  wire w7631;
  wire w7632;
  wire w7633;
  wire w7634;
  wire w7635;
  wire w7636;
  wire w7637;
  wire w7638;
  wire w7639;
  wire w7640;
  wire w7641;
  wire w7642;
  wire w7643;
  wire w7644;
  wire w7645;
  wire w7646;
  wire w7647;
  wire w7648;
  wire w7649;
  wire w7650;
  wire w7651;
  wire w7652;
  wire w7653;
  wire w7654;
  wire w7655;
  wire w7656;
  wire w7657;
  wire w7658;
  wire w7659;
  wire w7660;
  wire w7661;
  wire w7662;
  wire w7663;
  wire w7664;
  wire w7665;
  wire w7666;
  wire w7667;
  wire w7668;
  wire w7669;
  wire w7670;
  wire w7671;
  wire w7672;
  wire w7673;
  wire w7674;
  wire w7675;
  wire w7676;
  wire w7677;
  wire w7678;
  wire w7679;
  wire w7680;
  wire w7681;
  wire w7682;
  wire w7683;
  wire w7684;
  wire w7685;
  wire w7686;
  wire w7687;
  wire w7688;
  wire w7689;
  wire w7690;
  wire w7691;
  wire w7692;
  wire w7693;
  wire w7694;
  wire w7695;
  wire w7696;
  wire w7698;
  wire w7699;
  wire w7700;
  wire w7701;
  wire w7702;
  wire w7703;
  wire w7704;
  wire w7705;
  wire w7706;
  wire w7707;
  wire w7708;
  wire w7709;
  wire w7710;
  wire w7711;
  wire w7712;
  wire w7713;
  wire w7714;
  wire w7715;
  wire w7716;
  wire w7717;
  wire w7718;
  wire w7719;
  wire w7720;
  wire w7721;
  wire w7722;
  wire w7723;
  wire w7724;
  wire w7725;
  wire w7726;
  wire w7727;
  wire w7728;
  wire w7729;
  wire w7730;
  wire w7731;
  wire w7732;
  wire w7733;
  wire w7734;
  wire w7735;
  wire w7736;
  wire w7737;
  wire w7738;
  wire w7739;
  wire w7740;
  wire w7741;
  wire w7742;
  wire w7743;
  wire w7744;
  wire w7745;
  wire w7746;
  wire w7747;
  wire w7748;
  wire w7749;
  wire w7750;
  wire w7751;
  wire w7752;
  wire w7753;
  wire w7754;
  wire w7755;
  wire w7756;
  wire w7757;
  wire w7758;
  wire w7759;
  wire w7760;
  wire w7761;
  wire w7762;
  wire w7763;
  wire w7764;
  wire w7765;
  wire w7766;
  wire w7767;
  wire w7768;
  wire w7769;
  wire w7770;
  wire w7771;
  wire w7772;
  wire w7773;
  wire w7774;
  wire w7775;
  wire w7776;
  wire w7777;
  wire w7778;
  wire w7779;
  wire w7780;
  wire w7781;
  wire w7782;
  wire w7783;
  wire w7784;
  wire w7785;
  wire w7786;
  wire w7787;
  wire w7788;
  wire w7789;
  wire w7790;
  wire w7791;
  wire w7792;
  wire w7793;
  wire w7794;
  wire w7795;
  wire w7796;
  wire w7797;
  wire w7798;
  wire w7799;
  wire w7800;
  wire w7802;
  wire w7803;
  wire w7804;
  wire w7805;
  wire w7806;
  wire w7807;
  wire w7808;
  wire w7809;
  wire w7810;
  wire w7811;
  wire w7812;
  wire w7813;
  wire w7814;
  wire w7815;
  wire w7816;
  wire w7817;
  wire w7818;
  wire w7819;
  wire w7820;
  wire w7821;
  wire w7822;
  wire w7823;
  wire w7824;
  wire w7825;
  wire w7826;
  wire w7827;
  wire w7828;
  wire w7829;
  wire w7830;
  wire w7831;
  wire w7832;
  wire w7833;
  wire w7834;
  wire w7835;
  wire w7836;
  wire w7837;
  wire w7838;
  wire w7839;
  wire w7840;
  wire w7841;
  wire w7842;
  wire w7843;
  wire w7844;
  wire w7845;
  wire w7846;
  wire w7847;
  wire w7848;
  wire w7849;
  wire w7850;
  wire w7851;
  wire w7852;
  wire w7853;
  wire w7854;
  wire w7855;
  wire w7856;
  wire w7857;
  wire w7858;
  wire w7859;
  wire w7860;
  wire w7861;
  wire w7862;
  wire w7863;
  wire w7864;
  wire w7865;
  wire w7866;
  wire w7867;
  wire w7868;
  wire w7869;
  wire w7870;
  wire w7871;
  wire w7872;
  wire w7873;
  wire w7874;
  wire w7875;
  wire w7876;
  wire w7877;
  wire w7878;
  wire w7879;
  wire w7880;
  wire w7881;
  wire w7882;
  wire w7883;
  wire w7884;
  wire w7885;
  wire w7886;
  wire w7887;
  wire w7888;
  wire w7889;
  wire w7890;
  wire w7891;
  wire w7892;
  wire w7893;
  wire w7894;
  wire w7895;
  wire w7896;
  wire w7897;
  wire w7898;
  wire w7899;
  wire w7900;
  wire w7901;
  wire w7902;
  wire w7903;
  wire w7904;
  wire w7906;
  wire w7907;
  wire w7908;
  wire w7909;
  wire w7910;
  wire w7911;
  wire w7912;
  wire w7913;
  wire w7914;
  wire w7915;
  wire w7916;
  wire w7917;
  wire w7918;
  wire w7919;
  wire w7920;
  wire w7921;
  wire w7922;
  wire w7923;
  wire w7924;
  wire w7925;
  wire w7926;
  wire w7927;
  wire w7928;
  wire w7929;
  wire w7930;
  wire w7931;
  wire w7932;
  wire w7933;
  wire w7934;
  wire w7935;
  wire w7936;
  wire w7937;
  wire w7938;
  wire w7939;
  wire w7940;
  wire w7941;
  wire w7942;
  wire w7943;
  wire w7944;
  wire w7945;
  wire w7946;
  wire w7947;
  wire w7948;
  wire w7949;
  wire w7950;
  wire w7951;
  wire w7952;
  wire w7953;
  wire w7954;
  wire w7955;
  wire w7956;
  wire w7957;
  wire w7958;
  wire w7959;
  wire w7960;
  wire w7961;
  wire w7962;
  wire w7963;
  wire w7964;
  wire w7965;
  wire w7966;
  wire w7967;
  wire w7968;
  wire w7969;
  wire w7970;
  wire w7971;
  wire w7972;
  wire w7973;
  wire w7974;
  wire w7975;
  wire w7976;
  wire w7977;
  wire w7978;
  wire w7979;
  wire w7980;
  wire w7981;
  wire w7982;
  wire w7983;
  wire w7984;
  wire w7985;
  wire w7986;
  wire w7987;
  wire w7988;
  wire w7989;
  wire w7990;
  wire w7991;
  wire w7992;
  wire w7993;
  wire w7994;
  wire w7995;
  wire w7996;
  wire w7997;
  wire w7998;
  wire w7999;
  wire w8000;
  wire w8001;
  wire w8002;
  wire w8003;
  wire w8004;
  wire w8005;
  wire w8006;
  wire w8007;
  wire w8008;
  wire w8010;
  wire w8011;
  wire w8012;
  wire w8013;
  wire w8014;
  wire w8015;
  wire w8016;
  wire w8017;
  wire w8018;
  wire w8019;
  wire w8020;
  wire w8021;
  wire w8022;
  wire w8023;
  wire w8024;
  wire w8025;
  wire w8026;
  wire w8027;
  wire w8028;
  wire w8029;
  wire w8030;
  wire w8031;
  wire w8032;
  wire w8033;
  wire w8034;
  wire w8035;
  wire w8036;
  wire w8037;
  wire w8038;
  wire w8039;
  wire w8040;
  wire w8041;
  wire w8042;
  wire w8043;
  wire w8044;
  wire w8045;
  wire w8046;
  wire w8047;
  wire w8048;
  wire w8049;
  wire w8050;
  wire w8051;
  wire w8052;
  wire w8053;
  wire w8054;
  wire w8055;
  wire w8056;
  wire w8057;
  wire w8058;
  wire w8059;
  wire w8060;
  wire w8061;
  wire w8062;
  wire w8063;
  wire w8064;
  wire w8065;
  wire w8066;
  wire w8067;
  wire w8068;
  wire w8069;
  wire w8070;
  wire w8071;
  wire w8072;
  wire w8073;
  wire w8074;
  wire w8075;
  wire w8076;
  wire w8077;
  wire w8078;
  wire w8079;
  wire w8080;
  wire w8081;
  wire w8082;
  wire w8083;
  wire w8084;
  wire w8085;
  wire w8086;
  wire w8087;
  wire w8088;
  wire w8089;
  wire w8090;
  wire w8091;
  wire w8092;
  wire w8093;
  wire w8094;
  wire w8095;
  wire w8096;
  wire w8097;
  wire w8098;
  wire w8099;
  wire w8100;
  wire w8101;
  wire w8102;
  wire w8103;
  wire w8104;
  wire w8105;
  wire w8106;
  wire w8107;
  wire w8108;
  wire w8109;
  wire w8110;
  wire w8111;
  wire w8112;
  wire w8114;
  wire w8116;
  wire w8118;
  wire w8120;
  wire w8122;
  wire w8124;
  wire w8126;
  wire w8128;
  wire w8130;
  wire w8132;
  wire w8134;
  wire w8136;
  wire w8138;
  wire w8140;
  wire w8142;
  wire w8144;
  wire w8146;
  wire w8148;
  wire w8150;
  wire w8152;
  wire w8154;
  wire w8156;
  wire w8158;
  wire w8160;
  wire w8162;
  wire w8164;
  wire w8166;
  wire w8168;
  wire w8170;
  wire w8172;
  wire w8174;
  wire w8176;
  wire w8178;
  wire w8180;
  wire w8182;
  wire w8184;
  wire w8186;
  wire w8188;
  wire w8190;
  wire w8192;
  wire w8194;
  wire w8196;
  wire w8198;
  wire w8200;
  wire w8202;
  wire w8204;
  wire w8206;
  wire w8208;
  wire w8210;
  wire w8212;
  wire w8214;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w2810);
  FullAdder U1 (w2810, IN2[0], IN2[1], w2811, w2812);
  FullAdder U2 (w2812, IN3[0], IN3[1], w2813, w2814);
  FullAdder U3 (w2814, IN4[0], IN4[1], w2815, w2816);
  FullAdder U4 (w2816, IN5[0], IN5[1], w2817, w2818);
  FullAdder U5 (w2818, IN6[0], IN6[1], w2819, w2820);
  FullAdder U6 (w2820, IN7[0], IN7[1], w2821, w2822);
  FullAdder U7 (w2822, IN8[0], IN8[1], w2823, w2824);
  FullAdder U8 (w2824, IN9[0], IN9[1], w2825, w2826);
  FullAdder U9 (w2826, IN10[0], IN10[1], w2827, w2828);
  FullAdder U10 (w2828, IN11[0], IN11[1], w2829, w2830);
  FullAdder U11 (w2830, IN12[0], IN12[1], w2831, w2832);
  FullAdder U12 (w2832, IN13[0], IN13[1], w2833, w2834);
  FullAdder U13 (w2834, IN14[0], IN14[1], w2835, w2836);
  FullAdder U14 (w2836, IN15[0], IN15[1], w2837, w2838);
  FullAdder U15 (w2838, IN16[0], IN16[1], w2839, w2840);
  FullAdder U16 (w2840, IN17[0], IN17[1], w2841, w2842);
  FullAdder U17 (w2842, IN18[0], IN18[1], w2843, w2844);
  FullAdder U18 (w2844, IN19[0], IN19[1], w2845, w2846);
  FullAdder U19 (w2846, IN20[0], IN20[1], w2847, w2848);
  FullAdder U20 (w2848, IN21[0], IN21[1], w2849, w2850);
  FullAdder U21 (w2850, IN22[0], IN22[1], w2851, w2852);
  FullAdder U22 (w2852, IN23[0], IN23[1], w2853, w2854);
  FullAdder U23 (w2854, IN24[0], IN24[1], w2855, w2856);
  FullAdder U24 (w2856, IN25[0], IN25[1], w2857, w2858);
  FullAdder U25 (w2858, IN26[0], IN26[1], w2859, w2860);
  FullAdder U26 (w2860, IN27[0], IN27[1], w2861, w2862);
  FullAdder U27 (w2862, IN28[0], IN28[1], w2863, w2864);
  FullAdder U28 (w2864, IN29[0], IN29[1], w2865, w2866);
  FullAdder U29 (w2866, IN30[0], IN30[1], w2867, w2868);
  FullAdder U30 (w2868, IN31[0], IN31[1], w2869, w2870);
  FullAdder U31 (w2870, IN32[0], IN32[1], w2871, w2872);
  FullAdder U32 (w2872, IN33[0], IN33[1], w2873, w2874);
  FullAdder U33 (w2874, IN34[0], IN34[1], w2875, w2876);
  FullAdder U34 (w2876, IN35[0], IN35[1], w2877, w2878);
  FullAdder U35 (w2878, IN36[0], IN36[1], w2879, w2880);
  FullAdder U36 (w2880, IN37[0], IN37[1], w2881, w2882);
  FullAdder U37 (w2882, IN38[0], IN38[1], w2883, w2884);
  FullAdder U38 (w2884, IN39[0], IN39[1], w2885, w2886);
  FullAdder U39 (w2886, IN40[0], IN40[1], w2887, w2888);
  FullAdder U40 (w2888, IN41[0], IN41[1], w2889, w2890);
  FullAdder U41 (w2890, IN42[0], IN42[1], w2891, w2892);
  FullAdder U42 (w2892, IN43[0], IN43[1], w2893, w2894);
  FullAdder U43 (w2894, IN44[0], IN44[1], w2895, w2896);
  FullAdder U44 (w2896, IN45[0], IN45[1], w2897, w2898);
  FullAdder U45 (w2898, IN46[0], IN46[1], w2899, w2900);
  FullAdder U46 (w2900, IN47[0], IN47[1], w2901, w2902);
  FullAdder U47 (w2902, IN48[0], IN48[1], w2903, w2904);
  FullAdder U48 (w2904, IN49[0], IN49[1], w2905, w2906);
  FullAdder U49 (w2906, IN50[0], IN50[1], w2907, w2908);
  FullAdder U50 (w2908, IN51[0], IN51[1], w2909, w2910);
  FullAdder U51 (w2910, IN52[0], IN52[1], w2911, w2912);
  HalfAdder U52 (w2811, IN2[2], Out1[2], w2914);
  FullAdder U53 (w2914, w2813, IN3[2], w2915, w2916);
  FullAdder U54 (w2916, w2815, IN4[2], w2917, w2918);
  FullAdder U55 (w2918, w2817, IN5[2], w2919, w2920);
  FullAdder U56 (w2920, w2819, IN6[2], w2921, w2922);
  FullAdder U57 (w2922, w2821, IN7[2], w2923, w2924);
  FullAdder U58 (w2924, w2823, IN8[2], w2925, w2926);
  FullAdder U59 (w2926, w2825, IN9[2], w2927, w2928);
  FullAdder U60 (w2928, w2827, IN10[2], w2929, w2930);
  FullAdder U61 (w2930, w2829, IN11[2], w2931, w2932);
  FullAdder U62 (w2932, w2831, IN12[2], w2933, w2934);
  FullAdder U63 (w2934, w2833, IN13[2], w2935, w2936);
  FullAdder U64 (w2936, w2835, IN14[2], w2937, w2938);
  FullAdder U65 (w2938, w2837, IN15[2], w2939, w2940);
  FullAdder U66 (w2940, w2839, IN16[2], w2941, w2942);
  FullAdder U67 (w2942, w2841, IN17[2], w2943, w2944);
  FullAdder U68 (w2944, w2843, IN18[2], w2945, w2946);
  FullAdder U69 (w2946, w2845, IN19[2], w2947, w2948);
  FullAdder U70 (w2948, w2847, IN20[2], w2949, w2950);
  FullAdder U71 (w2950, w2849, IN21[2], w2951, w2952);
  FullAdder U72 (w2952, w2851, IN22[2], w2953, w2954);
  FullAdder U73 (w2954, w2853, IN23[2], w2955, w2956);
  FullAdder U74 (w2956, w2855, IN24[2], w2957, w2958);
  FullAdder U75 (w2958, w2857, IN25[2], w2959, w2960);
  FullAdder U76 (w2960, w2859, IN26[2], w2961, w2962);
  FullAdder U77 (w2962, w2861, IN27[2], w2963, w2964);
  FullAdder U78 (w2964, w2863, IN28[2], w2965, w2966);
  FullAdder U79 (w2966, w2865, IN29[2], w2967, w2968);
  FullAdder U80 (w2968, w2867, IN30[2], w2969, w2970);
  FullAdder U81 (w2970, w2869, IN31[2], w2971, w2972);
  FullAdder U82 (w2972, w2871, IN32[2], w2973, w2974);
  FullAdder U83 (w2974, w2873, IN33[2], w2975, w2976);
  FullAdder U84 (w2976, w2875, IN34[2], w2977, w2978);
  FullAdder U85 (w2978, w2877, IN35[2], w2979, w2980);
  FullAdder U86 (w2980, w2879, IN36[2], w2981, w2982);
  FullAdder U87 (w2982, w2881, IN37[2], w2983, w2984);
  FullAdder U88 (w2984, w2883, IN38[2], w2985, w2986);
  FullAdder U89 (w2986, w2885, IN39[2], w2987, w2988);
  FullAdder U90 (w2988, w2887, IN40[2], w2989, w2990);
  FullAdder U91 (w2990, w2889, IN41[2], w2991, w2992);
  FullAdder U92 (w2992, w2891, IN42[2], w2993, w2994);
  FullAdder U93 (w2994, w2893, IN43[2], w2995, w2996);
  FullAdder U94 (w2996, w2895, IN44[2], w2997, w2998);
  FullAdder U95 (w2998, w2897, IN45[2], w2999, w3000);
  FullAdder U96 (w3000, w2899, IN46[2], w3001, w3002);
  FullAdder U97 (w3002, w2901, IN47[2], w3003, w3004);
  FullAdder U98 (w3004, w2903, IN48[2], w3005, w3006);
  FullAdder U99 (w3006, w2905, IN49[2], w3007, w3008);
  FullAdder U100 (w3008, w2907, IN50[2], w3009, w3010);
  FullAdder U101 (w3010, w2909, IN51[2], w3011, w3012);
  FullAdder U102 (w3012, w2911, IN52[2], w3013, w3014);
  FullAdder U103 (w3014, w2912, IN53[0], w3015, w3016);
  HalfAdder U104 (w2915, IN3[3], Out1[3], w3018);
  FullAdder U105 (w3018, w2917, IN4[3], w3019, w3020);
  FullAdder U106 (w3020, w2919, IN5[3], w3021, w3022);
  FullAdder U107 (w3022, w2921, IN6[3], w3023, w3024);
  FullAdder U108 (w3024, w2923, IN7[3], w3025, w3026);
  FullAdder U109 (w3026, w2925, IN8[3], w3027, w3028);
  FullAdder U110 (w3028, w2927, IN9[3], w3029, w3030);
  FullAdder U111 (w3030, w2929, IN10[3], w3031, w3032);
  FullAdder U112 (w3032, w2931, IN11[3], w3033, w3034);
  FullAdder U113 (w3034, w2933, IN12[3], w3035, w3036);
  FullAdder U114 (w3036, w2935, IN13[3], w3037, w3038);
  FullAdder U115 (w3038, w2937, IN14[3], w3039, w3040);
  FullAdder U116 (w3040, w2939, IN15[3], w3041, w3042);
  FullAdder U117 (w3042, w2941, IN16[3], w3043, w3044);
  FullAdder U118 (w3044, w2943, IN17[3], w3045, w3046);
  FullAdder U119 (w3046, w2945, IN18[3], w3047, w3048);
  FullAdder U120 (w3048, w2947, IN19[3], w3049, w3050);
  FullAdder U121 (w3050, w2949, IN20[3], w3051, w3052);
  FullAdder U122 (w3052, w2951, IN21[3], w3053, w3054);
  FullAdder U123 (w3054, w2953, IN22[3], w3055, w3056);
  FullAdder U124 (w3056, w2955, IN23[3], w3057, w3058);
  FullAdder U125 (w3058, w2957, IN24[3], w3059, w3060);
  FullAdder U126 (w3060, w2959, IN25[3], w3061, w3062);
  FullAdder U127 (w3062, w2961, IN26[3], w3063, w3064);
  FullAdder U128 (w3064, w2963, IN27[3], w3065, w3066);
  FullAdder U129 (w3066, w2965, IN28[3], w3067, w3068);
  FullAdder U130 (w3068, w2967, IN29[3], w3069, w3070);
  FullAdder U131 (w3070, w2969, IN30[3], w3071, w3072);
  FullAdder U132 (w3072, w2971, IN31[3], w3073, w3074);
  FullAdder U133 (w3074, w2973, IN32[3], w3075, w3076);
  FullAdder U134 (w3076, w2975, IN33[3], w3077, w3078);
  FullAdder U135 (w3078, w2977, IN34[3], w3079, w3080);
  FullAdder U136 (w3080, w2979, IN35[3], w3081, w3082);
  FullAdder U137 (w3082, w2981, IN36[3], w3083, w3084);
  FullAdder U138 (w3084, w2983, IN37[3], w3085, w3086);
  FullAdder U139 (w3086, w2985, IN38[3], w3087, w3088);
  FullAdder U140 (w3088, w2987, IN39[3], w3089, w3090);
  FullAdder U141 (w3090, w2989, IN40[3], w3091, w3092);
  FullAdder U142 (w3092, w2991, IN41[3], w3093, w3094);
  FullAdder U143 (w3094, w2993, IN42[3], w3095, w3096);
  FullAdder U144 (w3096, w2995, IN43[3], w3097, w3098);
  FullAdder U145 (w3098, w2997, IN44[3], w3099, w3100);
  FullAdder U146 (w3100, w2999, IN45[3], w3101, w3102);
  FullAdder U147 (w3102, w3001, IN46[3], w3103, w3104);
  FullAdder U148 (w3104, w3003, IN47[3], w3105, w3106);
  FullAdder U149 (w3106, w3005, IN48[3], w3107, w3108);
  FullAdder U150 (w3108, w3007, IN49[3], w3109, w3110);
  FullAdder U151 (w3110, w3009, IN50[3], w3111, w3112);
  FullAdder U152 (w3112, w3011, IN51[3], w3113, w3114);
  FullAdder U153 (w3114, w3013, IN52[3], w3115, w3116);
  FullAdder U154 (w3116, w3015, IN53[1], w3117, w3118);
  FullAdder U155 (w3118, w3016, IN54[0], w3119, w3120);
  HalfAdder U156 (w3019, IN4[4], Out1[4], w3122);
  FullAdder U157 (w3122, w3021, IN5[4], w3123, w3124);
  FullAdder U158 (w3124, w3023, IN6[4], w3125, w3126);
  FullAdder U159 (w3126, w3025, IN7[4], w3127, w3128);
  FullAdder U160 (w3128, w3027, IN8[4], w3129, w3130);
  FullAdder U161 (w3130, w3029, IN9[4], w3131, w3132);
  FullAdder U162 (w3132, w3031, IN10[4], w3133, w3134);
  FullAdder U163 (w3134, w3033, IN11[4], w3135, w3136);
  FullAdder U164 (w3136, w3035, IN12[4], w3137, w3138);
  FullAdder U165 (w3138, w3037, IN13[4], w3139, w3140);
  FullAdder U166 (w3140, w3039, IN14[4], w3141, w3142);
  FullAdder U167 (w3142, w3041, IN15[4], w3143, w3144);
  FullAdder U168 (w3144, w3043, IN16[4], w3145, w3146);
  FullAdder U169 (w3146, w3045, IN17[4], w3147, w3148);
  FullAdder U170 (w3148, w3047, IN18[4], w3149, w3150);
  FullAdder U171 (w3150, w3049, IN19[4], w3151, w3152);
  FullAdder U172 (w3152, w3051, IN20[4], w3153, w3154);
  FullAdder U173 (w3154, w3053, IN21[4], w3155, w3156);
  FullAdder U174 (w3156, w3055, IN22[4], w3157, w3158);
  FullAdder U175 (w3158, w3057, IN23[4], w3159, w3160);
  FullAdder U176 (w3160, w3059, IN24[4], w3161, w3162);
  FullAdder U177 (w3162, w3061, IN25[4], w3163, w3164);
  FullAdder U178 (w3164, w3063, IN26[4], w3165, w3166);
  FullAdder U179 (w3166, w3065, IN27[4], w3167, w3168);
  FullAdder U180 (w3168, w3067, IN28[4], w3169, w3170);
  FullAdder U181 (w3170, w3069, IN29[4], w3171, w3172);
  FullAdder U182 (w3172, w3071, IN30[4], w3173, w3174);
  FullAdder U183 (w3174, w3073, IN31[4], w3175, w3176);
  FullAdder U184 (w3176, w3075, IN32[4], w3177, w3178);
  FullAdder U185 (w3178, w3077, IN33[4], w3179, w3180);
  FullAdder U186 (w3180, w3079, IN34[4], w3181, w3182);
  FullAdder U187 (w3182, w3081, IN35[4], w3183, w3184);
  FullAdder U188 (w3184, w3083, IN36[4], w3185, w3186);
  FullAdder U189 (w3186, w3085, IN37[4], w3187, w3188);
  FullAdder U190 (w3188, w3087, IN38[4], w3189, w3190);
  FullAdder U191 (w3190, w3089, IN39[4], w3191, w3192);
  FullAdder U192 (w3192, w3091, IN40[4], w3193, w3194);
  FullAdder U193 (w3194, w3093, IN41[4], w3195, w3196);
  FullAdder U194 (w3196, w3095, IN42[4], w3197, w3198);
  FullAdder U195 (w3198, w3097, IN43[4], w3199, w3200);
  FullAdder U196 (w3200, w3099, IN44[4], w3201, w3202);
  FullAdder U197 (w3202, w3101, IN45[4], w3203, w3204);
  FullAdder U198 (w3204, w3103, IN46[4], w3205, w3206);
  FullAdder U199 (w3206, w3105, IN47[4], w3207, w3208);
  FullAdder U200 (w3208, w3107, IN48[4], w3209, w3210);
  FullAdder U201 (w3210, w3109, IN49[4], w3211, w3212);
  FullAdder U202 (w3212, w3111, IN50[4], w3213, w3214);
  FullAdder U203 (w3214, w3113, IN51[4], w3215, w3216);
  FullAdder U204 (w3216, w3115, IN52[4], w3217, w3218);
  FullAdder U205 (w3218, w3117, IN53[2], w3219, w3220);
  FullAdder U206 (w3220, w3119, IN54[1], w3221, w3222);
  FullAdder U207 (w3222, w3120, IN55[0], w3223, w3224);
  HalfAdder U208 (w3123, IN5[5], Out1[5], w3226);
  FullAdder U209 (w3226, w3125, IN6[5], w3227, w3228);
  FullAdder U210 (w3228, w3127, IN7[5], w3229, w3230);
  FullAdder U211 (w3230, w3129, IN8[5], w3231, w3232);
  FullAdder U212 (w3232, w3131, IN9[5], w3233, w3234);
  FullAdder U213 (w3234, w3133, IN10[5], w3235, w3236);
  FullAdder U214 (w3236, w3135, IN11[5], w3237, w3238);
  FullAdder U215 (w3238, w3137, IN12[5], w3239, w3240);
  FullAdder U216 (w3240, w3139, IN13[5], w3241, w3242);
  FullAdder U217 (w3242, w3141, IN14[5], w3243, w3244);
  FullAdder U218 (w3244, w3143, IN15[5], w3245, w3246);
  FullAdder U219 (w3246, w3145, IN16[5], w3247, w3248);
  FullAdder U220 (w3248, w3147, IN17[5], w3249, w3250);
  FullAdder U221 (w3250, w3149, IN18[5], w3251, w3252);
  FullAdder U222 (w3252, w3151, IN19[5], w3253, w3254);
  FullAdder U223 (w3254, w3153, IN20[5], w3255, w3256);
  FullAdder U224 (w3256, w3155, IN21[5], w3257, w3258);
  FullAdder U225 (w3258, w3157, IN22[5], w3259, w3260);
  FullAdder U226 (w3260, w3159, IN23[5], w3261, w3262);
  FullAdder U227 (w3262, w3161, IN24[5], w3263, w3264);
  FullAdder U228 (w3264, w3163, IN25[5], w3265, w3266);
  FullAdder U229 (w3266, w3165, IN26[5], w3267, w3268);
  FullAdder U230 (w3268, w3167, IN27[5], w3269, w3270);
  FullAdder U231 (w3270, w3169, IN28[5], w3271, w3272);
  FullAdder U232 (w3272, w3171, IN29[5], w3273, w3274);
  FullAdder U233 (w3274, w3173, IN30[5], w3275, w3276);
  FullAdder U234 (w3276, w3175, IN31[5], w3277, w3278);
  FullAdder U235 (w3278, w3177, IN32[5], w3279, w3280);
  FullAdder U236 (w3280, w3179, IN33[5], w3281, w3282);
  FullAdder U237 (w3282, w3181, IN34[5], w3283, w3284);
  FullAdder U238 (w3284, w3183, IN35[5], w3285, w3286);
  FullAdder U239 (w3286, w3185, IN36[5], w3287, w3288);
  FullAdder U240 (w3288, w3187, IN37[5], w3289, w3290);
  FullAdder U241 (w3290, w3189, IN38[5], w3291, w3292);
  FullAdder U242 (w3292, w3191, IN39[5], w3293, w3294);
  FullAdder U243 (w3294, w3193, IN40[5], w3295, w3296);
  FullAdder U244 (w3296, w3195, IN41[5], w3297, w3298);
  FullAdder U245 (w3298, w3197, IN42[5], w3299, w3300);
  FullAdder U246 (w3300, w3199, IN43[5], w3301, w3302);
  FullAdder U247 (w3302, w3201, IN44[5], w3303, w3304);
  FullAdder U248 (w3304, w3203, IN45[5], w3305, w3306);
  FullAdder U249 (w3306, w3205, IN46[5], w3307, w3308);
  FullAdder U250 (w3308, w3207, IN47[5], w3309, w3310);
  FullAdder U251 (w3310, w3209, IN48[5], w3311, w3312);
  FullAdder U252 (w3312, w3211, IN49[5], w3313, w3314);
  FullAdder U253 (w3314, w3213, IN50[5], w3315, w3316);
  FullAdder U254 (w3316, w3215, IN51[5], w3317, w3318);
  FullAdder U255 (w3318, w3217, IN52[5], w3319, w3320);
  FullAdder U256 (w3320, w3219, IN53[3], w3321, w3322);
  FullAdder U257 (w3322, w3221, IN54[2], w3323, w3324);
  FullAdder U258 (w3324, w3223, IN55[1], w3325, w3326);
  FullAdder U259 (w3326, w3224, IN56[0], w3327, w3328);
  HalfAdder U260 (w3227, IN6[6], Out1[6], w3330);
  FullAdder U261 (w3330, w3229, IN7[6], w3331, w3332);
  FullAdder U262 (w3332, w3231, IN8[6], w3333, w3334);
  FullAdder U263 (w3334, w3233, IN9[6], w3335, w3336);
  FullAdder U264 (w3336, w3235, IN10[6], w3337, w3338);
  FullAdder U265 (w3338, w3237, IN11[6], w3339, w3340);
  FullAdder U266 (w3340, w3239, IN12[6], w3341, w3342);
  FullAdder U267 (w3342, w3241, IN13[6], w3343, w3344);
  FullAdder U268 (w3344, w3243, IN14[6], w3345, w3346);
  FullAdder U269 (w3346, w3245, IN15[6], w3347, w3348);
  FullAdder U270 (w3348, w3247, IN16[6], w3349, w3350);
  FullAdder U271 (w3350, w3249, IN17[6], w3351, w3352);
  FullAdder U272 (w3352, w3251, IN18[6], w3353, w3354);
  FullAdder U273 (w3354, w3253, IN19[6], w3355, w3356);
  FullAdder U274 (w3356, w3255, IN20[6], w3357, w3358);
  FullAdder U275 (w3358, w3257, IN21[6], w3359, w3360);
  FullAdder U276 (w3360, w3259, IN22[6], w3361, w3362);
  FullAdder U277 (w3362, w3261, IN23[6], w3363, w3364);
  FullAdder U278 (w3364, w3263, IN24[6], w3365, w3366);
  FullAdder U279 (w3366, w3265, IN25[6], w3367, w3368);
  FullAdder U280 (w3368, w3267, IN26[6], w3369, w3370);
  FullAdder U281 (w3370, w3269, IN27[6], w3371, w3372);
  FullAdder U282 (w3372, w3271, IN28[6], w3373, w3374);
  FullAdder U283 (w3374, w3273, IN29[6], w3375, w3376);
  FullAdder U284 (w3376, w3275, IN30[6], w3377, w3378);
  FullAdder U285 (w3378, w3277, IN31[6], w3379, w3380);
  FullAdder U286 (w3380, w3279, IN32[6], w3381, w3382);
  FullAdder U287 (w3382, w3281, IN33[6], w3383, w3384);
  FullAdder U288 (w3384, w3283, IN34[6], w3385, w3386);
  FullAdder U289 (w3386, w3285, IN35[6], w3387, w3388);
  FullAdder U290 (w3388, w3287, IN36[6], w3389, w3390);
  FullAdder U291 (w3390, w3289, IN37[6], w3391, w3392);
  FullAdder U292 (w3392, w3291, IN38[6], w3393, w3394);
  FullAdder U293 (w3394, w3293, IN39[6], w3395, w3396);
  FullAdder U294 (w3396, w3295, IN40[6], w3397, w3398);
  FullAdder U295 (w3398, w3297, IN41[6], w3399, w3400);
  FullAdder U296 (w3400, w3299, IN42[6], w3401, w3402);
  FullAdder U297 (w3402, w3301, IN43[6], w3403, w3404);
  FullAdder U298 (w3404, w3303, IN44[6], w3405, w3406);
  FullAdder U299 (w3406, w3305, IN45[6], w3407, w3408);
  FullAdder U300 (w3408, w3307, IN46[6], w3409, w3410);
  FullAdder U301 (w3410, w3309, IN47[6], w3411, w3412);
  FullAdder U302 (w3412, w3311, IN48[6], w3413, w3414);
  FullAdder U303 (w3414, w3313, IN49[6], w3415, w3416);
  FullAdder U304 (w3416, w3315, IN50[6], w3417, w3418);
  FullAdder U305 (w3418, w3317, IN51[6], w3419, w3420);
  FullAdder U306 (w3420, w3319, IN52[6], w3421, w3422);
  FullAdder U307 (w3422, w3321, IN53[4], w3423, w3424);
  FullAdder U308 (w3424, w3323, IN54[3], w3425, w3426);
  FullAdder U309 (w3426, w3325, IN55[2], w3427, w3428);
  FullAdder U310 (w3428, w3327, IN56[1], w3429, w3430);
  FullAdder U311 (w3430, w3328, IN57[0], w3431, w3432);
  HalfAdder U312 (w3331, IN7[7], Out1[7], w3434);
  FullAdder U313 (w3434, w3333, IN8[7], w3435, w3436);
  FullAdder U314 (w3436, w3335, IN9[7], w3437, w3438);
  FullAdder U315 (w3438, w3337, IN10[7], w3439, w3440);
  FullAdder U316 (w3440, w3339, IN11[7], w3441, w3442);
  FullAdder U317 (w3442, w3341, IN12[7], w3443, w3444);
  FullAdder U318 (w3444, w3343, IN13[7], w3445, w3446);
  FullAdder U319 (w3446, w3345, IN14[7], w3447, w3448);
  FullAdder U320 (w3448, w3347, IN15[7], w3449, w3450);
  FullAdder U321 (w3450, w3349, IN16[7], w3451, w3452);
  FullAdder U322 (w3452, w3351, IN17[7], w3453, w3454);
  FullAdder U323 (w3454, w3353, IN18[7], w3455, w3456);
  FullAdder U324 (w3456, w3355, IN19[7], w3457, w3458);
  FullAdder U325 (w3458, w3357, IN20[7], w3459, w3460);
  FullAdder U326 (w3460, w3359, IN21[7], w3461, w3462);
  FullAdder U327 (w3462, w3361, IN22[7], w3463, w3464);
  FullAdder U328 (w3464, w3363, IN23[7], w3465, w3466);
  FullAdder U329 (w3466, w3365, IN24[7], w3467, w3468);
  FullAdder U330 (w3468, w3367, IN25[7], w3469, w3470);
  FullAdder U331 (w3470, w3369, IN26[7], w3471, w3472);
  FullAdder U332 (w3472, w3371, IN27[7], w3473, w3474);
  FullAdder U333 (w3474, w3373, IN28[7], w3475, w3476);
  FullAdder U334 (w3476, w3375, IN29[7], w3477, w3478);
  FullAdder U335 (w3478, w3377, IN30[7], w3479, w3480);
  FullAdder U336 (w3480, w3379, IN31[7], w3481, w3482);
  FullAdder U337 (w3482, w3381, IN32[7], w3483, w3484);
  FullAdder U338 (w3484, w3383, IN33[7], w3485, w3486);
  FullAdder U339 (w3486, w3385, IN34[7], w3487, w3488);
  FullAdder U340 (w3488, w3387, IN35[7], w3489, w3490);
  FullAdder U341 (w3490, w3389, IN36[7], w3491, w3492);
  FullAdder U342 (w3492, w3391, IN37[7], w3493, w3494);
  FullAdder U343 (w3494, w3393, IN38[7], w3495, w3496);
  FullAdder U344 (w3496, w3395, IN39[7], w3497, w3498);
  FullAdder U345 (w3498, w3397, IN40[7], w3499, w3500);
  FullAdder U346 (w3500, w3399, IN41[7], w3501, w3502);
  FullAdder U347 (w3502, w3401, IN42[7], w3503, w3504);
  FullAdder U348 (w3504, w3403, IN43[7], w3505, w3506);
  FullAdder U349 (w3506, w3405, IN44[7], w3507, w3508);
  FullAdder U350 (w3508, w3407, IN45[7], w3509, w3510);
  FullAdder U351 (w3510, w3409, IN46[7], w3511, w3512);
  FullAdder U352 (w3512, w3411, IN47[7], w3513, w3514);
  FullAdder U353 (w3514, w3413, IN48[7], w3515, w3516);
  FullAdder U354 (w3516, w3415, IN49[7], w3517, w3518);
  FullAdder U355 (w3518, w3417, IN50[7], w3519, w3520);
  FullAdder U356 (w3520, w3419, IN51[7], w3521, w3522);
  FullAdder U357 (w3522, w3421, IN52[7], w3523, w3524);
  FullAdder U358 (w3524, w3423, IN53[5], w3525, w3526);
  FullAdder U359 (w3526, w3425, IN54[4], w3527, w3528);
  FullAdder U360 (w3528, w3427, IN55[3], w3529, w3530);
  FullAdder U361 (w3530, w3429, IN56[2], w3531, w3532);
  FullAdder U362 (w3532, w3431, IN57[1], w3533, w3534);
  FullAdder U363 (w3534, w3432, IN58[0], w3535, w3536);
  HalfAdder U364 (w3435, IN8[8], Out1[8], w3538);
  FullAdder U365 (w3538, w3437, IN9[8], w3539, w3540);
  FullAdder U366 (w3540, w3439, IN10[8], w3541, w3542);
  FullAdder U367 (w3542, w3441, IN11[8], w3543, w3544);
  FullAdder U368 (w3544, w3443, IN12[8], w3545, w3546);
  FullAdder U369 (w3546, w3445, IN13[8], w3547, w3548);
  FullAdder U370 (w3548, w3447, IN14[8], w3549, w3550);
  FullAdder U371 (w3550, w3449, IN15[8], w3551, w3552);
  FullAdder U372 (w3552, w3451, IN16[8], w3553, w3554);
  FullAdder U373 (w3554, w3453, IN17[8], w3555, w3556);
  FullAdder U374 (w3556, w3455, IN18[8], w3557, w3558);
  FullAdder U375 (w3558, w3457, IN19[8], w3559, w3560);
  FullAdder U376 (w3560, w3459, IN20[8], w3561, w3562);
  FullAdder U377 (w3562, w3461, IN21[8], w3563, w3564);
  FullAdder U378 (w3564, w3463, IN22[8], w3565, w3566);
  FullAdder U379 (w3566, w3465, IN23[8], w3567, w3568);
  FullAdder U380 (w3568, w3467, IN24[8], w3569, w3570);
  FullAdder U381 (w3570, w3469, IN25[8], w3571, w3572);
  FullAdder U382 (w3572, w3471, IN26[8], w3573, w3574);
  FullAdder U383 (w3574, w3473, IN27[8], w3575, w3576);
  FullAdder U384 (w3576, w3475, IN28[8], w3577, w3578);
  FullAdder U385 (w3578, w3477, IN29[8], w3579, w3580);
  FullAdder U386 (w3580, w3479, IN30[8], w3581, w3582);
  FullAdder U387 (w3582, w3481, IN31[8], w3583, w3584);
  FullAdder U388 (w3584, w3483, IN32[8], w3585, w3586);
  FullAdder U389 (w3586, w3485, IN33[8], w3587, w3588);
  FullAdder U390 (w3588, w3487, IN34[8], w3589, w3590);
  FullAdder U391 (w3590, w3489, IN35[8], w3591, w3592);
  FullAdder U392 (w3592, w3491, IN36[8], w3593, w3594);
  FullAdder U393 (w3594, w3493, IN37[8], w3595, w3596);
  FullAdder U394 (w3596, w3495, IN38[8], w3597, w3598);
  FullAdder U395 (w3598, w3497, IN39[8], w3599, w3600);
  FullAdder U396 (w3600, w3499, IN40[8], w3601, w3602);
  FullAdder U397 (w3602, w3501, IN41[8], w3603, w3604);
  FullAdder U398 (w3604, w3503, IN42[8], w3605, w3606);
  FullAdder U399 (w3606, w3505, IN43[8], w3607, w3608);
  FullAdder U400 (w3608, w3507, IN44[8], w3609, w3610);
  FullAdder U401 (w3610, w3509, IN45[8], w3611, w3612);
  FullAdder U402 (w3612, w3511, IN46[8], w3613, w3614);
  FullAdder U403 (w3614, w3513, IN47[8], w3615, w3616);
  FullAdder U404 (w3616, w3515, IN48[8], w3617, w3618);
  FullAdder U405 (w3618, w3517, IN49[8], w3619, w3620);
  FullAdder U406 (w3620, w3519, IN50[8], w3621, w3622);
  FullAdder U407 (w3622, w3521, IN51[8], w3623, w3624);
  FullAdder U408 (w3624, w3523, IN52[8], w3625, w3626);
  FullAdder U409 (w3626, w3525, IN53[6], w3627, w3628);
  FullAdder U410 (w3628, w3527, IN54[5], w3629, w3630);
  FullAdder U411 (w3630, w3529, IN55[4], w3631, w3632);
  FullAdder U412 (w3632, w3531, IN56[3], w3633, w3634);
  FullAdder U413 (w3634, w3533, IN57[2], w3635, w3636);
  FullAdder U414 (w3636, w3535, IN58[1], w3637, w3638);
  FullAdder U415 (w3638, w3536, IN59[0], w3639, w3640);
  HalfAdder U416 (w3539, IN9[9], Out1[9], w3642);
  FullAdder U417 (w3642, w3541, IN10[9], w3643, w3644);
  FullAdder U418 (w3644, w3543, IN11[9], w3645, w3646);
  FullAdder U419 (w3646, w3545, IN12[9], w3647, w3648);
  FullAdder U420 (w3648, w3547, IN13[9], w3649, w3650);
  FullAdder U421 (w3650, w3549, IN14[9], w3651, w3652);
  FullAdder U422 (w3652, w3551, IN15[9], w3653, w3654);
  FullAdder U423 (w3654, w3553, IN16[9], w3655, w3656);
  FullAdder U424 (w3656, w3555, IN17[9], w3657, w3658);
  FullAdder U425 (w3658, w3557, IN18[9], w3659, w3660);
  FullAdder U426 (w3660, w3559, IN19[9], w3661, w3662);
  FullAdder U427 (w3662, w3561, IN20[9], w3663, w3664);
  FullAdder U428 (w3664, w3563, IN21[9], w3665, w3666);
  FullAdder U429 (w3666, w3565, IN22[9], w3667, w3668);
  FullAdder U430 (w3668, w3567, IN23[9], w3669, w3670);
  FullAdder U431 (w3670, w3569, IN24[9], w3671, w3672);
  FullAdder U432 (w3672, w3571, IN25[9], w3673, w3674);
  FullAdder U433 (w3674, w3573, IN26[9], w3675, w3676);
  FullAdder U434 (w3676, w3575, IN27[9], w3677, w3678);
  FullAdder U435 (w3678, w3577, IN28[9], w3679, w3680);
  FullAdder U436 (w3680, w3579, IN29[9], w3681, w3682);
  FullAdder U437 (w3682, w3581, IN30[9], w3683, w3684);
  FullAdder U438 (w3684, w3583, IN31[9], w3685, w3686);
  FullAdder U439 (w3686, w3585, IN32[9], w3687, w3688);
  FullAdder U440 (w3688, w3587, IN33[9], w3689, w3690);
  FullAdder U441 (w3690, w3589, IN34[9], w3691, w3692);
  FullAdder U442 (w3692, w3591, IN35[9], w3693, w3694);
  FullAdder U443 (w3694, w3593, IN36[9], w3695, w3696);
  FullAdder U444 (w3696, w3595, IN37[9], w3697, w3698);
  FullAdder U445 (w3698, w3597, IN38[9], w3699, w3700);
  FullAdder U446 (w3700, w3599, IN39[9], w3701, w3702);
  FullAdder U447 (w3702, w3601, IN40[9], w3703, w3704);
  FullAdder U448 (w3704, w3603, IN41[9], w3705, w3706);
  FullAdder U449 (w3706, w3605, IN42[9], w3707, w3708);
  FullAdder U450 (w3708, w3607, IN43[9], w3709, w3710);
  FullAdder U451 (w3710, w3609, IN44[9], w3711, w3712);
  FullAdder U452 (w3712, w3611, IN45[9], w3713, w3714);
  FullAdder U453 (w3714, w3613, IN46[9], w3715, w3716);
  FullAdder U454 (w3716, w3615, IN47[9], w3717, w3718);
  FullAdder U455 (w3718, w3617, IN48[9], w3719, w3720);
  FullAdder U456 (w3720, w3619, IN49[9], w3721, w3722);
  FullAdder U457 (w3722, w3621, IN50[9], w3723, w3724);
  FullAdder U458 (w3724, w3623, IN51[9], w3725, w3726);
  FullAdder U459 (w3726, w3625, IN52[9], w3727, w3728);
  FullAdder U460 (w3728, w3627, IN53[7], w3729, w3730);
  FullAdder U461 (w3730, w3629, IN54[6], w3731, w3732);
  FullAdder U462 (w3732, w3631, IN55[5], w3733, w3734);
  FullAdder U463 (w3734, w3633, IN56[4], w3735, w3736);
  FullAdder U464 (w3736, w3635, IN57[3], w3737, w3738);
  FullAdder U465 (w3738, w3637, IN58[2], w3739, w3740);
  FullAdder U466 (w3740, w3639, IN59[1], w3741, w3742);
  FullAdder U467 (w3742, w3640, IN60[0], w3743, w3744);
  HalfAdder U468 (w3643, IN10[10], Out1[10], w3746);
  FullAdder U469 (w3746, w3645, IN11[10], w3747, w3748);
  FullAdder U470 (w3748, w3647, IN12[10], w3749, w3750);
  FullAdder U471 (w3750, w3649, IN13[10], w3751, w3752);
  FullAdder U472 (w3752, w3651, IN14[10], w3753, w3754);
  FullAdder U473 (w3754, w3653, IN15[10], w3755, w3756);
  FullAdder U474 (w3756, w3655, IN16[10], w3757, w3758);
  FullAdder U475 (w3758, w3657, IN17[10], w3759, w3760);
  FullAdder U476 (w3760, w3659, IN18[10], w3761, w3762);
  FullAdder U477 (w3762, w3661, IN19[10], w3763, w3764);
  FullAdder U478 (w3764, w3663, IN20[10], w3765, w3766);
  FullAdder U479 (w3766, w3665, IN21[10], w3767, w3768);
  FullAdder U480 (w3768, w3667, IN22[10], w3769, w3770);
  FullAdder U481 (w3770, w3669, IN23[10], w3771, w3772);
  FullAdder U482 (w3772, w3671, IN24[10], w3773, w3774);
  FullAdder U483 (w3774, w3673, IN25[10], w3775, w3776);
  FullAdder U484 (w3776, w3675, IN26[10], w3777, w3778);
  FullAdder U485 (w3778, w3677, IN27[10], w3779, w3780);
  FullAdder U486 (w3780, w3679, IN28[10], w3781, w3782);
  FullAdder U487 (w3782, w3681, IN29[10], w3783, w3784);
  FullAdder U488 (w3784, w3683, IN30[10], w3785, w3786);
  FullAdder U489 (w3786, w3685, IN31[10], w3787, w3788);
  FullAdder U490 (w3788, w3687, IN32[10], w3789, w3790);
  FullAdder U491 (w3790, w3689, IN33[10], w3791, w3792);
  FullAdder U492 (w3792, w3691, IN34[10], w3793, w3794);
  FullAdder U493 (w3794, w3693, IN35[10], w3795, w3796);
  FullAdder U494 (w3796, w3695, IN36[10], w3797, w3798);
  FullAdder U495 (w3798, w3697, IN37[10], w3799, w3800);
  FullAdder U496 (w3800, w3699, IN38[10], w3801, w3802);
  FullAdder U497 (w3802, w3701, IN39[10], w3803, w3804);
  FullAdder U498 (w3804, w3703, IN40[10], w3805, w3806);
  FullAdder U499 (w3806, w3705, IN41[10], w3807, w3808);
  FullAdder U500 (w3808, w3707, IN42[10], w3809, w3810);
  FullAdder U501 (w3810, w3709, IN43[10], w3811, w3812);
  FullAdder U502 (w3812, w3711, IN44[10], w3813, w3814);
  FullAdder U503 (w3814, w3713, IN45[10], w3815, w3816);
  FullAdder U504 (w3816, w3715, IN46[10], w3817, w3818);
  FullAdder U505 (w3818, w3717, IN47[10], w3819, w3820);
  FullAdder U506 (w3820, w3719, IN48[10], w3821, w3822);
  FullAdder U507 (w3822, w3721, IN49[10], w3823, w3824);
  FullAdder U508 (w3824, w3723, IN50[10], w3825, w3826);
  FullAdder U509 (w3826, w3725, IN51[10], w3827, w3828);
  FullAdder U510 (w3828, w3727, IN52[10], w3829, w3830);
  FullAdder U511 (w3830, w3729, IN53[8], w3831, w3832);
  FullAdder U512 (w3832, w3731, IN54[7], w3833, w3834);
  FullAdder U513 (w3834, w3733, IN55[6], w3835, w3836);
  FullAdder U514 (w3836, w3735, IN56[5], w3837, w3838);
  FullAdder U515 (w3838, w3737, IN57[4], w3839, w3840);
  FullAdder U516 (w3840, w3739, IN58[3], w3841, w3842);
  FullAdder U517 (w3842, w3741, IN59[2], w3843, w3844);
  FullAdder U518 (w3844, w3743, IN60[1], w3845, w3846);
  FullAdder U519 (w3846, w3744, IN61[0], w3847, w3848);
  HalfAdder U520 (w3747, IN11[11], Out1[11], w3850);
  FullAdder U521 (w3850, w3749, IN12[11], w3851, w3852);
  FullAdder U522 (w3852, w3751, IN13[11], w3853, w3854);
  FullAdder U523 (w3854, w3753, IN14[11], w3855, w3856);
  FullAdder U524 (w3856, w3755, IN15[11], w3857, w3858);
  FullAdder U525 (w3858, w3757, IN16[11], w3859, w3860);
  FullAdder U526 (w3860, w3759, IN17[11], w3861, w3862);
  FullAdder U527 (w3862, w3761, IN18[11], w3863, w3864);
  FullAdder U528 (w3864, w3763, IN19[11], w3865, w3866);
  FullAdder U529 (w3866, w3765, IN20[11], w3867, w3868);
  FullAdder U530 (w3868, w3767, IN21[11], w3869, w3870);
  FullAdder U531 (w3870, w3769, IN22[11], w3871, w3872);
  FullAdder U532 (w3872, w3771, IN23[11], w3873, w3874);
  FullAdder U533 (w3874, w3773, IN24[11], w3875, w3876);
  FullAdder U534 (w3876, w3775, IN25[11], w3877, w3878);
  FullAdder U535 (w3878, w3777, IN26[11], w3879, w3880);
  FullAdder U536 (w3880, w3779, IN27[11], w3881, w3882);
  FullAdder U537 (w3882, w3781, IN28[11], w3883, w3884);
  FullAdder U538 (w3884, w3783, IN29[11], w3885, w3886);
  FullAdder U539 (w3886, w3785, IN30[11], w3887, w3888);
  FullAdder U540 (w3888, w3787, IN31[11], w3889, w3890);
  FullAdder U541 (w3890, w3789, IN32[11], w3891, w3892);
  FullAdder U542 (w3892, w3791, IN33[11], w3893, w3894);
  FullAdder U543 (w3894, w3793, IN34[11], w3895, w3896);
  FullAdder U544 (w3896, w3795, IN35[11], w3897, w3898);
  FullAdder U545 (w3898, w3797, IN36[11], w3899, w3900);
  FullAdder U546 (w3900, w3799, IN37[11], w3901, w3902);
  FullAdder U547 (w3902, w3801, IN38[11], w3903, w3904);
  FullAdder U548 (w3904, w3803, IN39[11], w3905, w3906);
  FullAdder U549 (w3906, w3805, IN40[11], w3907, w3908);
  FullAdder U550 (w3908, w3807, IN41[11], w3909, w3910);
  FullAdder U551 (w3910, w3809, IN42[11], w3911, w3912);
  FullAdder U552 (w3912, w3811, IN43[11], w3913, w3914);
  FullAdder U553 (w3914, w3813, IN44[11], w3915, w3916);
  FullAdder U554 (w3916, w3815, IN45[11], w3917, w3918);
  FullAdder U555 (w3918, w3817, IN46[11], w3919, w3920);
  FullAdder U556 (w3920, w3819, IN47[11], w3921, w3922);
  FullAdder U557 (w3922, w3821, IN48[11], w3923, w3924);
  FullAdder U558 (w3924, w3823, IN49[11], w3925, w3926);
  FullAdder U559 (w3926, w3825, IN50[11], w3927, w3928);
  FullAdder U560 (w3928, w3827, IN51[11], w3929, w3930);
  FullAdder U561 (w3930, w3829, IN52[11], w3931, w3932);
  FullAdder U562 (w3932, w3831, IN53[9], w3933, w3934);
  FullAdder U563 (w3934, w3833, IN54[8], w3935, w3936);
  FullAdder U564 (w3936, w3835, IN55[7], w3937, w3938);
  FullAdder U565 (w3938, w3837, IN56[6], w3939, w3940);
  FullAdder U566 (w3940, w3839, IN57[5], w3941, w3942);
  FullAdder U567 (w3942, w3841, IN58[4], w3943, w3944);
  FullAdder U568 (w3944, w3843, IN59[3], w3945, w3946);
  FullAdder U569 (w3946, w3845, IN60[2], w3947, w3948);
  FullAdder U570 (w3948, w3847, IN61[1], w3949, w3950);
  FullAdder U571 (w3950, w3848, IN62[0], w3951, w3952);
  HalfAdder U572 (w3851, IN12[12], Out1[12], w3954);
  FullAdder U573 (w3954, w3853, IN13[12], w3955, w3956);
  FullAdder U574 (w3956, w3855, IN14[12], w3957, w3958);
  FullAdder U575 (w3958, w3857, IN15[12], w3959, w3960);
  FullAdder U576 (w3960, w3859, IN16[12], w3961, w3962);
  FullAdder U577 (w3962, w3861, IN17[12], w3963, w3964);
  FullAdder U578 (w3964, w3863, IN18[12], w3965, w3966);
  FullAdder U579 (w3966, w3865, IN19[12], w3967, w3968);
  FullAdder U580 (w3968, w3867, IN20[12], w3969, w3970);
  FullAdder U581 (w3970, w3869, IN21[12], w3971, w3972);
  FullAdder U582 (w3972, w3871, IN22[12], w3973, w3974);
  FullAdder U583 (w3974, w3873, IN23[12], w3975, w3976);
  FullAdder U584 (w3976, w3875, IN24[12], w3977, w3978);
  FullAdder U585 (w3978, w3877, IN25[12], w3979, w3980);
  FullAdder U586 (w3980, w3879, IN26[12], w3981, w3982);
  FullAdder U587 (w3982, w3881, IN27[12], w3983, w3984);
  FullAdder U588 (w3984, w3883, IN28[12], w3985, w3986);
  FullAdder U589 (w3986, w3885, IN29[12], w3987, w3988);
  FullAdder U590 (w3988, w3887, IN30[12], w3989, w3990);
  FullAdder U591 (w3990, w3889, IN31[12], w3991, w3992);
  FullAdder U592 (w3992, w3891, IN32[12], w3993, w3994);
  FullAdder U593 (w3994, w3893, IN33[12], w3995, w3996);
  FullAdder U594 (w3996, w3895, IN34[12], w3997, w3998);
  FullAdder U595 (w3998, w3897, IN35[12], w3999, w4000);
  FullAdder U596 (w4000, w3899, IN36[12], w4001, w4002);
  FullAdder U597 (w4002, w3901, IN37[12], w4003, w4004);
  FullAdder U598 (w4004, w3903, IN38[12], w4005, w4006);
  FullAdder U599 (w4006, w3905, IN39[12], w4007, w4008);
  FullAdder U600 (w4008, w3907, IN40[12], w4009, w4010);
  FullAdder U601 (w4010, w3909, IN41[12], w4011, w4012);
  FullAdder U602 (w4012, w3911, IN42[12], w4013, w4014);
  FullAdder U603 (w4014, w3913, IN43[12], w4015, w4016);
  FullAdder U604 (w4016, w3915, IN44[12], w4017, w4018);
  FullAdder U605 (w4018, w3917, IN45[12], w4019, w4020);
  FullAdder U606 (w4020, w3919, IN46[12], w4021, w4022);
  FullAdder U607 (w4022, w3921, IN47[12], w4023, w4024);
  FullAdder U608 (w4024, w3923, IN48[12], w4025, w4026);
  FullAdder U609 (w4026, w3925, IN49[12], w4027, w4028);
  FullAdder U610 (w4028, w3927, IN50[12], w4029, w4030);
  FullAdder U611 (w4030, w3929, IN51[12], w4031, w4032);
  FullAdder U612 (w4032, w3931, IN52[12], w4033, w4034);
  FullAdder U613 (w4034, w3933, IN53[10], w4035, w4036);
  FullAdder U614 (w4036, w3935, IN54[9], w4037, w4038);
  FullAdder U615 (w4038, w3937, IN55[8], w4039, w4040);
  FullAdder U616 (w4040, w3939, IN56[7], w4041, w4042);
  FullAdder U617 (w4042, w3941, IN57[6], w4043, w4044);
  FullAdder U618 (w4044, w3943, IN58[5], w4045, w4046);
  FullAdder U619 (w4046, w3945, IN59[4], w4047, w4048);
  FullAdder U620 (w4048, w3947, IN60[3], w4049, w4050);
  FullAdder U621 (w4050, w3949, IN61[2], w4051, w4052);
  FullAdder U622 (w4052, w3951, IN62[1], w4053, w4054);
  FullAdder U623 (w4054, w3952, IN63[0], w4055, w4056);
  HalfAdder U624 (w3955, IN13[13], Out1[13], w4058);
  FullAdder U625 (w4058, w3957, IN14[13], w4059, w4060);
  FullAdder U626 (w4060, w3959, IN15[13], w4061, w4062);
  FullAdder U627 (w4062, w3961, IN16[13], w4063, w4064);
  FullAdder U628 (w4064, w3963, IN17[13], w4065, w4066);
  FullAdder U629 (w4066, w3965, IN18[13], w4067, w4068);
  FullAdder U630 (w4068, w3967, IN19[13], w4069, w4070);
  FullAdder U631 (w4070, w3969, IN20[13], w4071, w4072);
  FullAdder U632 (w4072, w3971, IN21[13], w4073, w4074);
  FullAdder U633 (w4074, w3973, IN22[13], w4075, w4076);
  FullAdder U634 (w4076, w3975, IN23[13], w4077, w4078);
  FullAdder U635 (w4078, w3977, IN24[13], w4079, w4080);
  FullAdder U636 (w4080, w3979, IN25[13], w4081, w4082);
  FullAdder U637 (w4082, w3981, IN26[13], w4083, w4084);
  FullAdder U638 (w4084, w3983, IN27[13], w4085, w4086);
  FullAdder U639 (w4086, w3985, IN28[13], w4087, w4088);
  FullAdder U640 (w4088, w3987, IN29[13], w4089, w4090);
  FullAdder U641 (w4090, w3989, IN30[13], w4091, w4092);
  FullAdder U642 (w4092, w3991, IN31[13], w4093, w4094);
  FullAdder U643 (w4094, w3993, IN32[13], w4095, w4096);
  FullAdder U644 (w4096, w3995, IN33[13], w4097, w4098);
  FullAdder U645 (w4098, w3997, IN34[13], w4099, w4100);
  FullAdder U646 (w4100, w3999, IN35[13], w4101, w4102);
  FullAdder U647 (w4102, w4001, IN36[13], w4103, w4104);
  FullAdder U648 (w4104, w4003, IN37[13], w4105, w4106);
  FullAdder U649 (w4106, w4005, IN38[13], w4107, w4108);
  FullAdder U650 (w4108, w4007, IN39[13], w4109, w4110);
  FullAdder U651 (w4110, w4009, IN40[13], w4111, w4112);
  FullAdder U652 (w4112, w4011, IN41[13], w4113, w4114);
  FullAdder U653 (w4114, w4013, IN42[13], w4115, w4116);
  FullAdder U654 (w4116, w4015, IN43[13], w4117, w4118);
  FullAdder U655 (w4118, w4017, IN44[13], w4119, w4120);
  FullAdder U656 (w4120, w4019, IN45[13], w4121, w4122);
  FullAdder U657 (w4122, w4021, IN46[13], w4123, w4124);
  FullAdder U658 (w4124, w4023, IN47[13], w4125, w4126);
  FullAdder U659 (w4126, w4025, IN48[13], w4127, w4128);
  FullAdder U660 (w4128, w4027, IN49[13], w4129, w4130);
  FullAdder U661 (w4130, w4029, IN50[13], w4131, w4132);
  FullAdder U662 (w4132, w4031, IN51[13], w4133, w4134);
  FullAdder U663 (w4134, w4033, IN52[13], w4135, w4136);
  FullAdder U664 (w4136, w4035, IN53[11], w4137, w4138);
  FullAdder U665 (w4138, w4037, IN54[10], w4139, w4140);
  FullAdder U666 (w4140, w4039, IN55[9], w4141, w4142);
  FullAdder U667 (w4142, w4041, IN56[8], w4143, w4144);
  FullAdder U668 (w4144, w4043, IN57[7], w4145, w4146);
  FullAdder U669 (w4146, w4045, IN58[6], w4147, w4148);
  FullAdder U670 (w4148, w4047, IN59[5], w4149, w4150);
  FullAdder U671 (w4150, w4049, IN60[4], w4151, w4152);
  FullAdder U672 (w4152, w4051, IN61[3], w4153, w4154);
  FullAdder U673 (w4154, w4053, IN62[2], w4155, w4156);
  FullAdder U674 (w4156, w4055, IN63[1], w4157, w4158);
  FullAdder U675 (w4158, w4056, IN64[0], w4159, w4160);
  HalfAdder U676 (w4059, IN14[14], Out1[14], w4162);
  FullAdder U677 (w4162, w4061, IN15[14], w4163, w4164);
  FullAdder U678 (w4164, w4063, IN16[14], w4165, w4166);
  FullAdder U679 (w4166, w4065, IN17[14], w4167, w4168);
  FullAdder U680 (w4168, w4067, IN18[14], w4169, w4170);
  FullAdder U681 (w4170, w4069, IN19[14], w4171, w4172);
  FullAdder U682 (w4172, w4071, IN20[14], w4173, w4174);
  FullAdder U683 (w4174, w4073, IN21[14], w4175, w4176);
  FullAdder U684 (w4176, w4075, IN22[14], w4177, w4178);
  FullAdder U685 (w4178, w4077, IN23[14], w4179, w4180);
  FullAdder U686 (w4180, w4079, IN24[14], w4181, w4182);
  FullAdder U687 (w4182, w4081, IN25[14], w4183, w4184);
  FullAdder U688 (w4184, w4083, IN26[14], w4185, w4186);
  FullAdder U689 (w4186, w4085, IN27[14], w4187, w4188);
  FullAdder U690 (w4188, w4087, IN28[14], w4189, w4190);
  FullAdder U691 (w4190, w4089, IN29[14], w4191, w4192);
  FullAdder U692 (w4192, w4091, IN30[14], w4193, w4194);
  FullAdder U693 (w4194, w4093, IN31[14], w4195, w4196);
  FullAdder U694 (w4196, w4095, IN32[14], w4197, w4198);
  FullAdder U695 (w4198, w4097, IN33[14], w4199, w4200);
  FullAdder U696 (w4200, w4099, IN34[14], w4201, w4202);
  FullAdder U697 (w4202, w4101, IN35[14], w4203, w4204);
  FullAdder U698 (w4204, w4103, IN36[14], w4205, w4206);
  FullAdder U699 (w4206, w4105, IN37[14], w4207, w4208);
  FullAdder U700 (w4208, w4107, IN38[14], w4209, w4210);
  FullAdder U701 (w4210, w4109, IN39[14], w4211, w4212);
  FullAdder U702 (w4212, w4111, IN40[14], w4213, w4214);
  FullAdder U703 (w4214, w4113, IN41[14], w4215, w4216);
  FullAdder U704 (w4216, w4115, IN42[14], w4217, w4218);
  FullAdder U705 (w4218, w4117, IN43[14], w4219, w4220);
  FullAdder U706 (w4220, w4119, IN44[14], w4221, w4222);
  FullAdder U707 (w4222, w4121, IN45[14], w4223, w4224);
  FullAdder U708 (w4224, w4123, IN46[14], w4225, w4226);
  FullAdder U709 (w4226, w4125, IN47[14], w4227, w4228);
  FullAdder U710 (w4228, w4127, IN48[14], w4229, w4230);
  FullAdder U711 (w4230, w4129, IN49[14], w4231, w4232);
  FullAdder U712 (w4232, w4131, IN50[14], w4233, w4234);
  FullAdder U713 (w4234, w4133, IN51[14], w4235, w4236);
  FullAdder U714 (w4236, w4135, IN52[14], w4237, w4238);
  FullAdder U715 (w4238, w4137, IN53[12], w4239, w4240);
  FullAdder U716 (w4240, w4139, IN54[11], w4241, w4242);
  FullAdder U717 (w4242, w4141, IN55[10], w4243, w4244);
  FullAdder U718 (w4244, w4143, IN56[9], w4245, w4246);
  FullAdder U719 (w4246, w4145, IN57[8], w4247, w4248);
  FullAdder U720 (w4248, w4147, IN58[7], w4249, w4250);
  FullAdder U721 (w4250, w4149, IN59[6], w4251, w4252);
  FullAdder U722 (w4252, w4151, IN60[5], w4253, w4254);
  FullAdder U723 (w4254, w4153, IN61[4], w4255, w4256);
  FullAdder U724 (w4256, w4155, IN62[3], w4257, w4258);
  FullAdder U725 (w4258, w4157, IN63[2], w4259, w4260);
  FullAdder U726 (w4260, w4159, IN64[1], w4261, w4262);
  FullAdder U727 (w4262, w4160, IN65[0], w4263, w4264);
  HalfAdder U728 (w4163, IN15[15], Out1[15], w4266);
  FullAdder U729 (w4266, w4165, IN16[15], w4267, w4268);
  FullAdder U730 (w4268, w4167, IN17[15], w4269, w4270);
  FullAdder U731 (w4270, w4169, IN18[15], w4271, w4272);
  FullAdder U732 (w4272, w4171, IN19[15], w4273, w4274);
  FullAdder U733 (w4274, w4173, IN20[15], w4275, w4276);
  FullAdder U734 (w4276, w4175, IN21[15], w4277, w4278);
  FullAdder U735 (w4278, w4177, IN22[15], w4279, w4280);
  FullAdder U736 (w4280, w4179, IN23[15], w4281, w4282);
  FullAdder U737 (w4282, w4181, IN24[15], w4283, w4284);
  FullAdder U738 (w4284, w4183, IN25[15], w4285, w4286);
  FullAdder U739 (w4286, w4185, IN26[15], w4287, w4288);
  FullAdder U740 (w4288, w4187, IN27[15], w4289, w4290);
  FullAdder U741 (w4290, w4189, IN28[15], w4291, w4292);
  FullAdder U742 (w4292, w4191, IN29[15], w4293, w4294);
  FullAdder U743 (w4294, w4193, IN30[15], w4295, w4296);
  FullAdder U744 (w4296, w4195, IN31[15], w4297, w4298);
  FullAdder U745 (w4298, w4197, IN32[15], w4299, w4300);
  FullAdder U746 (w4300, w4199, IN33[15], w4301, w4302);
  FullAdder U747 (w4302, w4201, IN34[15], w4303, w4304);
  FullAdder U748 (w4304, w4203, IN35[15], w4305, w4306);
  FullAdder U749 (w4306, w4205, IN36[15], w4307, w4308);
  FullAdder U750 (w4308, w4207, IN37[15], w4309, w4310);
  FullAdder U751 (w4310, w4209, IN38[15], w4311, w4312);
  FullAdder U752 (w4312, w4211, IN39[15], w4313, w4314);
  FullAdder U753 (w4314, w4213, IN40[15], w4315, w4316);
  FullAdder U754 (w4316, w4215, IN41[15], w4317, w4318);
  FullAdder U755 (w4318, w4217, IN42[15], w4319, w4320);
  FullAdder U756 (w4320, w4219, IN43[15], w4321, w4322);
  FullAdder U757 (w4322, w4221, IN44[15], w4323, w4324);
  FullAdder U758 (w4324, w4223, IN45[15], w4325, w4326);
  FullAdder U759 (w4326, w4225, IN46[15], w4327, w4328);
  FullAdder U760 (w4328, w4227, IN47[15], w4329, w4330);
  FullAdder U761 (w4330, w4229, IN48[15], w4331, w4332);
  FullAdder U762 (w4332, w4231, IN49[15], w4333, w4334);
  FullAdder U763 (w4334, w4233, IN50[15], w4335, w4336);
  FullAdder U764 (w4336, w4235, IN51[15], w4337, w4338);
  FullAdder U765 (w4338, w4237, IN52[15], w4339, w4340);
  FullAdder U766 (w4340, w4239, IN53[13], w4341, w4342);
  FullAdder U767 (w4342, w4241, IN54[12], w4343, w4344);
  FullAdder U768 (w4344, w4243, IN55[11], w4345, w4346);
  FullAdder U769 (w4346, w4245, IN56[10], w4347, w4348);
  FullAdder U770 (w4348, w4247, IN57[9], w4349, w4350);
  FullAdder U771 (w4350, w4249, IN58[8], w4351, w4352);
  FullAdder U772 (w4352, w4251, IN59[7], w4353, w4354);
  FullAdder U773 (w4354, w4253, IN60[6], w4355, w4356);
  FullAdder U774 (w4356, w4255, IN61[5], w4357, w4358);
  FullAdder U775 (w4358, w4257, IN62[4], w4359, w4360);
  FullAdder U776 (w4360, w4259, IN63[3], w4361, w4362);
  FullAdder U777 (w4362, w4261, IN64[2], w4363, w4364);
  FullAdder U778 (w4364, w4263, IN65[1], w4365, w4366);
  FullAdder U779 (w4366, w4264, IN66[0], w4367, w4368);
  HalfAdder U780 (w4267, IN16[16], Out1[16], w4370);
  FullAdder U781 (w4370, w4269, IN17[16], w4371, w4372);
  FullAdder U782 (w4372, w4271, IN18[16], w4373, w4374);
  FullAdder U783 (w4374, w4273, IN19[16], w4375, w4376);
  FullAdder U784 (w4376, w4275, IN20[16], w4377, w4378);
  FullAdder U785 (w4378, w4277, IN21[16], w4379, w4380);
  FullAdder U786 (w4380, w4279, IN22[16], w4381, w4382);
  FullAdder U787 (w4382, w4281, IN23[16], w4383, w4384);
  FullAdder U788 (w4384, w4283, IN24[16], w4385, w4386);
  FullAdder U789 (w4386, w4285, IN25[16], w4387, w4388);
  FullAdder U790 (w4388, w4287, IN26[16], w4389, w4390);
  FullAdder U791 (w4390, w4289, IN27[16], w4391, w4392);
  FullAdder U792 (w4392, w4291, IN28[16], w4393, w4394);
  FullAdder U793 (w4394, w4293, IN29[16], w4395, w4396);
  FullAdder U794 (w4396, w4295, IN30[16], w4397, w4398);
  FullAdder U795 (w4398, w4297, IN31[16], w4399, w4400);
  FullAdder U796 (w4400, w4299, IN32[16], w4401, w4402);
  FullAdder U797 (w4402, w4301, IN33[16], w4403, w4404);
  FullAdder U798 (w4404, w4303, IN34[16], w4405, w4406);
  FullAdder U799 (w4406, w4305, IN35[16], w4407, w4408);
  FullAdder U800 (w4408, w4307, IN36[16], w4409, w4410);
  FullAdder U801 (w4410, w4309, IN37[16], w4411, w4412);
  FullAdder U802 (w4412, w4311, IN38[16], w4413, w4414);
  FullAdder U803 (w4414, w4313, IN39[16], w4415, w4416);
  FullAdder U804 (w4416, w4315, IN40[16], w4417, w4418);
  FullAdder U805 (w4418, w4317, IN41[16], w4419, w4420);
  FullAdder U806 (w4420, w4319, IN42[16], w4421, w4422);
  FullAdder U807 (w4422, w4321, IN43[16], w4423, w4424);
  FullAdder U808 (w4424, w4323, IN44[16], w4425, w4426);
  FullAdder U809 (w4426, w4325, IN45[16], w4427, w4428);
  FullAdder U810 (w4428, w4327, IN46[16], w4429, w4430);
  FullAdder U811 (w4430, w4329, IN47[16], w4431, w4432);
  FullAdder U812 (w4432, w4331, IN48[16], w4433, w4434);
  FullAdder U813 (w4434, w4333, IN49[16], w4435, w4436);
  FullAdder U814 (w4436, w4335, IN50[16], w4437, w4438);
  FullAdder U815 (w4438, w4337, IN51[16], w4439, w4440);
  FullAdder U816 (w4440, w4339, IN52[16], w4441, w4442);
  FullAdder U817 (w4442, w4341, IN53[14], w4443, w4444);
  FullAdder U818 (w4444, w4343, IN54[13], w4445, w4446);
  FullAdder U819 (w4446, w4345, IN55[12], w4447, w4448);
  FullAdder U820 (w4448, w4347, IN56[11], w4449, w4450);
  FullAdder U821 (w4450, w4349, IN57[10], w4451, w4452);
  FullAdder U822 (w4452, w4351, IN58[9], w4453, w4454);
  FullAdder U823 (w4454, w4353, IN59[8], w4455, w4456);
  FullAdder U824 (w4456, w4355, IN60[7], w4457, w4458);
  FullAdder U825 (w4458, w4357, IN61[6], w4459, w4460);
  FullAdder U826 (w4460, w4359, IN62[5], w4461, w4462);
  FullAdder U827 (w4462, w4361, IN63[4], w4463, w4464);
  FullAdder U828 (w4464, w4363, IN64[3], w4465, w4466);
  FullAdder U829 (w4466, w4365, IN65[2], w4467, w4468);
  FullAdder U830 (w4468, w4367, IN66[1], w4469, w4470);
  FullAdder U831 (w4470, w4368, IN67[0], w4471, w4472);
  HalfAdder U832 (w4371, IN17[17], Out1[17], w4474);
  FullAdder U833 (w4474, w4373, IN18[17], w4475, w4476);
  FullAdder U834 (w4476, w4375, IN19[17], w4477, w4478);
  FullAdder U835 (w4478, w4377, IN20[17], w4479, w4480);
  FullAdder U836 (w4480, w4379, IN21[17], w4481, w4482);
  FullAdder U837 (w4482, w4381, IN22[17], w4483, w4484);
  FullAdder U838 (w4484, w4383, IN23[17], w4485, w4486);
  FullAdder U839 (w4486, w4385, IN24[17], w4487, w4488);
  FullAdder U840 (w4488, w4387, IN25[17], w4489, w4490);
  FullAdder U841 (w4490, w4389, IN26[17], w4491, w4492);
  FullAdder U842 (w4492, w4391, IN27[17], w4493, w4494);
  FullAdder U843 (w4494, w4393, IN28[17], w4495, w4496);
  FullAdder U844 (w4496, w4395, IN29[17], w4497, w4498);
  FullAdder U845 (w4498, w4397, IN30[17], w4499, w4500);
  FullAdder U846 (w4500, w4399, IN31[17], w4501, w4502);
  FullAdder U847 (w4502, w4401, IN32[17], w4503, w4504);
  FullAdder U848 (w4504, w4403, IN33[17], w4505, w4506);
  FullAdder U849 (w4506, w4405, IN34[17], w4507, w4508);
  FullAdder U850 (w4508, w4407, IN35[17], w4509, w4510);
  FullAdder U851 (w4510, w4409, IN36[17], w4511, w4512);
  FullAdder U852 (w4512, w4411, IN37[17], w4513, w4514);
  FullAdder U853 (w4514, w4413, IN38[17], w4515, w4516);
  FullAdder U854 (w4516, w4415, IN39[17], w4517, w4518);
  FullAdder U855 (w4518, w4417, IN40[17], w4519, w4520);
  FullAdder U856 (w4520, w4419, IN41[17], w4521, w4522);
  FullAdder U857 (w4522, w4421, IN42[17], w4523, w4524);
  FullAdder U858 (w4524, w4423, IN43[17], w4525, w4526);
  FullAdder U859 (w4526, w4425, IN44[17], w4527, w4528);
  FullAdder U860 (w4528, w4427, IN45[17], w4529, w4530);
  FullAdder U861 (w4530, w4429, IN46[17], w4531, w4532);
  FullAdder U862 (w4532, w4431, IN47[17], w4533, w4534);
  FullAdder U863 (w4534, w4433, IN48[17], w4535, w4536);
  FullAdder U864 (w4536, w4435, IN49[17], w4537, w4538);
  FullAdder U865 (w4538, w4437, IN50[17], w4539, w4540);
  FullAdder U866 (w4540, w4439, IN51[17], w4541, w4542);
  FullAdder U867 (w4542, w4441, IN52[17], w4543, w4544);
  FullAdder U868 (w4544, w4443, IN53[15], w4545, w4546);
  FullAdder U869 (w4546, w4445, IN54[14], w4547, w4548);
  FullAdder U870 (w4548, w4447, IN55[13], w4549, w4550);
  FullAdder U871 (w4550, w4449, IN56[12], w4551, w4552);
  FullAdder U872 (w4552, w4451, IN57[11], w4553, w4554);
  FullAdder U873 (w4554, w4453, IN58[10], w4555, w4556);
  FullAdder U874 (w4556, w4455, IN59[9], w4557, w4558);
  FullAdder U875 (w4558, w4457, IN60[8], w4559, w4560);
  FullAdder U876 (w4560, w4459, IN61[7], w4561, w4562);
  FullAdder U877 (w4562, w4461, IN62[6], w4563, w4564);
  FullAdder U878 (w4564, w4463, IN63[5], w4565, w4566);
  FullAdder U879 (w4566, w4465, IN64[4], w4567, w4568);
  FullAdder U880 (w4568, w4467, IN65[3], w4569, w4570);
  FullAdder U881 (w4570, w4469, IN66[2], w4571, w4572);
  FullAdder U882 (w4572, w4471, IN67[1], w4573, w4574);
  FullAdder U883 (w4574, w4472, IN68[0], w4575, w4576);
  HalfAdder U884 (w4475, IN18[18], Out1[18], w4578);
  FullAdder U885 (w4578, w4477, IN19[18], w4579, w4580);
  FullAdder U886 (w4580, w4479, IN20[18], w4581, w4582);
  FullAdder U887 (w4582, w4481, IN21[18], w4583, w4584);
  FullAdder U888 (w4584, w4483, IN22[18], w4585, w4586);
  FullAdder U889 (w4586, w4485, IN23[18], w4587, w4588);
  FullAdder U890 (w4588, w4487, IN24[18], w4589, w4590);
  FullAdder U891 (w4590, w4489, IN25[18], w4591, w4592);
  FullAdder U892 (w4592, w4491, IN26[18], w4593, w4594);
  FullAdder U893 (w4594, w4493, IN27[18], w4595, w4596);
  FullAdder U894 (w4596, w4495, IN28[18], w4597, w4598);
  FullAdder U895 (w4598, w4497, IN29[18], w4599, w4600);
  FullAdder U896 (w4600, w4499, IN30[18], w4601, w4602);
  FullAdder U897 (w4602, w4501, IN31[18], w4603, w4604);
  FullAdder U898 (w4604, w4503, IN32[18], w4605, w4606);
  FullAdder U899 (w4606, w4505, IN33[18], w4607, w4608);
  FullAdder U900 (w4608, w4507, IN34[18], w4609, w4610);
  FullAdder U901 (w4610, w4509, IN35[18], w4611, w4612);
  FullAdder U902 (w4612, w4511, IN36[18], w4613, w4614);
  FullAdder U903 (w4614, w4513, IN37[18], w4615, w4616);
  FullAdder U904 (w4616, w4515, IN38[18], w4617, w4618);
  FullAdder U905 (w4618, w4517, IN39[18], w4619, w4620);
  FullAdder U906 (w4620, w4519, IN40[18], w4621, w4622);
  FullAdder U907 (w4622, w4521, IN41[18], w4623, w4624);
  FullAdder U908 (w4624, w4523, IN42[18], w4625, w4626);
  FullAdder U909 (w4626, w4525, IN43[18], w4627, w4628);
  FullAdder U910 (w4628, w4527, IN44[18], w4629, w4630);
  FullAdder U911 (w4630, w4529, IN45[18], w4631, w4632);
  FullAdder U912 (w4632, w4531, IN46[18], w4633, w4634);
  FullAdder U913 (w4634, w4533, IN47[18], w4635, w4636);
  FullAdder U914 (w4636, w4535, IN48[18], w4637, w4638);
  FullAdder U915 (w4638, w4537, IN49[18], w4639, w4640);
  FullAdder U916 (w4640, w4539, IN50[18], w4641, w4642);
  FullAdder U917 (w4642, w4541, IN51[18], w4643, w4644);
  FullAdder U918 (w4644, w4543, IN52[18], w4645, w4646);
  FullAdder U919 (w4646, w4545, IN53[16], w4647, w4648);
  FullAdder U920 (w4648, w4547, IN54[15], w4649, w4650);
  FullAdder U921 (w4650, w4549, IN55[14], w4651, w4652);
  FullAdder U922 (w4652, w4551, IN56[13], w4653, w4654);
  FullAdder U923 (w4654, w4553, IN57[12], w4655, w4656);
  FullAdder U924 (w4656, w4555, IN58[11], w4657, w4658);
  FullAdder U925 (w4658, w4557, IN59[10], w4659, w4660);
  FullAdder U926 (w4660, w4559, IN60[9], w4661, w4662);
  FullAdder U927 (w4662, w4561, IN61[8], w4663, w4664);
  FullAdder U928 (w4664, w4563, IN62[7], w4665, w4666);
  FullAdder U929 (w4666, w4565, IN63[6], w4667, w4668);
  FullAdder U930 (w4668, w4567, IN64[5], w4669, w4670);
  FullAdder U931 (w4670, w4569, IN65[4], w4671, w4672);
  FullAdder U932 (w4672, w4571, IN66[3], w4673, w4674);
  FullAdder U933 (w4674, w4573, IN67[2], w4675, w4676);
  FullAdder U934 (w4676, w4575, IN68[1], w4677, w4678);
  FullAdder U935 (w4678, w4576, IN69[0], w4679, w4680);
  HalfAdder U936 (w4579, IN19[19], Out1[19], w4682);
  FullAdder U937 (w4682, w4581, IN20[19], w4683, w4684);
  FullAdder U938 (w4684, w4583, IN21[19], w4685, w4686);
  FullAdder U939 (w4686, w4585, IN22[19], w4687, w4688);
  FullAdder U940 (w4688, w4587, IN23[19], w4689, w4690);
  FullAdder U941 (w4690, w4589, IN24[19], w4691, w4692);
  FullAdder U942 (w4692, w4591, IN25[19], w4693, w4694);
  FullAdder U943 (w4694, w4593, IN26[19], w4695, w4696);
  FullAdder U944 (w4696, w4595, IN27[19], w4697, w4698);
  FullAdder U945 (w4698, w4597, IN28[19], w4699, w4700);
  FullAdder U946 (w4700, w4599, IN29[19], w4701, w4702);
  FullAdder U947 (w4702, w4601, IN30[19], w4703, w4704);
  FullAdder U948 (w4704, w4603, IN31[19], w4705, w4706);
  FullAdder U949 (w4706, w4605, IN32[19], w4707, w4708);
  FullAdder U950 (w4708, w4607, IN33[19], w4709, w4710);
  FullAdder U951 (w4710, w4609, IN34[19], w4711, w4712);
  FullAdder U952 (w4712, w4611, IN35[19], w4713, w4714);
  FullAdder U953 (w4714, w4613, IN36[19], w4715, w4716);
  FullAdder U954 (w4716, w4615, IN37[19], w4717, w4718);
  FullAdder U955 (w4718, w4617, IN38[19], w4719, w4720);
  FullAdder U956 (w4720, w4619, IN39[19], w4721, w4722);
  FullAdder U957 (w4722, w4621, IN40[19], w4723, w4724);
  FullAdder U958 (w4724, w4623, IN41[19], w4725, w4726);
  FullAdder U959 (w4726, w4625, IN42[19], w4727, w4728);
  FullAdder U960 (w4728, w4627, IN43[19], w4729, w4730);
  FullAdder U961 (w4730, w4629, IN44[19], w4731, w4732);
  FullAdder U962 (w4732, w4631, IN45[19], w4733, w4734);
  FullAdder U963 (w4734, w4633, IN46[19], w4735, w4736);
  FullAdder U964 (w4736, w4635, IN47[19], w4737, w4738);
  FullAdder U965 (w4738, w4637, IN48[19], w4739, w4740);
  FullAdder U966 (w4740, w4639, IN49[19], w4741, w4742);
  FullAdder U967 (w4742, w4641, IN50[19], w4743, w4744);
  FullAdder U968 (w4744, w4643, IN51[19], w4745, w4746);
  FullAdder U969 (w4746, w4645, IN52[19], w4747, w4748);
  FullAdder U970 (w4748, w4647, IN53[17], w4749, w4750);
  FullAdder U971 (w4750, w4649, IN54[16], w4751, w4752);
  FullAdder U972 (w4752, w4651, IN55[15], w4753, w4754);
  FullAdder U973 (w4754, w4653, IN56[14], w4755, w4756);
  FullAdder U974 (w4756, w4655, IN57[13], w4757, w4758);
  FullAdder U975 (w4758, w4657, IN58[12], w4759, w4760);
  FullAdder U976 (w4760, w4659, IN59[11], w4761, w4762);
  FullAdder U977 (w4762, w4661, IN60[10], w4763, w4764);
  FullAdder U978 (w4764, w4663, IN61[9], w4765, w4766);
  FullAdder U979 (w4766, w4665, IN62[8], w4767, w4768);
  FullAdder U980 (w4768, w4667, IN63[7], w4769, w4770);
  FullAdder U981 (w4770, w4669, IN64[6], w4771, w4772);
  FullAdder U982 (w4772, w4671, IN65[5], w4773, w4774);
  FullAdder U983 (w4774, w4673, IN66[4], w4775, w4776);
  FullAdder U984 (w4776, w4675, IN67[3], w4777, w4778);
  FullAdder U985 (w4778, w4677, IN68[2], w4779, w4780);
  FullAdder U986 (w4780, w4679, IN69[1], w4781, w4782);
  FullAdder U987 (w4782, w4680, IN70[0], w4783, w4784);
  HalfAdder U988 (w4683, IN20[20], Out1[20], w4786);
  FullAdder U989 (w4786, w4685, IN21[20], w4787, w4788);
  FullAdder U990 (w4788, w4687, IN22[20], w4789, w4790);
  FullAdder U991 (w4790, w4689, IN23[20], w4791, w4792);
  FullAdder U992 (w4792, w4691, IN24[20], w4793, w4794);
  FullAdder U993 (w4794, w4693, IN25[20], w4795, w4796);
  FullAdder U994 (w4796, w4695, IN26[20], w4797, w4798);
  FullAdder U995 (w4798, w4697, IN27[20], w4799, w4800);
  FullAdder U996 (w4800, w4699, IN28[20], w4801, w4802);
  FullAdder U997 (w4802, w4701, IN29[20], w4803, w4804);
  FullAdder U998 (w4804, w4703, IN30[20], w4805, w4806);
  FullAdder U999 (w4806, w4705, IN31[20], w4807, w4808);
  FullAdder U1000 (w4808, w4707, IN32[20], w4809, w4810);
  FullAdder U1001 (w4810, w4709, IN33[20], w4811, w4812);
  FullAdder U1002 (w4812, w4711, IN34[20], w4813, w4814);
  FullAdder U1003 (w4814, w4713, IN35[20], w4815, w4816);
  FullAdder U1004 (w4816, w4715, IN36[20], w4817, w4818);
  FullAdder U1005 (w4818, w4717, IN37[20], w4819, w4820);
  FullAdder U1006 (w4820, w4719, IN38[20], w4821, w4822);
  FullAdder U1007 (w4822, w4721, IN39[20], w4823, w4824);
  FullAdder U1008 (w4824, w4723, IN40[20], w4825, w4826);
  FullAdder U1009 (w4826, w4725, IN41[20], w4827, w4828);
  FullAdder U1010 (w4828, w4727, IN42[20], w4829, w4830);
  FullAdder U1011 (w4830, w4729, IN43[20], w4831, w4832);
  FullAdder U1012 (w4832, w4731, IN44[20], w4833, w4834);
  FullAdder U1013 (w4834, w4733, IN45[20], w4835, w4836);
  FullAdder U1014 (w4836, w4735, IN46[20], w4837, w4838);
  FullAdder U1015 (w4838, w4737, IN47[20], w4839, w4840);
  FullAdder U1016 (w4840, w4739, IN48[20], w4841, w4842);
  FullAdder U1017 (w4842, w4741, IN49[20], w4843, w4844);
  FullAdder U1018 (w4844, w4743, IN50[20], w4845, w4846);
  FullAdder U1019 (w4846, w4745, IN51[20], w4847, w4848);
  FullAdder U1020 (w4848, w4747, IN52[20], w4849, w4850);
  FullAdder U1021 (w4850, w4749, IN53[18], w4851, w4852);
  FullAdder U1022 (w4852, w4751, IN54[17], w4853, w4854);
  FullAdder U1023 (w4854, w4753, IN55[16], w4855, w4856);
  FullAdder U1024 (w4856, w4755, IN56[15], w4857, w4858);
  FullAdder U1025 (w4858, w4757, IN57[14], w4859, w4860);
  FullAdder U1026 (w4860, w4759, IN58[13], w4861, w4862);
  FullAdder U1027 (w4862, w4761, IN59[12], w4863, w4864);
  FullAdder U1028 (w4864, w4763, IN60[11], w4865, w4866);
  FullAdder U1029 (w4866, w4765, IN61[10], w4867, w4868);
  FullAdder U1030 (w4868, w4767, IN62[9], w4869, w4870);
  FullAdder U1031 (w4870, w4769, IN63[8], w4871, w4872);
  FullAdder U1032 (w4872, w4771, IN64[7], w4873, w4874);
  FullAdder U1033 (w4874, w4773, IN65[6], w4875, w4876);
  FullAdder U1034 (w4876, w4775, IN66[5], w4877, w4878);
  FullAdder U1035 (w4878, w4777, IN67[4], w4879, w4880);
  FullAdder U1036 (w4880, w4779, IN68[3], w4881, w4882);
  FullAdder U1037 (w4882, w4781, IN69[2], w4883, w4884);
  FullAdder U1038 (w4884, w4783, IN70[1], w4885, w4886);
  FullAdder U1039 (w4886, w4784, IN71[0], w4887, w4888);
  HalfAdder U1040 (w4787, IN21[21], Out1[21], w4890);
  FullAdder U1041 (w4890, w4789, IN22[21], w4891, w4892);
  FullAdder U1042 (w4892, w4791, IN23[21], w4893, w4894);
  FullAdder U1043 (w4894, w4793, IN24[21], w4895, w4896);
  FullAdder U1044 (w4896, w4795, IN25[21], w4897, w4898);
  FullAdder U1045 (w4898, w4797, IN26[21], w4899, w4900);
  FullAdder U1046 (w4900, w4799, IN27[21], w4901, w4902);
  FullAdder U1047 (w4902, w4801, IN28[21], w4903, w4904);
  FullAdder U1048 (w4904, w4803, IN29[21], w4905, w4906);
  FullAdder U1049 (w4906, w4805, IN30[21], w4907, w4908);
  FullAdder U1050 (w4908, w4807, IN31[21], w4909, w4910);
  FullAdder U1051 (w4910, w4809, IN32[21], w4911, w4912);
  FullAdder U1052 (w4912, w4811, IN33[21], w4913, w4914);
  FullAdder U1053 (w4914, w4813, IN34[21], w4915, w4916);
  FullAdder U1054 (w4916, w4815, IN35[21], w4917, w4918);
  FullAdder U1055 (w4918, w4817, IN36[21], w4919, w4920);
  FullAdder U1056 (w4920, w4819, IN37[21], w4921, w4922);
  FullAdder U1057 (w4922, w4821, IN38[21], w4923, w4924);
  FullAdder U1058 (w4924, w4823, IN39[21], w4925, w4926);
  FullAdder U1059 (w4926, w4825, IN40[21], w4927, w4928);
  FullAdder U1060 (w4928, w4827, IN41[21], w4929, w4930);
  FullAdder U1061 (w4930, w4829, IN42[21], w4931, w4932);
  FullAdder U1062 (w4932, w4831, IN43[21], w4933, w4934);
  FullAdder U1063 (w4934, w4833, IN44[21], w4935, w4936);
  FullAdder U1064 (w4936, w4835, IN45[21], w4937, w4938);
  FullAdder U1065 (w4938, w4837, IN46[21], w4939, w4940);
  FullAdder U1066 (w4940, w4839, IN47[21], w4941, w4942);
  FullAdder U1067 (w4942, w4841, IN48[21], w4943, w4944);
  FullAdder U1068 (w4944, w4843, IN49[21], w4945, w4946);
  FullAdder U1069 (w4946, w4845, IN50[21], w4947, w4948);
  FullAdder U1070 (w4948, w4847, IN51[21], w4949, w4950);
  FullAdder U1071 (w4950, w4849, IN52[21], w4951, w4952);
  FullAdder U1072 (w4952, w4851, IN53[19], w4953, w4954);
  FullAdder U1073 (w4954, w4853, IN54[18], w4955, w4956);
  FullAdder U1074 (w4956, w4855, IN55[17], w4957, w4958);
  FullAdder U1075 (w4958, w4857, IN56[16], w4959, w4960);
  FullAdder U1076 (w4960, w4859, IN57[15], w4961, w4962);
  FullAdder U1077 (w4962, w4861, IN58[14], w4963, w4964);
  FullAdder U1078 (w4964, w4863, IN59[13], w4965, w4966);
  FullAdder U1079 (w4966, w4865, IN60[12], w4967, w4968);
  FullAdder U1080 (w4968, w4867, IN61[11], w4969, w4970);
  FullAdder U1081 (w4970, w4869, IN62[10], w4971, w4972);
  FullAdder U1082 (w4972, w4871, IN63[9], w4973, w4974);
  FullAdder U1083 (w4974, w4873, IN64[8], w4975, w4976);
  FullAdder U1084 (w4976, w4875, IN65[7], w4977, w4978);
  FullAdder U1085 (w4978, w4877, IN66[6], w4979, w4980);
  FullAdder U1086 (w4980, w4879, IN67[5], w4981, w4982);
  FullAdder U1087 (w4982, w4881, IN68[4], w4983, w4984);
  FullAdder U1088 (w4984, w4883, IN69[3], w4985, w4986);
  FullAdder U1089 (w4986, w4885, IN70[2], w4987, w4988);
  FullAdder U1090 (w4988, w4887, IN71[1], w4989, w4990);
  FullAdder U1091 (w4990, w4888, IN72[0], w4991, w4992);
  HalfAdder U1092 (w4891, IN22[22], Out1[22], w4994);
  FullAdder U1093 (w4994, w4893, IN23[22], w4995, w4996);
  FullAdder U1094 (w4996, w4895, IN24[22], w4997, w4998);
  FullAdder U1095 (w4998, w4897, IN25[22], w4999, w5000);
  FullAdder U1096 (w5000, w4899, IN26[22], w5001, w5002);
  FullAdder U1097 (w5002, w4901, IN27[22], w5003, w5004);
  FullAdder U1098 (w5004, w4903, IN28[22], w5005, w5006);
  FullAdder U1099 (w5006, w4905, IN29[22], w5007, w5008);
  FullAdder U1100 (w5008, w4907, IN30[22], w5009, w5010);
  FullAdder U1101 (w5010, w4909, IN31[22], w5011, w5012);
  FullAdder U1102 (w5012, w4911, IN32[22], w5013, w5014);
  FullAdder U1103 (w5014, w4913, IN33[22], w5015, w5016);
  FullAdder U1104 (w5016, w4915, IN34[22], w5017, w5018);
  FullAdder U1105 (w5018, w4917, IN35[22], w5019, w5020);
  FullAdder U1106 (w5020, w4919, IN36[22], w5021, w5022);
  FullAdder U1107 (w5022, w4921, IN37[22], w5023, w5024);
  FullAdder U1108 (w5024, w4923, IN38[22], w5025, w5026);
  FullAdder U1109 (w5026, w4925, IN39[22], w5027, w5028);
  FullAdder U1110 (w5028, w4927, IN40[22], w5029, w5030);
  FullAdder U1111 (w5030, w4929, IN41[22], w5031, w5032);
  FullAdder U1112 (w5032, w4931, IN42[22], w5033, w5034);
  FullAdder U1113 (w5034, w4933, IN43[22], w5035, w5036);
  FullAdder U1114 (w5036, w4935, IN44[22], w5037, w5038);
  FullAdder U1115 (w5038, w4937, IN45[22], w5039, w5040);
  FullAdder U1116 (w5040, w4939, IN46[22], w5041, w5042);
  FullAdder U1117 (w5042, w4941, IN47[22], w5043, w5044);
  FullAdder U1118 (w5044, w4943, IN48[22], w5045, w5046);
  FullAdder U1119 (w5046, w4945, IN49[22], w5047, w5048);
  FullAdder U1120 (w5048, w4947, IN50[22], w5049, w5050);
  FullAdder U1121 (w5050, w4949, IN51[22], w5051, w5052);
  FullAdder U1122 (w5052, w4951, IN52[22], w5053, w5054);
  FullAdder U1123 (w5054, w4953, IN53[20], w5055, w5056);
  FullAdder U1124 (w5056, w4955, IN54[19], w5057, w5058);
  FullAdder U1125 (w5058, w4957, IN55[18], w5059, w5060);
  FullAdder U1126 (w5060, w4959, IN56[17], w5061, w5062);
  FullAdder U1127 (w5062, w4961, IN57[16], w5063, w5064);
  FullAdder U1128 (w5064, w4963, IN58[15], w5065, w5066);
  FullAdder U1129 (w5066, w4965, IN59[14], w5067, w5068);
  FullAdder U1130 (w5068, w4967, IN60[13], w5069, w5070);
  FullAdder U1131 (w5070, w4969, IN61[12], w5071, w5072);
  FullAdder U1132 (w5072, w4971, IN62[11], w5073, w5074);
  FullAdder U1133 (w5074, w4973, IN63[10], w5075, w5076);
  FullAdder U1134 (w5076, w4975, IN64[9], w5077, w5078);
  FullAdder U1135 (w5078, w4977, IN65[8], w5079, w5080);
  FullAdder U1136 (w5080, w4979, IN66[7], w5081, w5082);
  FullAdder U1137 (w5082, w4981, IN67[6], w5083, w5084);
  FullAdder U1138 (w5084, w4983, IN68[5], w5085, w5086);
  FullAdder U1139 (w5086, w4985, IN69[4], w5087, w5088);
  FullAdder U1140 (w5088, w4987, IN70[3], w5089, w5090);
  FullAdder U1141 (w5090, w4989, IN71[2], w5091, w5092);
  FullAdder U1142 (w5092, w4991, IN72[1], w5093, w5094);
  FullAdder U1143 (w5094, w4992, IN73[0], w5095, w5096);
  HalfAdder U1144 (w4995, IN23[23], Out1[23], w5098);
  FullAdder U1145 (w5098, w4997, IN24[23], w5099, w5100);
  FullAdder U1146 (w5100, w4999, IN25[23], w5101, w5102);
  FullAdder U1147 (w5102, w5001, IN26[23], w5103, w5104);
  FullAdder U1148 (w5104, w5003, IN27[23], w5105, w5106);
  FullAdder U1149 (w5106, w5005, IN28[23], w5107, w5108);
  FullAdder U1150 (w5108, w5007, IN29[23], w5109, w5110);
  FullAdder U1151 (w5110, w5009, IN30[23], w5111, w5112);
  FullAdder U1152 (w5112, w5011, IN31[23], w5113, w5114);
  FullAdder U1153 (w5114, w5013, IN32[23], w5115, w5116);
  FullAdder U1154 (w5116, w5015, IN33[23], w5117, w5118);
  FullAdder U1155 (w5118, w5017, IN34[23], w5119, w5120);
  FullAdder U1156 (w5120, w5019, IN35[23], w5121, w5122);
  FullAdder U1157 (w5122, w5021, IN36[23], w5123, w5124);
  FullAdder U1158 (w5124, w5023, IN37[23], w5125, w5126);
  FullAdder U1159 (w5126, w5025, IN38[23], w5127, w5128);
  FullAdder U1160 (w5128, w5027, IN39[23], w5129, w5130);
  FullAdder U1161 (w5130, w5029, IN40[23], w5131, w5132);
  FullAdder U1162 (w5132, w5031, IN41[23], w5133, w5134);
  FullAdder U1163 (w5134, w5033, IN42[23], w5135, w5136);
  FullAdder U1164 (w5136, w5035, IN43[23], w5137, w5138);
  FullAdder U1165 (w5138, w5037, IN44[23], w5139, w5140);
  FullAdder U1166 (w5140, w5039, IN45[23], w5141, w5142);
  FullAdder U1167 (w5142, w5041, IN46[23], w5143, w5144);
  FullAdder U1168 (w5144, w5043, IN47[23], w5145, w5146);
  FullAdder U1169 (w5146, w5045, IN48[23], w5147, w5148);
  FullAdder U1170 (w5148, w5047, IN49[23], w5149, w5150);
  FullAdder U1171 (w5150, w5049, IN50[23], w5151, w5152);
  FullAdder U1172 (w5152, w5051, IN51[23], w5153, w5154);
  FullAdder U1173 (w5154, w5053, IN52[23], w5155, w5156);
  FullAdder U1174 (w5156, w5055, IN53[21], w5157, w5158);
  FullAdder U1175 (w5158, w5057, IN54[20], w5159, w5160);
  FullAdder U1176 (w5160, w5059, IN55[19], w5161, w5162);
  FullAdder U1177 (w5162, w5061, IN56[18], w5163, w5164);
  FullAdder U1178 (w5164, w5063, IN57[17], w5165, w5166);
  FullAdder U1179 (w5166, w5065, IN58[16], w5167, w5168);
  FullAdder U1180 (w5168, w5067, IN59[15], w5169, w5170);
  FullAdder U1181 (w5170, w5069, IN60[14], w5171, w5172);
  FullAdder U1182 (w5172, w5071, IN61[13], w5173, w5174);
  FullAdder U1183 (w5174, w5073, IN62[12], w5175, w5176);
  FullAdder U1184 (w5176, w5075, IN63[11], w5177, w5178);
  FullAdder U1185 (w5178, w5077, IN64[10], w5179, w5180);
  FullAdder U1186 (w5180, w5079, IN65[9], w5181, w5182);
  FullAdder U1187 (w5182, w5081, IN66[8], w5183, w5184);
  FullAdder U1188 (w5184, w5083, IN67[7], w5185, w5186);
  FullAdder U1189 (w5186, w5085, IN68[6], w5187, w5188);
  FullAdder U1190 (w5188, w5087, IN69[5], w5189, w5190);
  FullAdder U1191 (w5190, w5089, IN70[4], w5191, w5192);
  FullAdder U1192 (w5192, w5091, IN71[3], w5193, w5194);
  FullAdder U1193 (w5194, w5093, IN72[2], w5195, w5196);
  FullAdder U1194 (w5196, w5095, IN73[1], w5197, w5198);
  FullAdder U1195 (w5198, w5096, IN74[0], w5199, w5200);
  HalfAdder U1196 (w5099, IN24[24], Out1[24], w5202);
  FullAdder U1197 (w5202, w5101, IN25[24], w5203, w5204);
  FullAdder U1198 (w5204, w5103, IN26[24], w5205, w5206);
  FullAdder U1199 (w5206, w5105, IN27[24], w5207, w5208);
  FullAdder U1200 (w5208, w5107, IN28[24], w5209, w5210);
  FullAdder U1201 (w5210, w5109, IN29[24], w5211, w5212);
  FullAdder U1202 (w5212, w5111, IN30[24], w5213, w5214);
  FullAdder U1203 (w5214, w5113, IN31[24], w5215, w5216);
  FullAdder U1204 (w5216, w5115, IN32[24], w5217, w5218);
  FullAdder U1205 (w5218, w5117, IN33[24], w5219, w5220);
  FullAdder U1206 (w5220, w5119, IN34[24], w5221, w5222);
  FullAdder U1207 (w5222, w5121, IN35[24], w5223, w5224);
  FullAdder U1208 (w5224, w5123, IN36[24], w5225, w5226);
  FullAdder U1209 (w5226, w5125, IN37[24], w5227, w5228);
  FullAdder U1210 (w5228, w5127, IN38[24], w5229, w5230);
  FullAdder U1211 (w5230, w5129, IN39[24], w5231, w5232);
  FullAdder U1212 (w5232, w5131, IN40[24], w5233, w5234);
  FullAdder U1213 (w5234, w5133, IN41[24], w5235, w5236);
  FullAdder U1214 (w5236, w5135, IN42[24], w5237, w5238);
  FullAdder U1215 (w5238, w5137, IN43[24], w5239, w5240);
  FullAdder U1216 (w5240, w5139, IN44[24], w5241, w5242);
  FullAdder U1217 (w5242, w5141, IN45[24], w5243, w5244);
  FullAdder U1218 (w5244, w5143, IN46[24], w5245, w5246);
  FullAdder U1219 (w5246, w5145, IN47[24], w5247, w5248);
  FullAdder U1220 (w5248, w5147, IN48[24], w5249, w5250);
  FullAdder U1221 (w5250, w5149, IN49[24], w5251, w5252);
  FullAdder U1222 (w5252, w5151, IN50[24], w5253, w5254);
  FullAdder U1223 (w5254, w5153, IN51[24], w5255, w5256);
  FullAdder U1224 (w5256, w5155, IN52[24], w5257, w5258);
  FullAdder U1225 (w5258, w5157, IN53[22], w5259, w5260);
  FullAdder U1226 (w5260, w5159, IN54[21], w5261, w5262);
  FullAdder U1227 (w5262, w5161, IN55[20], w5263, w5264);
  FullAdder U1228 (w5264, w5163, IN56[19], w5265, w5266);
  FullAdder U1229 (w5266, w5165, IN57[18], w5267, w5268);
  FullAdder U1230 (w5268, w5167, IN58[17], w5269, w5270);
  FullAdder U1231 (w5270, w5169, IN59[16], w5271, w5272);
  FullAdder U1232 (w5272, w5171, IN60[15], w5273, w5274);
  FullAdder U1233 (w5274, w5173, IN61[14], w5275, w5276);
  FullAdder U1234 (w5276, w5175, IN62[13], w5277, w5278);
  FullAdder U1235 (w5278, w5177, IN63[12], w5279, w5280);
  FullAdder U1236 (w5280, w5179, IN64[11], w5281, w5282);
  FullAdder U1237 (w5282, w5181, IN65[10], w5283, w5284);
  FullAdder U1238 (w5284, w5183, IN66[9], w5285, w5286);
  FullAdder U1239 (w5286, w5185, IN67[8], w5287, w5288);
  FullAdder U1240 (w5288, w5187, IN68[7], w5289, w5290);
  FullAdder U1241 (w5290, w5189, IN69[6], w5291, w5292);
  FullAdder U1242 (w5292, w5191, IN70[5], w5293, w5294);
  FullAdder U1243 (w5294, w5193, IN71[4], w5295, w5296);
  FullAdder U1244 (w5296, w5195, IN72[3], w5297, w5298);
  FullAdder U1245 (w5298, w5197, IN73[2], w5299, w5300);
  FullAdder U1246 (w5300, w5199, IN74[1], w5301, w5302);
  FullAdder U1247 (w5302, w5200, IN75[0], w5303, w5304);
  HalfAdder U1248 (w5203, IN25[25], Out1[25], w5306);
  FullAdder U1249 (w5306, w5205, IN26[25], w5307, w5308);
  FullAdder U1250 (w5308, w5207, IN27[25], w5309, w5310);
  FullAdder U1251 (w5310, w5209, IN28[25], w5311, w5312);
  FullAdder U1252 (w5312, w5211, IN29[25], w5313, w5314);
  FullAdder U1253 (w5314, w5213, IN30[25], w5315, w5316);
  FullAdder U1254 (w5316, w5215, IN31[25], w5317, w5318);
  FullAdder U1255 (w5318, w5217, IN32[25], w5319, w5320);
  FullAdder U1256 (w5320, w5219, IN33[25], w5321, w5322);
  FullAdder U1257 (w5322, w5221, IN34[25], w5323, w5324);
  FullAdder U1258 (w5324, w5223, IN35[25], w5325, w5326);
  FullAdder U1259 (w5326, w5225, IN36[25], w5327, w5328);
  FullAdder U1260 (w5328, w5227, IN37[25], w5329, w5330);
  FullAdder U1261 (w5330, w5229, IN38[25], w5331, w5332);
  FullAdder U1262 (w5332, w5231, IN39[25], w5333, w5334);
  FullAdder U1263 (w5334, w5233, IN40[25], w5335, w5336);
  FullAdder U1264 (w5336, w5235, IN41[25], w5337, w5338);
  FullAdder U1265 (w5338, w5237, IN42[25], w5339, w5340);
  FullAdder U1266 (w5340, w5239, IN43[25], w5341, w5342);
  FullAdder U1267 (w5342, w5241, IN44[25], w5343, w5344);
  FullAdder U1268 (w5344, w5243, IN45[25], w5345, w5346);
  FullAdder U1269 (w5346, w5245, IN46[25], w5347, w5348);
  FullAdder U1270 (w5348, w5247, IN47[25], w5349, w5350);
  FullAdder U1271 (w5350, w5249, IN48[25], w5351, w5352);
  FullAdder U1272 (w5352, w5251, IN49[25], w5353, w5354);
  FullAdder U1273 (w5354, w5253, IN50[25], w5355, w5356);
  FullAdder U1274 (w5356, w5255, IN51[25], w5357, w5358);
  FullAdder U1275 (w5358, w5257, IN52[25], w5359, w5360);
  FullAdder U1276 (w5360, w5259, IN53[23], w5361, w5362);
  FullAdder U1277 (w5362, w5261, IN54[22], w5363, w5364);
  FullAdder U1278 (w5364, w5263, IN55[21], w5365, w5366);
  FullAdder U1279 (w5366, w5265, IN56[20], w5367, w5368);
  FullAdder U1280 (w5368, w5267, IN57[19], w5369, w5370);
  FullAdder U1281 (w5370, w5269, IN58[18], w5371, w5372);
  FullAdder U1282 (w5372, w5271, IN59[17], w5373, w5374);
  FullAdder U1283 (w5374, w5273, IN60[16], w5375, w5376);
  FullAdder U1284 (w5376, w5275, IN61[15], w5377, w5378);
  FullAdder U1285 (w5378, w5277, IN62[14], w5379, w5380);
  FullAdder U1286 (w5380, w5279, IN63[13], w5381, w5382);
  FullAdder U1287 (w5382, w5281, IN64[12], w5383, w5384);
  FullAdder U1288 (w5384, w5283, IN65[11], w5385, w5386);
  FullAdder U1289 (w5386, w5285, IN66[10], w5387, w5388);
  FullAdder U1290 (w5388, w5287, IN67[9], w5389, w5390);
  FullAdder U1291 (w5390, w5289, IN68[8], w5391, w5392);
  FullAdder U1292 (w5392, w5291, IN69[7], w5393, w5394);
  FullAdder U1293 (w5394, w5293, IN70[6], w5395, w5396);
  FullAdder U1294 (w5396, w5295, IN71[5], w5397, w5398);
  FullAdder U1295 (w5398, w5297, IN72[4], w5399, w5400);
  FullAdder U1296 (w5400, w5299, IN73[3], w5401, w5402);
  FullAdder U1297 (w5402, w5301, IN74[2], w5403, w5404);
  FullAdder U1298 (w5404, w5303, IN75[1], w5405, w5406);
  FullAdder U1299 (w5406, w5304, IN76[0], w5407, w5408);
  HalfAdder U1300 (w5307, IN26[26], Out1[26], w5410);
  FullAdder U1301 (w5410, w5309, IN27[26], w5411, w5412);
  FullAdder U1302 (w5412, w5311, IN28[26], w5413, w5414);
  FullAdder U1303 (w5414, w5313, IN29[26], w5415, w5416);
  FullAdder U1304 (w5416, w5315, IN30[26], w5417, w5418);
  FullAdder U1305 (w5418, w5317, IN31[26], w5419, w5420);
  FullAdder U1306 (w5420, w5319, IN32[26], w5421, w5422);
  FullAdder U1307 (w5422, w5321, IN33[26], w5423, w5424);
  FullAdder U1308 (w5424, w5323, IN34[26], w5425, w5426);
  FullAdder U1309 (w5426, w5325, IN35[26], w5427, w5428);
  FullAdder U1310 (w5428, w5327, IN36[26], w5429, w5430);
  FullAdder U1311 (w5430, w5329, IN37[26], w5431, w5432);
  FullAdder U1312 (w5432, w5331, IN38[26], w5433, w5434);
  FullAdder U1313 (w5434, w5333, IN39[26], w5435, w5436);
  FullAdder U1314 (w5436, w5335, IN40[26], w5437, w5438);
  FullAdder U1315 (w5438, w5337, IN41[26], w5439, w5440);
  FullAdder U1316 (w5440, w5339, IN42[26], w5441, w5442);
  FullAdder U1317 (w5442, w5341, IN43[26], w5443, w5444);
  FullAdder U1318 (w5444, w5343, IN44[26], w5445, w5446);
  FullAdder U1319 (w5446, w5345, IN45[26], w5447, w5448);
  FullAdder U1320 (w5448, w5347, IN46[26], w5449, w5450);
  FullAdder U1321 (w5450, w5349, IN47[26], w5451, w5452);
  FullAdder U1322 (w5452, w5351, IN48[26], w5453, w5454);
  FullAdder U1323 (w5454, w5353, IN49[26], w5455, w5456);
  FullAdder U1324 (w5456, w5355, IN50[26], w5457, w5458);
  FullAdder U1325 (w5458, w5357, IN51[26], w5459, w5460);
  FullAdder U1326 (w5460, w5359, IN52[26], w5461, w5462);
  FullAdder U1327 (w5462, w5361, IN53[24], w5463, w5464);
  FullAdder U1328 (w5464, w5363, IN54[23], w5465, w5466);
  FullAdder U1329 (w5466, w5365, IN55[22], w5467, w5468);
  FullAdder U1330 (w5468, w5367, IN56[21], w5469, w5470);
  FullAdder U1331 (w5470, w5369, IN57[20], w5471, w5472);
  FullAdder U1332 (w5472, w5371, IN58[19], w5473, w5474);
  FullAdder U1333 (w5474, w5373, IN59[18], w5475, w5476);
  FullAdder U1334 (w5476, w5375, IN60[17], w5477, w5478);
  FullAdder U1335 (w5478, w5377, IN61[16], w5479, w5480);
  FullAdder U1336 (w5480, w5379, IN62[15], w5481, w5482);
  FullAdder U1337 (w5482, w5381, IN63[14], w5483, w5484);
  FullAdder U1338 (w5484, w5383, IN64[13], w5485, w5486);
  FullAdder U1339 (w5486, w5385, IN65[12], w5487, w5488);
  FullAdder U1340 (w5488, w5387, IN66[11], w5489, w5490);
  FullAdder U1341 (w5490, w5389, IN67[10], w5491, w5492);
  FullAdder U1342 (w5492, w5391, IN68[9], w5493, w5494);
  FullAdder U1343 (w5494, w5393, IN69[8], w5495, w5496);
  FullAdder U1344 (w5496, w5395, IN70[7], w5497, w5498);
  FullAdder U1345 (w5498, w5397, IN71[6], w5499, w5500);
  FullAdder U1346 (w5500, w5399, IN72[5], w5501, w5502);
  FullAdder U1347 (w5502, w5401, IN73[4], w5503, w5504);
  FullAdder U1348 (w5504, w5403, IN74[3], w5505, w5506);
  FullAdder U1349 (w5506, w5405, IN75[2], w5507, w5508);
  FullAdder U1350 (w5508, w5407, IN76[1], w5509, w5510);
  FullAdder U1351 (w5510, w5408, IN77[0], w5511, w5512);
  HalfAdder U1352 (w5411, IN27[27], Out1[27], w5514);
  FullAdder U1353 (w5514, w5413, IN28[27], w5515, w5516);
  FullAdder U1354 (w5516, w5415, IN29[27], w5517, w5518);
  FullAdder U1355 (w5518, w5417, IN30[27], w5519, w5520);
  FullAdder U1356 (w5520, w5419, IN31[27], w5521, w5522);
  FullAdder U1357 (w5522, w5421, IN32[27], w5523, w5524);
  FullAdder U1358 (w5524, w5423, IN33[27], w5525, w5526);
  FullAdder U1359 (w5526, w5425, IN34[27], w5527, w5528);
  FullAdder U1360 (w5528, w5427, IN35[27], w5529, w5530);
  FullAdder U1361 (w5530, w5429, IN36[27], w5531, w5532);
  FullAdder U1362 (w5532, w5431, IN37[27], w5533, w5534);
  FullAdder U1363 (w5534, w5433, IN38[27], w5535, w5536);
  FullAdder U1364 (w5536, w5435, IN39[27], w5537, w5538);
  FullAdder U1365 (w5538, w5437, IN40[27], w5539, w5540);
  FullAdder U1366 (w5540, w5439, IN41[27], w5541, w5542);
  FullAdder U1367 (w5542, w5441, IN42[27], w5543, w5544);
  FullAdder U1368 (w5544, w5443, IN43[27], w5545, w5546);
  FullAdder U1369 (w5546, w5445, IN44[27], w5547, w5548);
  FullAdder U1370 (w5548, w5447, IN45[27], w5549, w5550);
  FullAdder U1371 (w5550, w5449, IN46[27], w5551, w5552);
  FullAdder U1372 (w5552, w5451, IN47[27], w5553, w5554);
  FullAdder U1373 (w5554, w5453, IN48[27], w5555, w5556);
  FullAdder U1374 (w5556, w5455, IN49[27], w5557, w5558);
  FullAdder U1375 (w5558, w5457, IN50[27], w5559, w5560);
  FullAdder U1376 (w5560, w5459, IN51[27], w5561, w5562);
  FullAdder U1377 (w5562, w5461, IN52[27], w5563, w5564);
  FullAdder U1378 (w5564, w5463, IN53[25], w5565, w5566);
  FullAdder U1379 (w5566, w5465, IN54[24], w5567, w5568);
  FullAdder U1380 (w5568, w5467, IN55[23], w5569, w5570);
  FullAdder U1381 (w5570, w5469, IN56[22], w5571, w5572);
  FullAdder U1382 (w5572, w5471, IN57[21], w5573, w5574);
  FullAdder U1383 (w5574, w5473, IN58[20], w5575, w5576);
  FullAdder U1384 (w5576, w5475, IN59[19], w5577, w5578);
  FullAdder U1385 (w5578, w5477, IN60[18], w5579, w5580);
  FullAdder U1386 (w5580, w5479, IN61[17], w5581, w5582);
  FullAdder U1387 (w5582, w5481, IN62[16], w5583, w5584);
  FullAdder U1388 (w5584, w5483, IN63[15], w5585, w5586);
  FullAdder U1389 (w5586, w5485, IN64[14], w5587, w5588);
  FullAdder U1390 (w5588, w5487, IN65[13], w5589, w5590);
  FullAdder U1391 (w5590, w5489, IN66[12], w5591, w5592);
  FullAdder U1392 (w5592, w5491, IN67[11], w5593, w5594);
  FullAdder U1393 (w5594, w5493, IN68[10], w5595, w5596);
  FullAdder U1394 (w5596, w5495, IN69[9], w5597, w5598);
  FullAdder U1395 (w5598, w5497, IN70[8], w5599, w5600);
  FullAdder U1396 (w5600, w5499, IN71[7], w5601, w5602);
  FullAdder U1397 (w5602, w5501, IN72[6], w5603, w5604);
  FullAdder U1398 (w5604, w5503, IN73[5], w5605, w5606);
  FullAdder U1399 (w5606, w5505, IN74[4], w5607, w5608);
  FullAdder U1400 (w5608, w5507, IN75[3], w5609, w5610);
  FullAdder U1401 (w5610, w5509, IN76[2], w5611, w5612);
  FullAdder U1402 (w5612, w5511, IN77[1], w5613, w5614);
  FullAdder U1403 (w5614, w5512, IN78[0], w5615, w5616);
  HalfAdder U1404 (w5515, IN28[28], Out1[28], w5618);
  FullAdder U1405 (w5618, w5517, IN29[28], w5619, w5620);
  FullAdder U1406 (w5620, w5519, IN30[28], w5621, w5622);
  FullAdder U1407 (w5622, w5521, IN31[28], w5623, w5624);
  FullAdder U1408 (w5624, w5523, IN32[28], w5625, w5626);
  FullAdder U1409 (w5626, w5525, IN33[28], w5627, w5628);
  FullAdder U1410 (w5628, w5527, IN34[28], w5629, w5630);
  FullAdder U1411 (w5630, w5529, IN35[28], w5631, w5632);
  FullAdder U1412 (w5632, w5531, IN36[28], w5633, w5634);
  FullAdder U1413 (w5634, w5533, IN37[28], w5635, w5636);
  FullAdder U1414 (w5636, w5535, IN38[28], w5637, w5638);
  FullAdder U1415 (w5638, w5537, IN39[28], w5639, w5640);
  FullAdder U1416 (w5640, w5539, IN40[28], w5641, w5642);
  FullAdder U1417 (w5642, w5541, IN41[28], w5643, w5644);
  FullAdder U1418 (w5644, w5543, IN42[28], w5645, w5646);
  FullAdder U1419 (w5646, w5545, IN43[28], w5647, w5648);
  FullAdder U1420 (w5648, w5547, IN44[28], w5649, w5650);
  FullAdder U1421 (w5650, w5549, IN45[28], w5651, w5652);
  FullAdder U1422 (w5652, w5551, IN46[28], w5653, w5654);
  FullAdder U1423 (w5654, w5553, IN47[28], w5655, w5656);
  FullAdder U1424 (w5656, w5555, IN48[28], w5657, w5658);
  FullAdder U1425 (w5658, w5557, IN49[28], w5659, w5660);
  FullAdder U1426 (w5660, w5559, IN50[28], w5661, w5662);
  FullAdder U1427 (w5662, w5561, IN51[28], w5663, w5664);
  FullAdder U1428 (w5664, w5563, IN52[28], w5665, w5666);
  FullAdder U1429 (w5666, w5565, IN53[26], w5667, w5668);
  FullAdder U1430 (w5668, w5567, IN54[25], w5669, w5670);
  FullAdder U1431 (w5670, w5569, IN55[24], w5671, w5672);
  FullAdder U1432 (w5672, w5571, IN56[23], w5673, w5674);
  FullAdder U1433 (w5674, w5573, IN57[22], w5675, w5676);
  FullAdder U1434 (w5676, w5575, IN58[21], w5677, w5678);
  FullAdder U1435 (w5678, w5577, IN59[20], w5679, w5680);
  FullAdder U1436 (w5680, w5579, IN60[19], w5681, w5682);
  FullAdder U1437 (w5682, w5581, IN61[18], w5683, w5684);
  FullAdder U1438 (w5684, w5583, IN62[17], w5685, w5686);
  FullAdder U1439 (w5686, w5585, IN63[16], w5687, w5688);
  FullAdder U1440 (w5688, w5587, IN64[15], w5689, w5690);
  FullAdder U1441 (w5690, w5589, IN65[14], w5691, w5692);
  FullAdder U1442 (w5692, w5591, IN66[13], w5693, w5694);
  FullAdder U1443 (w5694, w5593, IN67[12], w5695, w5696);
  FullAdder U1444 (w5696, w5595, IN68[11], w5697, w5698);
  FullAdder U1445 (w5698, w5597, IN69[10], w5699, w5700);
  FullAdder U1446 (w5700, w5599, IN70[9], w5701, w5702);
  FullAdder U1447 (w5702, w5601, IN71[8], w5703, w5704);
  FullAdder U1448 (w5704, w5603, IN72[7], w5705, w5706);
  FullAdder U1449 (w5706, w5605, IN73[6], w5707, w5708);
  FullAdder U1450 (w5708, w5607, IN74[5], w5709, w5710);
  FullAdder U1451 (w5710, w5609, IN75[4], w5711, w5712);
  FullAdder U1452 (w5712, w5611, IN76[3], w5713, w5714);
  FullAdder U1453 (w5714, w5613, IN77[2], w5715, w5716);
  FullAdder U1454 (w5716, w5615, IN78[1], w5717, w5718);
  FullAdder U1455 (w5718, w5616, IN79[0], w5719, w5720);
  HalfAdder U1456 (w5619, IN29[29], Out1[29], w5722);
  FullAdder U1457 (w5722, w5621, IN30[29], w5723, w5724);
  FullAdder U1458 (w5724, w5623, IN31[29], w5725, w5726);
  FullAdder U1459 (w5726, w5625, IN32[29], w5727, w5728);
  FullAdder U1460 (w5728, w5627, IN33[29], w5729, w5730);
  FullAdder U1461 (w5730, w5629, IN34[29], w5731, w5732);
  FullAdder U1462 (w5732, w5631, IN35[29], w5733, w5734);
  FullAdder U1463 (w5734, w5633, IN36[29], w5735, w5736);
  FullAdder U1464 (w5736, w5635, IN37[29], w5737, w5738);
  FullAdder U1465 (w5738, w5637, IN38[29], w5739, w5740);
  FullAdder U1466 (w5740, w5639, IN39[29], w5741, w5742);
  FullAdder U1467 (w5742, w5641, IN40[29], w5743, w5744);
  FullAdder U1468 (w5744, w5643, IN41[29], w5745, w5746);
  FullAdder U1469 (w5746, w5645, IN42[29], w5747, w5748);
  FullAdder U1470 (w5748, w5647, IN43[29], w5749, w5750);
  FullAdder U1471 (w5750, w5649, IN44[29], w5751, w5752);
  FullAdder U1472 (w5752, w5651, IN45[29], w5753, w5754);
  FullAdder U1473 (w5754, w5653, IN46[29], w5755, w5756);
  FullAdder U1474 (w5756, w5655, IN47[29], w5757, w5758);
  FullAdder U1475 (w5758, w5657, IN48[29], w5759, w5760);
  FullAdder U1476 (w5760, w5659, IN49[29], w5761, w5762);
  FullAdder U1477 (w5762, w5661, IN50[29], w5763, w5764);
  FullAdder U1478 (w5764, w5663, IN51[29], w5765, w5766);
  FullAdder U1479 (w5766, w5665, IN52[29], w5767, w5768);
  FullAdder U1480 (w5768, w5667, IN53[27], w5769, w5770);
  FullAdder U1481 (w5770, w5669, IN54[26], w5771, w5772);
  FullAdder U1482 (w5772, w5671, IN55[25], w5773, w5774);
  FullAdder U1483 (w5774, w5673, IN56[24], w5775, w5776);
  FullAdder U1484 (w5776, w5675, IN57[23], w5777, w5778);
  FullAdder U1485 (w5778, w5677, IN58[22], w5779, w5780);
  FullAdder U1486 (w5780, w5679, IN59[21], w5781, w5782);
  FullAdder U1487 (w5782, w5681, IN60[20], w5783, w5784);
  FullAdder U1488 (w5784, w5683, IN61[19], w5785, w5786);
  FullAdder U1489 (w5786, w5685, IN62[18], w5787, w5788);
  FullAdder U1490 (w5788, w5687, IN63[17], w5789, w5790);
  FullAdder U1491 (w5790, w5689, IN64[16], w5791, w5792);
  FullAdder U1492 (w5792, w5691, IN65[15], w5793, w5794);
  FullAdder U1493 (w5794, w5693, IN66[14], w5795, w5796);
  FullAdder U1494 (w5796, w5695, IN67[13], w5797, w5798);
  FullAdder U1495 (w5798, w5697, IN68[12], w5799, w5800);
  FullAdder U1496 (w5800, w5699, IN69[11], w5801, w5802);
  FullAdder U1497 (w5802, w5701, IN70[10], w5803, w5804);
  FullAdder U1498 (w5804, w5703, IN71[9], w5805, w5806);
  FullAdder U1499 (w5806, w5705, IN72[8], w5807, w5808);
  FullAdder U1500 (w5808, w5707, IN73[7], w5809, w5810);
  FullAdder U1501 (w5810, w5709, IN74[6], w5811, w5812);
  FullAdder U1502 (w5812, w5711, IN75[5], w5813, w5814);
  FullAdder U1503 (w5814, w5713, IN76[4], w5815, w5816);
  FullAdder U1504 (w5816, w5715, IN77[3], w5817, w5818);
  FullAdder U1505 (w5818, w5717, IN78[2], w5819, w5820);
  FullAdder U1506 (w5820, w5719, IN79[1], w5821, w5822);
  FullAdder U1507 (w5822, w5720, IN80[0], w5823, w5824);
  HalfAdder U1508 (w5723, IN30[30], Out1[30], w5826);
  FullAdder U1509 (w5826, w5725, IN31[30], w5827, w5828);
  FullAdder U1510 (w5828, w5727, IN32[30], w5829, w5830);
  FullAdder U1511 (w5830, w5729, IN33[30], w5831, w5832);
  FullAdder U1512 (w5832, w5731, IN34[30], w5833, w5834);
  FullAdder U1513 (w5834, w5733, IN35[30], w5835, w5836);
  FullAdder U1514 (w5836, w5735, IN36[30], w5837, w5838);
  FullAdder U1515 (w5838, w5737, IN37[30], w5839, w5840);
  FullAdder U1516 (w5840, w5739, IN38[30], w5841, w5842);
  FullAdder U1517 (w5842, w5741, IN39[30], w5843, w5844);
  FullAdder U1518 (w5844, w5743, IN40[30], w5845, w5846);
  FullAdder U1519 (w5846, w5745, IN41[30], w5847, w5848);
  FullAdder U1520 (w5848, w5747, IN42[30], w5849, w5850);
  FullAdder U1521 (w5850, w5749, IN43[30], w5851, w5852);
  FullAdder U1522 (w5852, w5751, IN44[30], w5853, w5854);
  FullAdder U1523 (w5854, w5753, IN45[30], w5855, w5856);
  FullAdder U1524 (w5856, w5755, IN46[30], w5857, w5858);
  FullAdder U1525 (w5858, w5757, IN47[30], w5859, w5860);
  FullAdder U1526 (w5860, w5759, IN48[30], w5861, w5862);
  FullAdder U1527 (w5862, w5761, IN49[30], w5863, w5864);
  FullAdder U1528 (w5864, w5763, IN50[30], w5865, w5866);
  FullAdder U1529 (w5866, w5765, IN51[30], w5867, w5868);
  FullAdder U1530 (w5868, w5767, IN52[30], w5869, w5870);
  FullAdder U1531 (w5870, w5769, IN53[28], w5871, w5872);
  FullAdder U1532 (w5872, w5771, IN54[27], w5873, w5874);
  FullAdder U1533 (w5874, w5773, IN55[26], w5875, w5876);
  FullAdder U1534 (w5876, w5775, IN56[25], w5877, w5878);
  FullAdder U1535 (w5878, w5777, IN57[24], w5879, w5880);
  FullAdder U1536 (w5880, w5779, IN58[23], w5881, w5882);
  FullAdder U1537 (w5882, w5781, IN59[22], w5883, w5884);
  FullAdder U1538 (w5884, w5783, IN60[21], w5885, w5886);
  FullAdder U1539 (w5886, w5785, IN61[20], w5887, w5888);
  FullAdder U1540 (w5888, w5787, IN62[19], w5889, w5890);
  FullAdder U1541 (w5890, w5789, IN63[18], w5891, w5892);
  FullAdder U1542 (w5892, w5791, IN64[17], w5893, w5894);
  FullAdder U1543 (w5894, w5793, IN65[16], w5895, w5896);
  FullAdder U1544 (w5896, w5795, IN66[15], w5897, w5898);
  FullAdder U1545 (w5898, w5797, IN67[14], w5899, w5900);
  FullAdder U1546 (w5900, w5799, IN68[13], w5901, w5902);
  FullAdder U1547 (w5902, w5801, IN69[12], w5903, w5904);
  FullAdder U1548 (w5904, w5803, IN70[11], w5905, w5906);
  FullAdder U1549 (w5906, w5805, IN71[10], w5907, w5908);
  FullAdder U1550 (w5908, w5807, IN72[9], w5909, w5910);
  FullAdder U1551 (w5910, w5809, IN73[8], w5911, w5912);
  FullAdder U1552 (w5912, w5811, IN74[7], w5913, w5914);
  FullAdder U1553 (w5914, w5813, IN75[6], w5915, w5916);
  FullAdder U1554 (w5916, w5815, IN76[5], w5917, w5918);
  FullAdder U1555 (w5918, w5817, IN77[4], w5919, w5920);
  FullAdder U1556 (w5920, w5819, IN78[3], w5921, w5922);
  FullAdder U1557 (w5922, w5821, IN79[2], w5923, w5924);
  FullAdder U1558 (w5924, w5823, IN80[1], w5925, w5926);
  FullAdder U1559 (w5926, w5824, IN81[0], w5927, w5928);
  HalfAdder U1560 (w5827, IN31[31], Out1[31], w5930);
  FullAdder U1561 (w5930, w5829, IN32[31], w5931, w5932);
  FullAdder U1562 (w5932, w5831, IN33[31], w5933, w5934);
  FullAdder U1563 (w5934, w5833, IN34[31], w5935, w5936);
  FullAdder U1564 (w5936, w5835, IN35[31], w5937, w5938);
  FullAdder U1565 (w5938, w5837, IN36[31], w5939, w5940);
  FullAdder U1566 (w5940, w5839, IN37[31], w5941, w5942);
  FullAdder U1567 (w5942, w5841, IN38[31], w5943, w5944);
  FullAdder U1568 (w5944, w5843, IN39[31], w5945, w5946);
  FullAdder U1569 (w5946, w5845, IN40[31], w5947, w5948);
  FullAdder U1570 (w5948, w5847, IN41[31], w5949, w5950);
  FullAdder U1571 (w5950, w5849, IN42[31], w5951, w5952);
  FullAdder U1572 (w5952, w5851, IN43[31], w5953, w5954);
  FullAdder U1573 (w5954, w5853, IN44[31], w5955, w5956);
  FullAdder U1574 (w5956, w5855, IN45[31], w5957, w5958);
  FullAdder U1575 (w5958, w5857, IN46[31], w5959, w5960);
  FullAdder U1576 (w5960, w5859, IN47[31], w5961, w5962);
  FullAdder U1577 (w5962, w5861, IN48[31], w5963, w5964);
  FullAdder U1578 (w5964, w5863, IN49[31], w5965, w5966);
  FullAdder U1579 (w5966, w5865, IN50[31], w5967, w5968);
  FullAdder U1580 (w5968, w5867, IN51[31], w5969, w5970);
  FullAdder U1581 (w5970, w5869, IN52[31], w5971, w5972);
  FullAdder U1582 (w5972, w5871, IN53[29], w5973, w5974);
  FullAdder U1583 (w5974, w5873, IN54[28], w5975, w5976);
  FullAdder U1584 (w5976, w5875, IN55[27], w5977, w5978);
  FullAdder U1585 (w5978, w5877, IN56[26], w5979, w5980);
  FullAdder U1586 (w5980, w5879, IN57[25], w5981, w5982);
  FullAdder U1587 (w5982, w5881, IN58[24], w5983, w5984);
  FullAdder U1588 (w5984, w5883, IN59[23], w5985, w5986);
  FullAdder U1589 (w5986, w5885, IN60[22], w5987, w5988);
  FullAdder U1590 (w5988, w5887, IN61[21], w5989, w5990);
  FullAdder U1591 (w5990, w5889, IN62[20], w5991, w5992);
  FullAdder U1592 (w5992, w5891, IN63[19], w5993, w5994);
  FullAdder U1593 (w5994, w5893, IN64[18], w5995, w5996);
  FullAdder U1594 (w5996, w5895, IN65[17], w5997, w5998);
  FullAdder U1595 (w5998, w5897, IN66[16], w5999, w6000);
  FullAdder U1596 (w6000, w5899, IN67[15], w6001, w6002);
  FullAdder U1597 (w6002, w5901, IN68[14], w6003, w6004);
  FullAdder U1598 (w6004, w5903, IN69[13], w6005, w6006);
  FullAdder U1599 (w6006, w5905, IN70[12], w6007, w6008);
  FullAdder U1600 (w6008, w5907, IN71[11], w6009, w6010);
  FullAdder U1601 (w6010, w5909, IN72[10], w6011, w6012);
  FullAdder U1602 (w6012, w5911, IN73[9], w6013, w6014);
  FullAdder U1603 (w6014, w5913, IN74[8], w6015, w6016);
  FullAdder U1604 (w6016, w5915, IN75[7], w6017, w6018);
  FullAdder U1605 (w6018, w5917, IN76[6], w6019, w6020);
  FullAdder U1606 (w6020, w5919, IN77[5], w6021, w6022);
  FullAdder U1607 (w6022, w5921, IN78[4], w6023, w6024);
  FullAdder U1608 (w6024, w5923, IN79[3], w6025, w6026);
  FullAdder U1609 (w6026, w5925, IN80[2], w6027, w6028);
  FullAdder U1610 (w6028, w5927, IN81[1], w6029, w6030);
  FullAdder U1611 (w6030, w5928, IN82[0], w6031, w6032);
  HalfAdder U1612 (w5931, IN32[32], Out1[32], w6034);
  FullAdder U1613 (w6034, w5933, IN33[32], w6035, w6036);
  FullAdder U1614 (w6036, w5935, IN34[32], w6037, w6038);
  FullAdder U1615 (w6038, w5937, IN35[32], w6039, w6040);
  FullAdder U1616 (w6040, w5939, IN36[32], w6041, w6042);
  FullAdder U1617 (w6042, w5941, IN37[32], w6043, w6044);
  FullAdder U1618 (w6044, w5943, IN38[32], w6045, w6046);
  FullAdder U1619 (w6046, w5945, IN39[32], w6047, w6048);
  FullAdder U1620 (w6048, w5947, IN40[32], w6049, w6050);
  FullAdder U1621 (w6050, w5949, IN41[32], w6051, w6052);
  FullAdder U1622 (w6052, w5951, IN42[32], w6053, w6054);
  FullAdder U1623 (w6054, w5953, IN43[32], w6055, w6056);
  FullAdder U1624 (w6056, w5955, IN44[32], w6057, w6058);
  FullAdder U1625 (w6058, w5957, IN45[32], w6059, w6060);
  FullAdder U1626 (w6060, w5959, IN46[32], w6061, w6062);
  FullAdder U1627 (w6062, w5961, IN47[32], w6063, w6064);
  FullAdder U1628 (w6064, w5963, IN48[32], w6065, w6066);
  FullAdder U1629 (w6066, w5965, IN49[32], w6067, w6068);
  FullAdder U1630 (w6068, w5967, IN50[32], w6069, w6070);
  FullAdder U1631 (w6070, w5969, IN51[32], w6071, w6072);
  FullAdder U1632 (w6072, w5971, IN52[32], w6073, w6074);
  FullAdder U1633 (w6074, w5973, IN53[30], w6075, w6076);
  FullAdder U1634 (w6076, w5975, IN54[29], w6077, w6078);
  FullAdder U1635 (w6078, w5977, IN55[28], w6079, w6080);
  FullAdder U1636 (w6080, w5979, IN56[27], w6081, w6082);
  FullAdder U1637 (w6082, w5981, IN57[26], w6083, w6084);
  FullAdder U1638 (w6084, w5983, IN58[25], w6085, w6086);
  FullAdder U1639 (w6086, w5985, IN59[24], w6087, w6088);
  FullAdder U1640 (w6088, w5987, IN60[23], w6089, w6090);
  FullAdder U1641 (w6090, w5989, IN61[22], w6091, w6092);
  FullAdder U1642 (w6092, w5991, IN62[21], w6093, w6094);
  FullAdder U1643 (w6094, w5993, IN63[20], w6095, w6096);
  FullAdder U1644 (w6096, w5995, IN64[19], w6097, w6098);
  FullAdder U1645 (w6098, w5997, IN65[18], w6099, w6100);
  FullAdder U1646 (w6100, w5999, IN66[17], w6101, w6102);
  FullAdder U1647 (w6102, w6001, IN67[16], w6103, w6104);
  FullAdder U1648 (w6104, w6003, IN68[15], w6105, w6106);
  FullAdder U1649 (w6106, w6005, IN69[14], w6107, w6108);
  FullAdder U1650 (w6108, w6007, IN70[13], w6109, w6110);
  FullAdder U1651 (w6110, w6009, IN71[12], w6111, w6112);
  FullAdder U1652 (w6112, w6011, IN72[11], w6113, w6114);
  FullAdder U1653 (w6114, w6013, IN73[10], w6115, w6116);
  FullAdder U1654 (w6116, w6015, IN74[9], w6117, w6118);
  FullAdder U1655 (w6118, w6017, IN75[8], w6119, w6120);
  FullAdder U1656 (w6120, w6019, IN76[7], w6121, w6122);
  FullAdder U1657 (w6122, w6021, IN77[6], w6123, w6124);
  FullAdder U1658 (w6124, w6023, IN78[5], w6125, w6126);
  FullAdder U1659 (w6126, w6025, IN79[4], w6127, w6128);
  FullAdder U1660 (w6128, w6027, IN80[3], w6129, w6130);
  FullAdder U1661 (w6130, w6029, IN81[2], w6131, w6132);
  FullAdder U1662 (w6132, w6031, IN82[1], w6133, w6134);
  FullAdder U1663 (w6134, w6032, IN83[0], w6135, w6136);
  HalfAdder U1664 (w6035, IN33[33], Out1[33], w6138);
  FullAdder U1665 (w6138, w6037, IN34[33], w6139, w6140);
  FullAdder U1666 (w6140, w6039, IN35[33], w6141, w6142);
  FullAdder U1667 (w6142, w6041, IN36[33], w6143, w6144);
  FullAdder U1668 (w6144, w6043, IN37[33], w6145, w6146);
  FullAdder U1669 (w6146, w6045, IN38[33], w6147, w6148);
  FullAdder U1670 (w6148, w6047, IN39[33], w6149, w6150);
  FullAdder U1671 (w6150, w6049, IN40[33], w6151, w6152);
  FullAdder U1672 (w6152, w6051, IN41[33], w6153, w6154);
  FullAdder U1673 (w6154, w6053, IN42[33], w6155, w6156);
  FullAdder U1674 (w6156, w6055, IN43[33], w6157, w6158);
  FullAdder U1675 (w6158, w6057, IN44[33], w6159, w6160);
  FullAdder U1676 (w6160, w6059, IN45[33], w6161, w6162);
  FullAdder U1677 (w6162, w6061, IN46[33], w6163, w6164);
  FullAdder U1678 (w6164, w6063, IN47[33], w6165, w6166);
  FullAdder U1679 (w6166, w6065, IN48[33], w6167, w6168);
  FullAdder U1680 (w6168, w6067, IN49[33], w6169, w6170);
  FullAdder U1681 (w6170, w6069, IN50[33], w6171, w6172);
  FullAdder U1682 (w6172, w6071, IN51[33], w6173, w6174);
  FullAdder U1683 (w6174, w6073, IN52[33], w6175, w6176);
  FullAdder U1684 (w6176, w6075, IN53[31], w6177, w6178);
  FullAdder U1685 (w6178, w6077, IN54[30], w6179, w6180);
  FullAdder U1686 (w6180, w6079, IN55[29], w6181, w6182);
  FullAdder U1687 (w6182, w6081, IN56[28], w6183, w6184);
  FullAdder U1688 (w6184, w6083, IN57[27], w6185, w6186);
  FullAdder U1689 (w6186, w6085, IN58[26], w6187, w6188);
  FullAdder U1690 (w6188, w6087, IN59[25], w6189, w6190);
  FullAdder U1691 (w6190, w6089, IN60[24], w6191, w6192);
  FullAdder U1692 (w6192, w6091, IN61[23], w6193, w6194);
  FullAdder U1693 (w6194, w6093, IN62[22], w6195, w6196);
  FullAdder U1694 (w6196, w6095, IN63[21], w6197, w6198);
  FullAdder U1695 (w6198, w6097, IN64[20], w6199, w6200);
  FullAdder U1696 (w6200, w6099, IN65[19], w6201, w6202);
  FullAdder U1697 (w6202, w6101, IN66[18], w6203, w6204);
  FullAdder U1698 (w6204, w6103, IN67[17], w6205, w6206);
  FullAdder U1699 (w6206, w6105, IN68[16], w6207, w6208);
  FullAdder U1700 (w6208, w6107, IN69[15], w6209, w6210);
  FullAdder U1701 (w6210, w6109, IN70[14], w6211, w6212);
  FullAdder U1702 (w6212, w6111, IN71[13], w6213, w6214);
  FullAdder U1703 (w6214, w6113, IN72[12], w6215, w6216);
  FullAdder U1704 (w6216, w6115, IN73[11], w6217, w6218);
  FullAdder U1705 (w6218, w6117, IN74[10], w6219, w6220);
  FullAdder U1706 (w6220, w6119, IN75[9], w6221, w6222);
  FullAdder U1707 (w6222, w6121, IN76[8], w6223, w6224);
  FullAdder U1708 (w6224, w6123, IN77[7], w6225, w6226);
  FullAdder U1709 (w6226, w6125, IN78[6], w6227, w6228);
  FullAdder U1710 (w6228, w6127, IN79[5], w6229, w6230);
  FullAdder U1711 (w6230, w6129, IN80[4], w6231, w6232);
  FullAdder U1712 (w6232, w6131, IN81[3], w6233, w6234);
  FullAdder U1713 (w6234, w6133, IN82[2], w6235, w6236);
  FullAdder U1714 (w6236, w6135, IN83[1], w6237, w6238);
  FullAdder U1715 (w6238, w6136, IN84[0], w6239, w6240);
  HalfAdder U1716 (w6139, IN34[34], Out1[34], w6242);
  FullAdder U1717 (w6242, w6141, IN35[34], w6243, w6244);
  FullAdder U1718 (w6244, w6143, IN36[34], w6245, w6246);
  FullAdder U1719 (w6246, w6145, IN37[34], w6247, w6248);
  FullAdder U1720 (w6248, w6147, IN38[34], w6249, w6250);
  FullAdder U1721 (w6250, w6149, IN39[34], w6251, w6252);
  FullAdder U1722 (w6252, w6151, IN40[34], w6253, w6254);
  FullAdder U1723 (w6254, w6153, IN41[34], w6255, w6256);
  FullAdder U1724 (w6256, w6155, IN42[34], w6257, w6258);
  FullAdder U1725 (w6258, w6157, IN43[34], w6259, w6260);
  FullAdder U1726 (w6260, w6159, IN44[34], w6261, w6262);
  FullAdder U1727 (w6262, w6161, IN45[34], w6263, w6264);
  FullAdder U1728 (w6264, w6163, IN46[34], w6265, w6266);
  FullAdder U1729 (w6266, w6165, IN47[34], w6267, w6268);
  FullAdder U1730 (w6268, w6167, IN48[34], w6269, w6270);
  FullAdder U1731 (w6270, w6169, IN49[34], w6271, w6272);
  FullAdder U1732 (w6272, w6171, IN50[34], w6273, w6274);
  FullAdder U1733 (w6274, w6173, IN51[34], w6275, w6276);
  FullAdder U1734 (w6276, w6175, IN52[34], w6277, w6278);
  FullAdder U1735 (w6278, w6177, IN53[32], w6279, w6280);
  FullAdder U1736 (w6280, w6179, IN54[31], w6281, w6282);
  FullAdder U1737 (w6282, w6181, IN55[30], w6283, w6284);
  FullAdder U1738 (w6284, w6183, IN56[29], w6285, w6286);
  FullAdder U1739 (w6286, w6185, IN57[28], w6287, w6288);
  FullAdder U1740 (w6288, w6187, IN58[27], w6289, w6290);
  FullAdder U1741 (w6290, w6189, IN59[26], w6291, w6292);
  FullAdder U1742 (w6292, w6191, IN60[25], w6293, w6294);
  FullAdder U1743 (w6294, w6193, IN61[24], w6295, w6296);
  FullAdder U1744 (w6296, w6195, IN62[23], w6297, w6298);
  FullAdder U1745 (w6298, w6197, IN63[22], w6299, w6300);
  FullAdder U1746 (w6300, w6199, IN64[21], w6301, w6302);
  FullAdder U1747 (w6302, w6201, IN65[20], w6303, w6304);
  FullAdder U1748 (w6304, w6203, IN66[19], w6305, w6306);
  FullAdder U1749 (w6306, w6205, IN67[18], w6307, w6308);
  FullAdder U1750 (w6308, w6207, IN68[17], w6309, w6310);
  FullAdder U1751 (w6310, w6209, IN69[16], w6311, w6312);
  FullAdder U1752 (w6312, w6211, IN70[15], w6313, w6314);
  FullAdder U1753 (w6314, w6213, IN71[14], w6315, w6316);
  FullAdder U1754 (w6316, w6215, IN72[13], w6317, w6318);
  FullAdder U1755 (w6318, w6217, IN73[12], w6319, w6320);
  FullAdder U1756 (w6320, w6219, IN74[11], w6321, w6322);
  FullAdder U1757 (w6322, w6221, IN75[10], w6323, w6324);
  FullAdder U1758 (w6324, w6223, IN76[9], w6325, w6326);
  FullAdder U1759 (w6326, w6225, IN77[8], w6327, w6328);
  FullAdder U1760 (w6328, w6227, IN78[7], w6329, w6330);
  FullAdder U1761 (w6330, w6229, IN79[6], w6331, w6332);
  FullAdder U1762 (w6332, w6231, IN80[5], w6333, w6334);
  FullAdder U1763 (w6334, w6233, IN81[4], w6335, w6336);
  FullAdder U1764 (w6336, w6235, IN82[3], w6337, w6338);
  FullAdder U1765 (w6338, w6237, IN83[2], w6339, w6340);
  FullAdder U1766 (w6340, w6239, IN84[1], w6341, w6342);
  FullAdder U1767 (w6342, w6240, IN85[0], w6343, w6344);
  HalfAdder U1768 (w6243, IN35[35], Out1[35], w6346);
  FullAdder U1769 (w6346, w6245, IN36[35], w6347, w6348);
  FullAdder U1770 (w6348, w6247, IN37[35], w6349, w6350);
  FullAdder U1771 (w6350, w6249, IN38[35], w6351, w6352);
  FullAdder U1772 (w6352, w6251, IN39[35], w6353, w6354);
  FullAdder U1773 (w6354, w6253, IN40[35], w6355, w6356);
  FullAdder U1774 (w6356, w6255, IN41[35], w6357, w6358);
  FullAdder U1775 (w6358, w6257, IN42[35], w6359, w6360);
  FullAdder U1776 (w6360, w6259, IN43[35], w6361, w6362);
  FullAdder U1777 (w6362, w6261, IN44[35], w6363, w6364);
  FullAdder U1778 (w6364, w6263, IN45[35], w6365, w6366);
  FullAdder U1779 (w6366, w6265, IN46[35], w6367, w6368);
  FullAdder U1780 (w6368, w6267, IN47[35], w6369, w6370);
  FullAdder U1781 (w6370, w6269, IN48[35], w6371, w6372);
  FullAdder U1782 (w6372, w6271, IN49[35], w6373, w6374);
  FullAdder U1783 (w6374, w6273, IN50[35], w6375, w6376);
  FullAdder U1784 (w6376, w6275, IN51[35], w6377, w6378);
  FullAdder U1785 (w6378, w6277, IN52[35], w6379, w6380);
  FullAdder U1786 (w6380, w6279, IN53[33], w6381, w6382);
  FullAdder U1787 (w6382, w6281, IN54[32], w6383, w6384);
  FullAdder U1788 (w6384, w6283, IN55[31], w6385, w6386);
  FullAdder U1789 (w6386, w6285, IN56[30], w6387, w6388);
  FullAdder U1790 (w6388, w6287, IN57[29], w6389, w6390);
  FullAdder U1791 (w6390, w6289, IN58[28], w6391, w6392);
  FullAdder U1792 (w6392, w6291, IN59[27], w6393, w6394);
  FullAdder U1793 (w6394, w6293, IN60[26], w6395, w6396);
  FullAdder U1794 (w6396, w6295, IN61[25], w6397, w6398);
  FullAdder U1795 (w6398, w6297, IN62[24], w6399, w6400);
  FullAdder U1796 (w6400, w6299, IN63[23], w6401, w6402);
  FullAdder U1797 (w6402, w6301, IN64[22], w6403, w6404);
  FullAdder U1798 (w6404, w6303, IN65[21], w6405, w6406);
  FullAdder U1799 (w6406, w6305, IN66[20], w6407, w6408);
  FullAdder U1800 (w6408, w6307, IN67[19], w6409, w6410);
  FullAdder U1801 (w6410, w6309, IN68[18], w6411, w6412);
  FullAdder U1802 (w6412, w6311, IN69[17], w6413, w6414);
  FullAdder U1803 (w6414, w6313, IN70[16], w6415, w6416);
  FullAdder U1804 (w6416, w6315, IN71[15], w6417, w6418);
  FullAdder U1805 (w6418, w6317, IN72[14], w6419, w6420);
  FullAdder U1806 (w6420, w6319, IN73[13], w6421, w6422);
  FullAdder U1807 (w6422, w6321, IN74[12], w6423, w6424);
  FullAdder U1808 (w6424, w6323, IN75[11], w6425, w6426);
  FullAdder U1809 (w6426, w6325, IN76[10], w6427, w6428);
  FullAdder U1810 (w6428, w6327, IN77[9], w6429, w6430);
  FullAdder U1811 (w6430, w6329, IN78[8], w6431, w6432);
  FullAdder U1812 (w6432, w6331, IN79[7], w6433, w6434);
  FullAdder U1813 (w6434, w6333, IN80[6], w6435, w6436);
  FullAdder U1814 (w6436, w6335, IN81[5], w6437, w6438);
  FullAdder U1815 (w6438, w6337, IN82[4], w6439, w6440);
  FullAdder U1816 (w6440, w6339, IN83[3], w6441, w6442);
  FullAdder U1817 (w6442, w6341, IN84[2], w6443, w6444);
  FullAdder U1818 (w6444, w6343, IN85[1], w6445, w6446);
  FullAdder U1819 (w6446, w6344, IN86[0], w6447, w6448);
  HalfAdder U1820 (w6347, IN36[36], Out1[36], w6450);
  FullAdder U1821 (w6450, w6349, IN37[36], w6451, w6452);
  FullAdder U1822 (w6452, w6351, IN38[36], w6453, w6454);
  FullAdder U1823 (w6454, w6353, IN39[36], w6455, w6456);
  FullAdder U1824 (w6456, w6355, IN40[36], w6457, w6458);
  FullAdder U1825 (w6458, w6357, IN41[36], w6459, w6460);
  FullAdder U1826 (w6460, w6359, IN42[36], w6461, w6462);
  FullAdder U1827 (w6462, w6361, IN43[36], w6463, w6464);
  FullAdder U1828 (w6464, w6363, IN44[36], w6465, w6466);
  FullAdder U1829 (w6466, w6365, IN45[36], w6467, w6468);
  FullAdder U1830 (w6468, w6367, IN46[36], w6469, w6470);
  FullAdder U1831 (w6470, w6369, IN47[36], w6471, w6472);
  FullAdder U1832 (w6472, w6371, IN48[36], w6473, w6474);
  FullAdder U1833 (w6474, w6373, IN49[36], w6475, w6476);
  FullAdder U1834 (w6476, w6375, IN50[36], w6477, w6478);
  FullAdder U1835 (w6478, w6377, IN51[36], w6479, w6480);
  FullAdder U1836 (w6480, w6379, IN52[36], w6481, w6482);
  FullAdder U1837 (w6482, w6381, IN53[34], w6483, w6484);
  FullAdder U1838 (w6484, w6383, IN54[33], w6485, w6486);
  FullAdder U1839 (w6486, w6385, IN55[32], w6487, w6488);
  FullAdder U1840 (w6488, w6387, IN56[31], w6489, w6490);
  FullAdder U1841 (w6490, w6389, IN57[30], w6491, w6492);
  FullAdder U1842 (w6492, w6391, IN58[29], w6493, w6494);
  FullAdder U1843 (w6494, w6393, IN59[28], w6495, w6496);
  FullAdder U1844 (w6496, w6395, IN60[27], w6497, w6498);
  FullAdder U1845 (w6498, w6397, IN61[26], w6499, w6500);
  FullAdder U1846 (w6500, w6399, IN62[25], w6501, w6502);
  FullAdder U1847 (w6502, w6401, IN63[24], w6503, w6504);
  FullAdder U1848 (w6504, w6403, IN64[23], w6505, w6506);
  FullAdder U1849 (w6506, w6405, IN65[22], w6507, w6508);
  FullAdder U1850 (w6508, w6407, IN66[21], w6509, w6510);
  FullAdder U1851 (w6510, w6409, IN67[20], w6511, w6512);
  FullAdder U1852 (w6512, w6411, IN68[19], w6513, w6514);
  FullAdder U1853 (w6514, w6413, IN69[18], w6515, w6516);
  FullAdder U1854 (w6516, w6415, IN70[17], w6517, w6518);
  FullAdder U1855 (w6518, w6417, IN71[16], w6519, w6520);
  FullAdder U1856 (w6520, w6419, IN72[15], w6521, w6522);
  FullAdder U1857 (w6522, w6421, IN73[14], w6523, w6524);
  FullAdder U1858 (w6524, w6423, IN74[13], w6525, w6526);
  FullAdder U1859 (w6526, w6425, IN75[12], w6527, w6528);
  FullAdder U1860 (w6528, w6427, IN76[11], w6529, w6530);
  FullAdder U1861 (w6530, w6429, IN77[10], w6531, w6532);
  FullAdder U1862 (w6532, w6431, IN78[9], w6533, w6534);
  FullAdder U1863 (w6534, w6433, IN79[8], w6535, w6536);
  FullAdder U1864 (w6536, w6435, IN80[7], w6537, w6538);
  FullAdder U1865 (w6538, w6437, IN81[6], w6539, w6540);
  FullAdder U1866 (w6540, w6439, IN82[5], w6541, w6542);
  FullAdder U1867 (w6542, w6441, IN83[4], w6543, w6544);
  FullAdder U1868 (w6544, w6443, IN84[3], w6545, w6546);
  FullAdder U1869 (w6546, w6445, IN85[2], w6547, w6548);
  FullAdder U1870 (w6548, w6447, IN86[1], w6549, w6550);
  FullAdder U1871 (w6550, w6448, IN87[0], w6551, w6552);
  HalfAdder U1872 (w6451, IN37[37], Out1[37], w6554);
  FullAdder U1873 (w6554, w6453, IN38[37], w6555, w6556);
  FullAdder U1874 (w6556, w6455, IN39[37], w6557, w6558);
  FullAdder U1875 (w6558, w6457, IN40[37], w6559, w6560);
  FullAdder U1876 (w6560, w6459, IN41[37], w6561, w6562);
  FullAdder U1877 (w6562, w6461, IN42[37], w6563, w6564);
  FullAdder U1878 (w6564, w6463, IN43[37], w6565, w6566);
  FullAdder U1879 (w6566, w6465, IN44[37], w6567, w6568);
  FullAdder U1880 (w6568, w6467, IN45[37], w6569, w6570);
  FullAdder U1881 (w6570, w6469, IN46[37], w6571, w6572);
  FullAdder U1882 (w6572, w6471, IN47[37], w6573, w6574);
  FullAdder U1883 (w6574, w6473, IN48[37], w6575, w6576);
  FullAdder U1884 (w6576, w6475, IN49[37], w6577, w6578);
  FullAdder U1885 (w6578, w6477, IN50[37], w6579, w6580);
  FullAdder U1886 (w6580, w6479, IN51[37], w6581, w6582);
  FullAdder U1887 (w6582, w6481, IN52[37], w6583, w6584);
  FullAdder U1888 (w6584, w6483, IN53[35], w6585, w6586);
  FullAdder U1889 (w6586, w6485, IN54[34], w6587, w6588);
  FullAdder U1890 (w6588, w6487, IN55[33], w6589, w6590);
  FullAdder U1891 (w6590, w6489, IN56[32], w6591, w6592);
  FullAdder U1892 (w6592, w6491, IN57[31], w6593, w6594);
  FullAdder U1893 (w6594, w6493, IN58[30], w6595, w6596);
  FullAdder U1894 (w6596, w6495, IN59[29], w6597, w6598);
  FullAdder U1895 (w6598, w6497, IN60[28], w6599, w6600);
  FullAdder U1896 (w6600, w6499, IN61[27], w6601, w6602);
  FullAdder U1897 (w6602, w6501, IN62[26], w6603, w6604);
  FullAdder U1898 (w6604, w6503, IN63[25], w6605, w6606);
  FullAdder U1899 (w6606, w6505, IN64[24], w6607, w6608);
  FullAdder U1900 (w6608, w6507, IN65[23], w6609, w6610);
  FullAdder U1901 (w6610, w6509, IN66[22], w6611, w6612);
  FullAdder U1902 (w6612, w6511, IN67[21], w6613, w6614);
  FullAdder U1903 (w6614, w6513, IN68[20], w6615, w6616);
  FullAdder U1904 (w6616, w6515, IN69[19], w6617, w6618);
  FullAdder U1905 (w6618, w6517, IN70[18], w6619, w6620);
  FullAdder U1906 (w6620, w6519, IN71[17], w6621, w6622);
  FullAdder U1907 (w6622, w6521, IN72[16], w6623, w6624);
  FullAdder U1908 (w6624, w6523, IN73[15], w6625, w6626);
  FullAdder U1909 (w6626, w6525, IN74[14], w6627, w6628);
  FullAdder U1910 (w6628, w6527, IN75[13], w6629, w6630);
  FullAdder U1911 (w6630, w6529, IN76[12], w6631, w6632);
  FullAdder U1912 (w6632, w6531, IN77[11], w6633, w6634);
  FullAdder U1913 (w6634, w6533, IN78[10], w6635, w6636);
  FullAdder U1914 (w6636, w6535, IN79[9], w6637, w6638);
  FullAdder U1915 (w6638, w6537, IN80[8], w6639, w6640);
  FullAdder U1916 (w6640, w6539, IN81[7], w6641, w6642);
  FullAdder U1917 (w6642, w6541, IN82[6], w6643, w6644);
  FullAdder U1918 (w6644, w6543, IN83[5], w6645, w6646);
  FullAdder U1919 (w6646, w6545, IN84[4], w6647, w6648);
  FullAdder U1920 (w6648, w6547, IN85[3], w6649, w6650);
  FullAdder U1921 (w6650, w6549, IN86[2], w6651, w6652);
  FullAdder U1922 (w6652, w6551, IN87[1], w6653, w6654);
  FullAdder U1923 (w6654, w6552, IN88[0], w6655, w6656);
  HalfAdder U1924 (w6555, IN38[38], Out1[38], w6658);
  FullAdder U1925 (w6658, w6557, IN39[38], w6659, w6660);
  FullAdder U1926 (w6660, w6559, IN40[38], w6661, w6662);
  FullAdder U1927 (w6662, w6561, IN41[38], w6663, w6664);
  FullAdder U1928 (w6664, w6563, IN42[38], w6665, w6666);
  FullAdder U1929 (w6666, w6565, IN43[38], w6667, w6668);
  FullAdder U1930 (w6668, w6567, IN44[38], w6669, w6670);
  FullAdder U1931 (w6670, w6569, IN45[38], w6671, w6672);
  FullAdder U1932 (w6672, w6571, IN46[38], w6673, w6674);
  FullAdder U1933 (w6674, w6573, IN47[38], w6675, w6676);
  FullAdder U1934 (w6676, w6575, IN48[38], w6677, w6678);
  FullAdder U1935 (w6678, w6577, IN49[38], w6679, w6680);
  FullAdder U1936 (w6680, w6579, IN50[38], w6681, w6682);
  FullAdder U1937 (w6682, w6581, IN51[38], w6683, w6684);
  FullAdder U1938 (w6684, w6583, IN52[38], w6685, w6686);
  FullAdder U1939 (w6686, w6585, IN53[36], w6687, w6688);
  FullAdder U1940 (w6688, w6587, IN54[35], w6689, w6690);
  FullAdder U1941 (w6690, w6589, IN55[34], w6691, w6692);
  FullAdder U1942 (w6692, w6591, IN56[33], w6693, w6694);
  FullAdder U1943 (w6694, w6593, IN57[32], w6695, w6696);
  FullAdder U1944 (w6696, w6595, IN58[31], w6697, w6698);
  FullAdder U1945 (w6698, w6597, IN59[30], w6699, w6700);
  FullAdder U1946 (w6700, w6599, IN60[29], w6701, w6702);
  FullAdder U1947 (w6702, w6601, IN61[28], w6703, w6704);
  FullAdder U1948 (w6704, w6603, IN62[27], w6705, w6706);
  FullAdder U1949 (w6706, w6605, IN63[26], w6707, w6708);
  FullAdder U1950 (w6708, w6607, IN64[25], w6709, w6710);
  FullAdder U1951 (w6710, w6609, IN65[24], w6711, w6712);
  FullAdder U1952 (w6712, w6611, IN66[23], w6713, w6714);
  FullAdder U1953 (w6714, w6613, IN67[22], w6715, w6716);
  FullAdder U1954 (w6716, w6615, IN68[21], w6717, w6718);
  FullAdder U1955 (w6718, w6617, IN69[20], w6719, w6720);
  FullAdder U1956 (w6720, w6619, IN70[19], w6721, w6722);
  FullAdder U1957 (w6722, w6621, IN71[18], w6723, w6724);
  FullAdder U1958 (w6724, w6623, IN72[17], w6725, w6726);
  FullAdder U1959 (w6726, w6625, IN73[16], w6727, w6728);
  FullAdder U1960 (w6728, w6627, IN74[15], w6729, w6730);
  FullAdder U1961 (w6730, w6629, IN75[14], w6731, w6732);
  FullAdder U1962 (w6732, w6631, IN76[13], w6733, w6734);
  FullAdder U1963 (w6734, w6633, IN77[12], w6735, w6736);
  FullAdder U1964 (w6736, w6635, IN78[11], w6737, w6738);
  FullAdder U1965 (w6738, w6637, IN79[10], w6739, w6740);
  FullAdder U1966 (w6740, w6639, IN80[9], w6741, w6742);
  FullAdder U1967 (w6742, w6641, IN81[8], w6743, w6744);
  FullAdder U1968 (w6744, w6643, IN82[7], w6745, w6746);
  FullAdder U1969 (w6746, w6645, IN83[6], w6747, w6748);
  FullAdder U1970 (w6748, w6647, IN84[5], w6749, w6750);
  FullAdder U1971 (w6750, w6649, IN85[4], w6751, w6752);
  FullAdder U1972 (w6752, w6651, IN86[3], w6753, w6754);
  FullAdder U1973 (w6754, w6653, IN87[2], w6755, w6756);
  FullAdder U1974 (w6756, w6655, IN88[1], w6757, w6758);
  FullAdder U1975 (w6758, w6656, IN89[0], w6759, w6760);
  HalfAdder U1976 (w6659, IN39[39], Out1[39], w6762);
  FullAdder U1977 (w6762, w6661, IN40[39], w6763, w6764);
  FullAdder U1978 (w6764, w6663, IN41[39], w6765, w6766);
  FullAdder U1979 (w6766, w6665, IN42[39], w6767, w6768);
  FullAdder U1980 (w6768, w6667, IN43[39], w6769, w6770);
  FullAdder U1981 (w6770, w6669, IN44[39], w6771, w6772);
  FullAdder U1982 (w6772, w6671, IN45[39], w6773, w6774);
  FullAdder U1983 (w6774, w6673, IN46[39], w6775, w6776);
  FullAdder U1984 (w6776, w6675, IN47[39], w6777, w6778);
  FullAdder U1985 (w6778, w6677, IN48[39], w6779, w6780);
  FullAdder U1986 (w6780, w6679, IN49[39], w6781, w6782);
  FullAdder U1987 (w6782, w6681, IN50[39], w6783, w6784);
  FullAdder U1988 (w6784, w6683, IN51[39], w6785, w6786);
  FullAdder U1989 (w6786, w6685, IN52[39], w6787, w6788);
  FullAdder U1990 (w6788, w6687, IN53[37], w6789, w6790);
  FullAdder U1991 (w6790, w6689, IN54[36], w6791, w6792);
  FullAdder U1992 (w6792, w6691, IN55[35], w6793, w6794);
  FullAdder U1993 (w6794, w6693, IN56[34], w6795, w6796);
  FullAdder U1994 (w6796, w6695, IN57[33], w6797, w6798);
  FullAdder U1995 (w6798, w6697, IN58[32], w6799, w6800);
  FullAdder U1996 (w6800, w6699, IN59[31], w6801, w6802);
  FullAdder U1997 (w6802, w6701, IN60[30], w6803, w6804);
  FullAdder U1998 (w6804, w6703, IN61[29], w6805, w6806);
  FullAdder U1999 (w6806, w6705, IN62[28], w6807, w6808);
  FullAdder U2000 (w6808, w6707, IN63[27], w6809, w6810);
  FullAdder U2001 (w6810, w6709, IN64[26], w6811, w6812);
  FullAdder U2002 (w6812, w6711, IN65[25], w6813, w6814);
  FullAdder U2003 (w6814, w6713, IN66[24], w6815, w6816);
  FullAdder U2004 (w6816, w6715, IN67[23], w6817, w6818);
  FullAdder U2005 (w6818, w6717, IN68[22], w6819, w6820);
  FullAdder U2006 (w6820, w6719, IN69[21], w6821, w6822);
  FullAdder U2007 (w6822, w6721, IN70[20], w6823, w6824);
  FullAdder U2008 (w6824, w6723, IN71[19], w6825, w6826);
  FullAdder U2009 (w6826, w6725, IN72[18], w6827, w6828);
  FullAdder U2010 (w6828, w6727, IN73[17], w6829, w6830);
  FullAdder U2011 (w6830, w6729, IN74[16], w6831, w6832);
  FullAdder U2012 (w6832, w6731, IN75[15], w6833, w6834);
  FullAdder U2013 (w6834, w6733, IN76[14], w6835, w6836);
  FullAdder U2014 (w6836, w6735, IN77[13], w6837, w6838);
  FullAdder U2015 (w6838, w6737, IN78[12], w6839, w6840);
  FullAdder U2016 (w6840, w6739, IN79[11], w6841, w6842);
  FullAdder U2017 (w6842, w6741, IN80[10], w6843, w6844);
  FullAdder U2018 (w6844, w6743, IN81[9], w6845, w6846);
  FullAdder U2019 (w6846, w6745, IN82[8], w6847, w6848);
  FullAdder U2020 (w6848, w6747, IN83[7], w6849, w6850);
  FullAdder U2021 (w6850, w6749, IN84[6], w6851, w6852);
  FullAdder U2022 (w6852, w6751, IN85[5], w6853, w6854);
  FullAdder U2023 (w6854, w6753, IN86[4], w6855, w6856);
  FullAdder U2024 (w6856, w6755, IN87[3], w6857, w6858);
  FullAdder U2025 (w6858, w6757, IN88[2], w6859, w6860);
  FullAdder U2026 (w6860, w6759, IN89[1], w6861, w6862);
  FullAdder U2027 (w6862, w6760, IN90[0], w6863, w6864);
  HalfAdder U2028 (w6763, IN40[40], Out1[40], w6866);
  FullAdder U2029 (w6866, w6765, IN41[40], w6867, w6868);
  FullAdder U2030 (w6868, w6767, IN42[40], w6869, w6870);
  FullAdder U2031 (w6870, w6769, IN43[40], w6871, w6872);
  FullAdder U2032 (w6872, w6771, IN44[40], w6873, w6874);
  FullAdder U2033 (w6874, w6773, IN45[40], w6875, w6876);
  FullAdder U2034 (w6876, w6775, IN46[40], w6877, w6878);
  FullAdder U2035 (w6878, w6777, IN47[40], w6879, w6880);
  FullAdder U2036 (w6880, w6779, IN48[40], w6881, w6882);
  FullAdder U2037 (w6882, w6781, IN49[40], w6883, w6884);
  FullAdder U2038 (w6884, w6783, IN50[40], w6885, w6886);
  FullAdder U2039 (w6886, w6785, IN51[40], w6887, w6888);
  FullAdder U2040 (w6888, w6787, IN52[40], w6889, w6890);
  FullAdder U2041 (w6890, w6789, IN53[38], w6891, w6892);
  FullAdder U2042 (w6892, w6791, IN54[37], w6893, w6894);
  FullAdder U2043 (w6894, w6793, IN55[36], w6895, w6896);
  FullAdder U2044 (w6896, w6795, IN56[35], w6897, w6898);
  FullAdder U2045 (w6898, w6797, IN57[34], w6899, w6900);
  FullAdder U2046 (w6900, w6799, IN58[33], w6901, w6902);
  FullAdder U2047 (w6902, w6801, IN59[32], w6903, w6904);
  FullAdder U2048 (w6904, w6803, IN60[31], w6905, w6906);
  FullAdder U2049 (w6906, w6805, IN61[30], w6907, w6908);
  FullAdder U2050 (w6908, w6807, IN62[29], w6909, w6910);
  FullAdder U2051 (w6910, w6809, IN63[28], w6911, w6912);
  FullAdder U2052 (w6912, w6811, IN64[27], w6913, w6914);
  FullAdder U2053 (w6914, w6813, IN65[26], w6915, w6916);
  FullAdder U2054 (w6916, w6815, IN66[25], w6917, w6918);
  FullAdder U2055 (w6918, w6817, IN67[24], w6919, w6920);
  FullAdder U2056 (w6920, w6819, IN68[23], w6921, w6922);
  FullAdder U2057 (w6922, w6821, IN69[22], w6923, w6924);
  FullAdder U2058 (w6924, w6823, IN70[21], w6925, w6926);
  FullAdder U2059 (w6926, w6825, IN71[20], w6927, w6928);
  FullAdder U2060 (w6928, w6827, IN72[19], w6929, w6930);
  FullAdder U2061 (w6930, w6829, IN73[18], w6931, w6932);
  FullAdder U2062 (w6932, w6831, IN74[17], w6933, w6934);
  FullAdder U2063 (w6934, w6833, IN75[16], w6935, w6936);
  FullAdder U2064 (w6936, w6835, IN76[15], w6937, w6938);
  FullAdder U2065 (w6938, w6837, IN77[14], w6939, w6940);
  FullAdder U2066 (w6940, w6839, IN78[13], w6941, w6942);
  FullAdder U2067 (w6942, w6841, IN79[12], w6943, w6944);
  FullAdder U2068 (w6944, w6843, IN80[11], w6945, w6946);
  FullAdder U2069 (w6946, w6845, IN81[10], w6947, w6948);
  FullAdder U2070 (w6948, w6847, IN82[9], w6949, w6950);
  FullAdder U2071 (w6950, w6849, IN83[8], w6951, w6952);
  FullAdder U2072 (w6952, w6851, IN84[7], w6953, w6954);
  FullAdder U2073 (w6954, w6853, IN85[6], w6955, w6956);
  FullAdder U2074 (w6956, w6855, IN86[5], w6957, w6958);
  FullAdder U2075 (w6958, w6857, IN87[4], w6959, w6960);
  FullAdder U2076 (w6960, w6859, IN88[3], w6961, w6962);
  FullAdder U2077 (w6962, w6861, IN89[2], w6963, w6964);
  FullAdder U2078 (w6964, w6863, IN90[1], w6965, w6966);
  FullAdder U2079 (w6966, w6864, IN91[0], w6967, w6968);
  HalfAdder U2080 (w6867, IN41[41], Out1[41], w6970);
  FullAdder U2081 (w6970, w6869, IN42[41], w6971, w6972);
  FullAdder U2082 (w6972, w6871, IN43[41], w6973, w6974);
  FullAdder U2083 (w6974, w6873, IN44[41], w6975, w6976);
  FullAdder U2084 (w6976, w6875, IN45[41], w6977, w6978);
  FullAdder U2085 (w6978, w6877, IN46[41], w6979, w6980);
  FullAdder U2086 (w6980, w6879, IN47[41], w6981, w6982);
  FullAdder U2087 (w6982, w6881, IN48[41], w6983, w6984);
  FullAdder U2088 (w6984, w6883, IN49[41], w6985, w6986);
  FullAdder U2089 (w6986, w6885, IN50[41], w6987, w6988);
  FullAdder U2090 (w6988, w6887, IN51[41], w6989, w6990);
  FullAdder U2091 (w6990, w6889, IN52[41], w6991, w6992);
  FullAdder U2092 (w6992, w6891, IN53[39], w6993, w6994);
  FullAdder U2093 (w6994, w6893, IN54[38], w6995, w6996);
  FullAdder U2094 (w6996, w6895, IN55[37], w6997, w6998);
  FullAdder U2095 (w6998, w6897, IN56[36], w6999, w7000);
  FullAdder U2096 (w7000, w6899, IN57[35], w7001, w7002);
  FullAdder U2097 (w7002, w6901, IN58[34], w7003, w7004);
  FullAdder U2098 (w7004, w6903, IN59[33], w7005, w7006);
  FullAdder U2099 (w7006, w6905, IN60[32], w7007, w7008);
  FullAdder U2100 (w7008, w6907, IN61[31], w7009, w7010);
  FullAdder U2101 (w7010, w6909, IN62[30], w7011, w7012);
  FullAdder U2102 (w7012, w6911, IN63[29], w7013, w7014);
  FullAdder U2103 (w7014, w6913, IN64[28], w7015, w7016);
  FullAdder U2104 (w7016, w6915, IN65[27], w7017, w7018);
  FullAdder U2105 (w7018, w6917, IN66[26], w7019, w7020);
  FullAdder U2106 (w7020, w6919, IN67[25], w7021, w7022);
  FullAdder U2107 (w7022, w6921, IN68[24], w7023, w7024);
  FullAdder U2108 (w7024, w6923, IN69[23], w7025, w7026);
  FullAdder U2109 (w7026, w6925, IN70[22], w7027, w7028);
  FullAdder U2110 (w7028, w6927, IN71[21], w7029, w7030);
  FullAdder U2111 (w7030, w6929, IN72[20], w7031, w7032);
  FullAdder U2112 (w7032, w6931, IN73[19], w7033, w7034);
  FullAdder U2113 (w7034, w6933, IN74[18], w7035, w7036);
  FullAdder U2114 (w7036, w6935, IN75[17], w7037, w7038);
  FullAdder U2115 (w7038, w6937, IN76[16], w7039, w7040);
  FullAdder U2116 (w7040, w6939, IN77[15], w7041, w7042);
  FullAdder U2117 (w7042, w6941, IN78[14], w7043, w7044);
  FullAdder U2118 (w7044, w6943, IN79[13], w7045, w7046);
  FullAdder U2119 (w7046, w6945, IN80[12], w7047, w7048);
  FullAdder U2120 (w7048, w6947, IN81[11], w7049, w7050);
  FullAdder U2121 (w7050, w6949, IN82[10], w7051, w7052);
  FullAdder U2122 (w7052, w6951, IN83[9], w7053, w7054);
  FullAdder U2123 (w7054, w6953, IN84[8], w7055, w7056);
  FullAdder U2124 (w7056, w6955, IN85[7], w7057, w7058);
  FullAdder U2125 (w7058, w6957, IN86[6], w7059, w7060);
  FullAdder U2126 (w7060, w6959, IN87[5], w7061, w7062);
  FullAdder U2127 (w7062, w6961, IN88[4], w7063, w7064);
  FullAdder U2128 (w7064, w6963, IN89[3], w7065, w7066);
  FullAdder U2129 (w7066, w6965, IN90[2], w7067, w7068);
  FullAdder U2130 (w7068, w6967, IN91[1], w7069, w7070);
  FullAdder U2131 (w7070, w6968, IN92[0], w7071, w7072);
  HalfAdder U2132 (w6971, IN42[42], Out1[42], w7074);
  FullAdder U2133 (w7074, w6973, IN43[42], w7075, w7076);
  FullAdder U2134 (w7076, w6975, IN44[42], w7077, w7078);
  FullAdder U2135 (w7078, w6977, IN45[42], w7079, w7080);
  FullAdder U2136 (w7080, w6979, IN46[42], w7081, w7082);
  FullAdder U2137 (w7082, w6981, IN47[42], w7083, w7084);
  FullAdder U2138 (w7084, w6983, IN48[42], w7085, w7086);
  FullAdder U2139 (w7086, w6985, IN49[42], w7087, w7088);
  FullAdder U2140 (w7088, w6987, IN50[42], w7089, w7090);
  FullAdder U2141 (w7090, w6989, IN51[42], w7091, w7092);
  FullAdder U2142 (w7092, w6991, IN52[42], w7093, w7094);
  FullAdder U2143 (w7094, w6993, IN53[40], w7095, w7096);
  FullAdder U2144 (w7096, w6995, IN54[39], w7097, w7098);
  FullAdder U2145 (w7098, w6997, IN55[38], w7099, w7100);
  FullAdder U2146 (w7100, w6999, IN56[37], w7101, w7102);
  FullAdder U2147 (w7102, w7001, IN57[36], w7103, w7104);
  FullAdder U2148 (w7104, w7003, IN58[35], w7105, w7106);
  FullAdder U2149 (w7106, w7005, IN59[34], w7107, w7108);
  FullAdder U2150 (w7108, w7007, IN60[33], w7109, w7110);
  FullAdder U2151 (w7110, w7009, IN61[32], w7111, w7112);
  FullAdder U2152 (w7112, w7011, IN62[31], w7113, w7114);
  FullAdder U2153 (w7114, w7013, IN63[30], w7115, w7116);
  FullAdder U2154 (w7116, w7015, IN64[29], w7117, w7118);
  FullAdder U2155 (w7118, w7017, IN65[28], w7119, w7120);
  FullAdder U2156 (w7120, w7019, IN66[27], w7121, w7122);
  FullAdder U2157 (w7122, w7021, IN67[26], w7123, w7124);
  FullAdder U2158 (w7124, w7023, IN68[25], w7125, w7126);
  FullAdder U2159 (w7126, w7025, IN69[24], w7127, w7128);
  FullAdder U2160 (w7128, w7027, IN70[23], w7129, w7130);
  FullAdder U2161 (w7130, w7029, IN71[22], w7131, w7132);
  FullAdder U2162 (w7132, w7031, IN72[21], w7133, w7134);
  FullAdder U2163 (w7134, w7033, IN73[20], w7135, w7136);
  FullAdder U2164 (w7136, w7035, IN74[19], w7137, w7138);
  FullAdder U2165 (w7138, w7037, IN75[18], w7139, w7140);
  FullAdder U2166 (w7140, w7039, IN76[17], w7141, w7142);
  FullAdder U2167 (w7142, w7041, IN77[16], w7143, w7144);
  FullAdder U2168 (w7144, w7043, IN78[15], w7145, w7146);
  FullAdder U2169 (w7146, w7045, IN79[14], w7147, w7148);
  FullAdder U2170 (w7148, w7047, IN80[13], w7149, w7150);
  FullAdder U2171 (w7150, w7049, IN81[12], w7151, w7152);
  FullAdder U2172 (w7152, w7051, IN82[11], w7153, w7154);
  FullAdder U2173 (w7154, w7053, IN83[10], w7155, w7156);
  FullAdder U2174 (w7156, w7055, IN84[9], w7157, w7158);
  FullAdder U2175 (w7158, w7057, IN85[8], w7159, w7160);
  FullAdder U2176 (w7160, w7059, IN86[7], w7161, w7162);
  FullAdder U2177 (w7162, w7061, IN87[6], w7163, w7164);
  FullAdder U2178 (w7164, w7063, IN88[5], w7165, w7166);
  FullAdder U2179 (w7166, w7065, IN89[4], w7167, w7168);
  FullAdder U2180 (w7168, w7067, IN90[3], w7169, w7170);
  FullAdder U2181 (w7170, w7069, IN91[2], w7171, w7172);
  FullAdder U2182 (w7172, w7071, IN92[1], w7173, w7174);
  FullAdder U2183 (w7174, w7072, IN93[0], w7175, w7176);
  HalfAdder U2184 (w7075, IN43[43], Out1[43], w7178);
  FullAdder U2185 (w7178, w7077, IN44[43], w7179, w7180);
  FullAdder U2186 (w7180, w7079, IN45[43], w7181, w7182);
  FullAdder U2187 (w7182, w7081, IN46[43], w7183, w7184);
  FullAdder U2188 (w7184, w7083, IN47[43], w7185, w7186);
  FullAdder U2189 (w7186, w7085, IN48[43], w7187, w7188);
  FullAdder U2190 (w7188, w7087, IN49[43], w7189, w7190);
  FullAdder U2191 (w7190, w7089, IN50[43], w7191, w7192);
  FullAdder U2192 (w7192, w7091, IN51[43], w7193, w7194);
  FullAdder U2193 (w7194, w7093, IN52[43], w7195, w7196);
  FullAdder U2194 (w7196, w7095, IN53[41], w7197, w7198);
  FullAdder U2195 (w7198, w7097, IN54[40], w7199, w7200);
  FullAdder U2196 (w7200, w7099, IN55[39], w7201, w7202);
  FullAdder U2197 (w7202, w7101, IN56[38], w7203, w7204);
  FullAdder U2198 (w7204, w7103, IN57[37], w7205, w7206);
  FullAdder U2199 (w7206, w7105, IN58[36], w7207, w7208);
  FullAdder U2200 (w7208, w7107, IN59[35], w7209, w7210);
  FullAdder U2201 (w7210, w7109, IN60[34], w7211, w7212);
  FullAdder U2202 (w7212, w7111, IN61[33], w7213, w7214);
  FullAdder U2203 (w7214, w7113, IN62[32], w7215, w7216);
  FullAdder U2204 (w7216, w7115, IN63[31], w7217, w7218);
  FullAdder U2205 (w7218, w7117, IN64[30], w7219, w7220);
  FullAdder U2206 (w7220, w7119, IN65[29], w7221, w7222);
  FullAdder U2207 (w7222, w7121, IN66[28], w7223, w7224);
  FullAdder U2208 (w7224, w7123, IN67[27], w7225, w7226);
  FullAdder U2209 (w7226, w7125, IN68[26], w7227, w7228);
  FullAdder U2210 (w7228, w7127, IN69[25], w7229, w7230);
  FullAdder U2211 (w7230, w7129, IN70[24], w7231, w7232);
  FullAdder U2212 (w7232, w7131, IN71[23], w7233, w7234);
  FullAdder U2213 (w7234, w7133, IN72[22], w7235, w7236);
  FullAdder U2214 (w7236, w7135, IN73[21], w7237, w7238);
  FullAdder U2215 (w7238, w7137, IN74[20], w7239, w7240);
  FullAdder U2216 (w7240, w7139, IN75[19], w7241, w7242);
  FullAdder U2217 (w7242, w7141, IN76[18], w7243, w7244);
  FullAdder U2218 (w7244, w7143, IN77[17], w7245, w7246);
  FullAdder U2219 (w7246, w7145, IN78[16], w7247, w7248);
  FullAdder U2220 (w7248, w7147, IN79[15], w7249, w7250);
  FullAdder U2221 (w7250, w7149, IN80[14], w7251, w7252);
  FullAdder U2222 (w7252, w7151, IN81[13], w7253, w7254);
  FullAdder U2223 (w7254, w7153, IN82[12], w7255, w7256);
  FullAdder U2224 (w7256, w7155, IN83[11], w7257, w7258);
  FullAdder U2225 (w7258, w7157, IN84[10], w7259, w7260);
  FullAdder U2226 (w7260, w7159, IN85[9], w7261, w7262);
  FullAdder U2227 (w7262, w7161, IN86[8], w7263, w7264);
  FullAdder U2228 (w7264, w7163, IN87[7], w7265, w7266);
  FullAdder U2229 (w7266, w7165, IN88[6], w7267, w7268);
  FullAdder U2230 (w7268, w7167, IN89[5], w7269, w7270);
  FullAdder U2231 (w7270, w7169, IN90[4], w7271, w7272);
  FullAdder U2232 (w7272, w7171, IN91[3], w7273, w7274);
  FullAdder U2233 (w7274, w7173, IN92[2], w7275, w7276);
  FullAdder U2234 (w7276, w7175, IN93[1], w7277, w7278);
  FullAdder U2235 (w7278, w7176, IN94[0], w7279, w7280);
  HalfAdder U2236 (w7179, IN44[44], Out1[44], w7282);
  FullAdder U2237 (w7282, w7181, IN45[44], w7283, w7284);
  FullAdder U2238 (w7284, w7183, IN46[44], w7285, w7286);
  FullAdder U2239 (w7286, w7185, IN47[44], w7287, w7288);
  FullAdder U2240 (w7288, w7187, IN48[44], w7289, w7290);
  FullAdder U2241 (w7290, w7189, IN49[44], w7291, w7292);
  FullAdder U2242 (w7292, w7191, IN50[44], w7293, w7294);
  FullAdder U2243 (w7294, w7193, IN51[44], w7295, w7296);
  FullAdder U2244 (w7296, w7195, IN52[44], w7297, w7298);
  FullAdder U2245 (w7298, w7197, IN53[42], w7299, w7300);
  FullAdder U2246 (w7300, w7199, IN54[41], w7301, w7302);
  FullAdder U2247 (w7302, w7201, IN55[40], w7303, w7304);
  FullAdder U2248 (w7304, w7203, IN56[39], w7305, w7306);
  FullAdder U2249 (w7306, w7205, IN57[38], w7307, w7308);
  FullAdder U2250 (w7308, w7207, IN58[37], w7309, w7310);
  FullAdder U2251 (w7310, w7209, IN59[36], w7311, w7312);
  FullAdder U2252 (w7312, w7211, IN60[35], w7313, w7314);
  FullAdder U2253 (w7314, w7213, IN61[34], w7315, w7316);
  FullAdder U2254 (w7316, w7215, IN62[33], w7317, w7318);
  FullAdder U2255 (w7318, w7217, IN63[32], w7319, w7320);
  FullAdder U2256 (w7320, w7219, IN64[31], w7321, w7322);
  FullAdder U2257 (w7322, w7221, IN65[30], w7323, w7324);
  FullAdder U2258 (w7324, w7223, IN66[29], w7325, w7326);
  FullAdder U2259 (w7326, w7225, IN67[28], w7327, w7328);
  FullAdder U2260 (w7328, w7227, IN68[27], w7329, w7330);
  FullAdder U2261 (w7330, w7229, IN69[26], w7331, w7332);
  FullAdder U2262 (w7332, w7231, IN70[25], w7333, w7334);
  FullAdder U2263 (w7334, w7233, IN71[24], w7335, w7336);
  FullAdder U2264 (w7336, w7235, IN72[23], w7337, w7338);
  FullAdder U2265 (w7338, w7237, IN73[22], w7339, w7340);
  FullAdder U2266 (w7340, w7239, IN74[21], w7341, w7342);
  FullAdder U2267 (w7342, w7241, IN75[20], w7343, w7344);
  FullAdder U2268 (w7344, w7243, IN76[19], w7345, w7346);
  FullAdder U2269 (w7346, w7245, IN77[18], w7347, w7348);
  FullAdder U2270 (w7348, w7247, IN78[17], w7349, w7350);
  FullAdder U2271 (w7350, w7249, IN79[16], w7351, w7352);
  FullAdder U2272 (w7352, w7251, IN80[15], w7353, w7354);
  FullAdder U2273 (w7354, w7253, IN81[14], w7355, w7356);
  FullAdder U2274 (w7356, w7255, IN82[13], w7357, w7358);
  FullAdder U2275 (w7358, w7257, IN83[12], w7359, w7360);
  FullAdder U2276 (w7360, w7259, IN84[11], w7361, w7362);
  FullAdder U2277 (w7362, w7261, IN85[10], w7363, w7364);
  FullAdder U2278 (w7364, w7263, IN86[9], w7365, w7366);
  FullAdder U2279 (w7366, w7265, IN87[8], w7367, w7368);
  FullAdder U2280 (w7368, w7267, IN88[7], w7369, w7370);
  FullAdder U2281 (w7370, w7269, IN89[6], w7371, w7372);
  FullAdder U2282 (w7372, w7271, IN90[5], w7373, w7374);
  FullAdder U2283 (w7374, w7273, IN91[4], w7375, w7376);
  FullAdder U2284 (w7376, w7275, IN92[3], w7377, w7378);
  FullAdder U2285 (w7378, w7277, IN93[2], w7379, w7380);
  FullAdder U2286 (w7380, w7279, IN94[1], w7381, w7382);
  FullAdder U2287 (w7382, w7280, IN95[0], w7383, w7384);
  HalfAdder U2288 (w7283, IN45[45], Out1[45], w7386);
  FullAdder U2289 (w7386, w7285, IN46[45], w7387, w7388);
  FullAdder U2290 (w7388, w7287, IN47[45], w7389, w7390);
  FullAdder U2291 (w7390, w7289, IN48[45], w7391, w7392);
  FullAdder U2292 (w7392, w7291, IN49[45], w7393, w7394);
  FullAdder U2293 (w7394, w7293, IN50[45], w7395, w7396);
  FullAdder U2294 (w7396, w7295, IN51[45], w7397, w7398);
  FullAdder U2295 (w7398, w7297, IN52[45], w7399, w7400);
  FullAdder U2296 (w7400, w7299, IN53[43], w7401, w7402);
  FullAdder U2297 (w7402, w7301, IN54[42], w7403, w7404);
  FullAdder U2298 (w7404, w7303, IN55[41], w7405, w7406);
  FullAdder U2299 (w7406, w7305, IN56[40], w7407, w7408);
  FullAdder U2300 (w7408, w7307, IN57[39], w7409, w7410);
  FullAdder U2301 (w7410, w7309, IN58[38], w7411, w7412);
  FullAdder U2302 (w7412, w7311, IN59[37], w7413, w7414);
  FullAdder U2303 (w7414, w7313, IN60[36], w7415, w7416);
  FullAdder U2304 (w7416, w7315, IN61[35], w7417, w7418);
  FullAdder U2305 (w7418, w7317, IN62[34], w7419, w7420);
  FullAdder U2306 (w7420, w7319, IN63[33], w7421, w7422);
  FullAdder U2307 (w7422, w7321, IN64[32], w7423, w7424);
  FullAdder U2308 (w7424, w7323, IN65[31], w7425, w7426);
  FullAdder U2309 (w7426, w7325, IN66[30], w7427, w7428);
  FullAdder U2310 (w7428, w7327, IN67[29], w7429, w7430);
  FullAdder U2311 (w7430, w7329, IN68[28], w7431, w7432);
  FullAdder U2312 (w7432, w7331, IN69[27], w7433, w7434);
  FullAdder U2313 (w7434, w7333, IN70[26], w7435, w7436);
  FullAdder U2314 (w7436, w7335, IN71[25], w7437, w7438);
  FullAdder U2315 (w7438, w7337, IN72[24], w7439, w7440);
  FullAdder U2316 (w7440, w7339, IN73[23], w7441, w7442);
  FullAdder U2317 (w7442, w7341, IN74[22], w7443, w7444);
  FullAdder U2318 (w7444, w7343, IN75[21], w7445, w7446);
  FullAdder U2319 (w7446, w7345, IN76[20], w7447, w7448);
  FullAdder U2320 (w7448, w7347, IN77[19], w7449, w7450);
  FullAdder U2321 (w7450, w7349, IN78[18], w7451, w7452);
  FullAdder U2322 (w7452, w7351, IN79[17], w7453, w7454);
  FullAdder U2323 (w7454, w7353, IN80[16], w7455, w7456);
  FullAdder U2324 (w7456, w7355, IN81[15], w7457, w7458);
  FullAdder U2325 (w7458, w7357, IN82[14], w7459, w7460);
  FullAdder U2326 (w7460, w7359, IN83[13], w7461, w7462);
  FullAdder U2327 (w7462, w7361, IN84[12], w7463, w7464);
  FullAdder U2328 (w7464, w7363, IN85[11], w7465, w7466);
  FullAdder U2329 (w7466, w7365, IN86[10], w7467, w7468);
  FullAdder U2330 (w7468, w7367, IN87[9], w7469, w7470);
  FullAdder U2331 (w7470, w7369, IN88[8], w7471, w7472);
  FullAdder U2332 (w7472, w7371, IN89[7], w7473, w7474);
  FullAdder U2333 (w7474, w7373, IN90[6], w7475, w7476);
  FullAdder U2334 (w7476, w7375, IN91[5], w7477, w7478);
  FullAdder U2335 (w7478, w7377, IN92[4], w7479, w7480);
  FullAdder U2336 (w7480, w7379, IN93[3], w7481, w7482);
  FullAdder U2337 (w7482, w7381, IN94[2], w7483, w7484);
  FullAdder U2338 (w7484, w7383, IN95[1], w7485, w7486);
  FullAdder U2339 (w7486, w7384, IN96[0], w7487, w7488);
  HalfAdder U2340 (w7387, IN46[46], Out1[46], w7490);
  FullAdder U2341 (w7490, w7389, IN47[46], w7491, w7492);
  FullAdder U2342 (w7492, w7391, IN48[46], w7493, w7494);
  FullAdder U2343 (w7494, w7393, IN49[46], w7495, w7496);
  FullAdder U2344 (w7496, w7395, IN50[46], w7497, w7498);
  FullAdder U2345 (w7498, w7397, IN51[46], w7499, w7500);
  FullAdder U2346 (w7500, w7399, IN52[46], w7501, w7502);
  FullAdder U2347 (w7502, w7401, IN53[44], w7503, w7504);
  FullAdder U2348 (w7504, w7403, IN54[43], w7505, w7506);
  FullAdder U2349 (w7506, w7405, IN55[42], w7507, w7508);
  FullAdder U2350 (w7508, w7407, IN56[41], w7509, w7510);
  FullAdder U2351 (w7510, w7409, IN57[40], w7511, w7512);
  FullAdder U2352 (w7512, w7411, IN58[39], w7513, w7514);
  FullAdder U2353 (w7514, w7413, IN59[38], w7515, w7516);
  FullAdder U2354 (w7516, w7415, IN60[37], w7517, w7518);
  FullAdder U2355 (w7518, w7417, IN61[36], w7519, w7520);
  FullAdder U2356 (w7520, w7419, IN62[35], w7521, w7522);
  FullAdder U2357 (w7522, w7421, IN63[34], w7523, w7524);
  FullAdder U2358 (w7524, w7423, IN64[33], w7525, w7526);
  FullAdder U2359 (w7526, w7425, IN65[32], w7527, w7528);
  FullAdder U2360 (w7528, w7427, IN66[31], w7529, w7530);
  FullAdder U2361 (w7530, w7429, IN67[30], w7531, w7532);
  FullAdder U2362 (w7532, w7431, IN68[29], w7533, w7534);
  FullAdder U2363 (w7534, w7433, IN69[28], w7535, w7536);
  FullAdder U2364 (w7536, w7435, IN70[27], w7537, w7538);
  FullAdder U2365 (w7538, w7437, IN71[26], w7539, w7540);
  FullAdder U2366 (w7540, w7439, IN72[25], w7541, w7542);
  FullAdder U2367 (w7542, w7441, IN73[24], w7543, w7544);
  FullAdder U2368 (w7544, w7443, IN74[23], w7545, w7546);
  FullAdder U2369 (w7546, w7445, IN75[22], w7547, w7548);
  FullAdder U2370 (w7548, w7447, IN76[21], w7549, w7550);
  FullAdder U2371 (w7550, w7449, IN77[20], w7551, w7552);
  FullAdder U2372 (w7552, w7451, IN78[19], w7553, w7554);
  FullAdder U2373 (w7554, w7453, IN79[18], w7555, w7556);
  FullAdder U2374 (w7556, w7455, IN80[17], w7557, w7558);
  FullAdder U2375 (w7558, w7457, IN81[16], w7559, w7560);
  FullAdder U2376 (w7560, w7459, IN82[15], w7561, w7562);
  FullAdder U2377 (w7562, w7461, IN83[14], w7563, w7564);
  FullAdder U2378 (w7564, w7463, IN84[13], w7565, w7566);
  FullAdder U2379 (w7566, w7465, IN85[12], w7567, w7568);
  FullAdder U2380 (w7568, w7467, IN86[11], w7569, w7570);
  FullAdder U2381 (w7570, w7469, IN87[10], w7571, w7572);
  FullAdder U2382 (w7572, w7471, IN88[9], w7573, w7574);
  FullAdder U2383 (w7574, w7473, IN89[8], w7575, w7576);
  FullAdder U2384 (w7576, w7475, IN90[7], w7577, w7578);
  FullAdder U2385 (w7578, w7477, IN91[6], w7579, w7580);
  FullAdder U2386 (w7580, w7479, IN92[5], w7581, w7582);
  FullAdder U2387 (w7582, w7481, IN93[4], w7583, w7584);
  FullAdder U2388 (w7584, w7483, IN94[3], w7585, w7586);
  FullAdder U2389 (w7586, w7485, IN95[2], w7587, w7588);
  FullAdder U2390 (w7588, w7487, IN96[1], w7589, w7590);
  FullAdder U2391 (w7590, w7488, IN97[0], w7591, w7592);
  HalfAdder U2392 (w7491, IN47[47], Out1[47], w7594);
  FullAdder U2393 (w7594, w7493, IN48[47], w7595, w7596);
  FullAdder U2394 (w7596, w7495, IN49[47], w7597, w7598);
  FullAdder U2395 (w7598, w7497, IN50[47], w7599, w7600);
  FullAdder U2396 (w7600, w7499, IN51[47], w7601, w7602);
  FullAdder U2397 (w7602, w7501, IN52[47], w7603, w7604);
  FullAdder U2398 (w7604, w7503, IN53[45], w7605, w7606);
  FullAdder U2399 (w7606, w7505, IN54[44], w7607, w7608);
  FullAdder U2400 (w7608, w7507, IN55[43], w7609, w7610);
  FullAdder U2401 (w7610, w7509, IN56[42], w7611, w7612);
  FullAdder U2402 (w7612, w7511, IN57[41], w7613, w7614);
  FullAdder U2403 (w7614, w7513, IN58[40], w7615, w7616);
  FullAdder U2404 (w7616, w7515, IN59[39], w7617, w7618);
  FullAdder U2405 (w7618, w7517, IN60[38], w7619, w7620);
  FullAdder U2406 (w7620, w7519, IN61[37], w7621, w7622);
  FullAdder U2407 (w7622, w7521, IN62[36], w7623, w7624);
  FullAdder U2408 (w7624, w7523, IN63[35], w7625, w7626);
  FullAdder U2409 (w7626, w7525, IN64[34], w7627, w7628);
  FullAdder U2410 (w7628, w7527, IN65[33], w7629, w7630);
  FullAdder U2411 (w7630, w7529, IN66[32], w7631, w7632);
  FullAdder U2412 (w7632, w7531, IN67[31], w7633, w7634);
  FullAdder U2413 (w7634, w7533, IN68[30], w7635, w7636);
  FullAdder U2414 (w7636, w7535, IN69[29], w7637, w7638);
  FullAdder U2415 (w7638, w7537, IN70[28], w7639, w7640);
  FullAdder U2416 (w7640, w7539, IN71[27], w7641, w7642);
  FullAdder U2417 (w7642, w7541, IN72[26], w7643, w7644);
  FullAdder U2418 (w7644, w7543, IN73[25], w7645, w7646);
  FullAdder U2419 (w7646, w7545, IN74[24], w7647, w7648);
  FullAdder U2420 (w7648, w7547, IN75[23], w7649, w7650);
  FullAdder U2421 (w7650, w7549, IN76[22], w7651, w7652);
  FullAdder U2422 (w7652, w7551, IN77[21], w7653, w7654);
  FullAdder U2423 (w7654, w7553, IN78[20], w7655, w7656);
  FullAdder U2424 (w7656, w7555, IN79[19], w7657, w7658);
  FullAdder U2425 (w7658, w7557, IN80[18], w7659, w7660);
  FullAdder U2426 (w7660, w7559, IN81[17], w7661, w7662);
  FullAdder U2427 (w7662, w7561, IN82[16], w7663, w7664);
  FullAdder U2428 (w7664, w7563, IN83[15], w7665, w7666);
  FullAdder U2429 (w7666, w7565, IN84[14], w7667, w7668);
  FullAdder U2430 (w7668, w7567, IN85[13], w7669, w7670);
  FullAdder U2431 (w7670, w7569, IN86[12], w7671, w7672);
  FullAdder U2432 (w7672, w7571, IN87[11], w7673, w7674);
  FullAdder U2433 (w7674, w7573, IN88[10], w7675, w7676);
  FullAdder U2434 (w7676, w7575, IN89[9], w7677, w7678);
  FullAdder U2435 (w7678, w7577, IN90[8], w7679, w7680);
  FullAdder U2436 (w7680, w7579, IN91[7], w7681, w7682);
  FullAdder U2437 (w7682, w7581, IN92[6], w7683, w7684);
  FullAdder U2438 (w7684, w7583, IN93[5], w7685, w7686);
  FullAdder U2439 (w7686, w7585, IN94[4], w7687, w7688);
  FullAdder U2440 (w7688, w7587, IN95[3], w7689, w7690);
  FullAdder U2441 (w7690, w7589, IN96[2], w7691, w7692);
  FullAdder U2442 (w7692, w7591, IN97[1], w7693, w7694);
  FullAdder U2443 (w7694, w7592, IN98[0], w7695, w7696);
  HalfAdder U2444 (w7595, IN48[48], Out1[48], w7698);
  FullAdder U2445 (w7698, w7597, IN49[48], w7699, w7700);
  FullAdder U2446 (w7700, w7599, IN50[48], w7701, w7702);
  FullAdder U2447 (w7702, w7601, IN51[48], w7703, w7704);
  FullAdder U2448 (w7704, w7603, IN52[48], w7705, w7706);
  FullAdder U2449 (w7706, w7605, IN53[46], w7707, w7708);
  FullAdder U2450 (w7708, w7607, IN54[45], w7709, w7710);
  FullAdder U2451 (w7710, w7609, IN55[44], w7711, w7712);
  FullAdder U2452 (w7712, w7611, IN56[43], w7713, w7714);
  FullAdder U2453 (w7714, w7613, IN57[42], w7715, w7716);
  FullAdder U2454 (w7716, w7615, IN58[41], w7717, w7718);
  FullAdder U2455 (w7718, w7617, IN59[40], w7719, w7720);
  FullAdder U2456 (w7720, w7619, IN60[39], w7721, w7722);
  FullAdder U2457 (w7722, w7621, IN61[38], w7723, w7724);
  FullAdder U2458 (w7724, w7623, IN62[37], w7725, w7726);
  FullAdder U2459 (w7726, w7625, IN63[36], w7727, w7728);
  FullAdder U2460 (w7728, w7627, IN64[35], w7729, w7730);
  FullAdder U2461 (w7730, w7629, IN65[34], w7731, w7732);
  FullAdder U2462 (w7732, w7631, IN66[33], w7733, w7734);
  FullAdder U2463 (w7734, w7633, IN67[32], w7735, w7736);
  FullAdder U2464 (w7736, w7635, IN68[31], w7737, w7738);
  FullAdder U2465 (w7738, w7637, IN69[30], w7739, w7740);
  FullAdder U2466 (w7740, w7639, IN70[29], w7741, w7742);
  FullAdder U2467 (w7742, w7641, IN71[28], w7743, w7744);
  FullAdder U2468 (w7744, w7643, IN72[27], w7745, w7746);
  FullAdder U2469 (w7746, w7645, IN73[26], w7747, w7748);
  FullAdder U2470 (w7748, w7647, IN74[25], w7749, w7750);
  FullAdder U2471 (w7750, w7649, IN75[24], w7751, w7752);
  FullAdder U2472 (w7752, w7651, IN76[23], w7753, w7754);
  FullAdder U2473 (w7754, w7653, IN77[22], w7755, w7756);
  FullAdder U2474 (w7756, w7655, IN78[21], w7757, w7758);
  FullAdder U2475 (w7758, w7657, IN79[20], w7759, w7760);
  FullAdder U2476 (w7760, w7659, IN80[19], w7761, w7762);
  FullAdder U2477 (w7762, w7661, IN81[18], w7763, w7764);
  FullAdder U2478 (w7764, w7663, IN82[17], w7765, w7766);
  FullAdder U2479 (w7766, w7665, IN83[16], w7767, w7768);
  FullAdder U2480 (w7768, w7667, IN84[15], w7769, w7770);
  FullAdder U2481 (w7770, w7669, IN85[14], w7771, w7772);
  FullAdder U2482 (w7772, w7671, IN86[13], w7773, w7774);
  FullAdder U2483 (w7774, w7673, IN87[12], w7775, w7776);
  FullAdder U2484 (w7776, w7675, IN88[11], w7777, w7778);
  FullAdder U2485 (w7778, w7677, IN89[10], w7779, w7780);
  FullAdder U2486 (w7780, w7679, IN90[9], w7781, w7782);
  FullAdder U2487 (w7782, w7681, IN91[8], w7783, w7784);
  FullAdder U2488 (w7784, w7683, IN92[7], w7785, w7786);
  FullAdder U2489 (w7786, w7685, IN93[6], w7787, w7788);
  FullAdder U2490 (w7788, w7687, IN94[5], w7789, w7790);
  FullAdder U2491 (w7790, w7689, IN95[4], w7791, w7792);
  FullAdder U2492 (w7792, w7691, IN96[3], w7793, w7794);
  FullAdder U2493 (w7794, w7693, IN97[2], w7795, w7796);
  FullAdder U2494 (w7796, w7695, IN98[1], w7797, w7798);
  FullAdder U2495 (w7798, w7696, IN99[0], w7799, w7800);
  HalfAdder U2496 (w7699, IN49[49], Out1[49], w7802);
  FullAdder U2497 (w7802, w7701, IN50[49], w7803, w7804);
  FullAdder U2498 (w7804, w7703, IN51[49], w7805, w7806);
  FullAdder U2499 (w7806, w7705, IN52[49], w7807, w7808);
  FullAdder U2500 (w7808, w7707, IN53[47], w7809, w7810);
  FullAdder U2501 (w7810, w7709, IN54[46], w7811, w7812);
  FullAdder U2502 (w7812, w7711, IN55[45], w7813, w7814);
  FullAdder U2503 (w7814, w7713, IN56[44], w7815, w7816);
  FullAdder U2504 (w7816, w7715, IN57[43], w7817, w7818);
  FullAdder U2505 (w7818, w7717, IN58[42], w7819, w7820);
  FullAdder U2506 (w7820, w7719, IN59[41], w7821, w7822);
  FullAdder U2507 (w7822, w7721, IN60[40], w7823, w7824);
  FullAdder U2508 (w7824, w7723, IN61[39], w7825, w7826);
  FullAdder U2509 (w7826, w7725, IN62[38], w7827, w7828);
  FullAdder U2510 (w7828, w7727, IN63[37], w7829, w7830);
  FullAdder U2511 (w7830, w7729, IN64[36], w7831, w7832);
  FullAdder U2512 (w7832, w7731, IN65[35], w7833, w7834);
  FullAdder U2513 (w7834, w7733, IN66[34], w7835, w7836);
  FullAdder U2514 (w7836, w7735, IN67[33], w7837, w7838);
  FullAdder U2515 (w7838, w7737, IN68[32], w7839, w7840);
  FullAdder U2516 (w7840, w7739, IN69[31], w7841, w7842);
  FullAdder U2517 (w7842, w7741, IN70[30], w7843, w7844);
  FullAdder U2518 (w7844, w7743, IN71[29], w7845, w7846);
  FullAdder U2519 (w7846, w7745, IN72[28], w7847, w7848);
  FullAdder U2520 (w7848, w7747, IN73[27], w7849, w7850);
  FullAdder U2521 (w7850, w7749, IN74[26], w7851, w7852);
  FullAdder U2522 (w7852, w7751, IN75[25], w7853, w7854);
  FullAdder U2523 (w7854, w7753, IN76[24], w7855, w7856);
  FullAdder U2524 (w7856, w7755, IN77[23], w7857, w7858);
  FullAdder U2525 (w7858, w7757, IN78[22], w7859, w7860);
  FullAdder U2526 (w7860, w7759, IN79[21], w7861, w7862);
  FullAdder U2527 (w7862, w7761, IN80[20], w7863, w7864);
  FullAdder U2528 (w7864, w7763, IN81[19], w7865, w7866);
  FullAdder U2529 (w7866, w7765, IN82[18], w7867, w7868);
  FullAdder U2530 (w7868, w7767, IN83[17], w7869, w7870);
  FullAdder U2531 (w7870, w7769, IN84[16], w7871, w7872);
  FullAdder U2532 (w7872, w7771, IN85[15], w7873, w7874);
  FullAdder U2533 (w7874, w7773, IN86[14], w7875, w7876);
  FullAdder U2534 (w7876, w7775, IN87[13], w7877, w7878);
  FullAdder U2535 (w7878, w7777, IN88[12], w7879, w7880);
  FullAdder U2536 (w7880, w7779, IN89[11], w7881, w7882);
  FullAdder U2537 (w7882, w7781, IN90[10], w7883, w7884);
  FullAdder U2538 (w7884, w7783, IN91[9], w7885, w7886);
  FullAdder U2539 (w7886, w7785, IN92[8], w7887, w7888);
  FullAdder U2540 (w7888, w7787, IN93[7], w7889, w7890);
  FullAdder U2541 (w7890, w7789, IN94[6], w7891, w7892);
  FullAdder U2542 (w7892, w7791, IN95[5], w7893, w7894);
  FullAdder U2543 (w7894, w7793, IN96[4], w7895, w7896);
  FullAdder U2544 (w7896, w7795, IN97[3], w7897, w7898);
  FullAdder U2545 (w7898, w7797, IN98[2], w7899, w7900);
  FullAdder U2546 (w7900, w7799, IN99[1], w7901, w7902);
  FullAdder U2547 (w7902, w7800, IN100[0], w7903, w7904);
  HalfAdder U2548 (w7803, IN50[50], Out1[50], w7906);
  FullAdder U2549 (w7906, w7805, IN51[50], w7907, w7908);
  FullAdder U2550 (w7908, w7807, IN52[50], w7909, w7910);
  FullAdder U2551 (w7910, w7809, IN53[48], w7911, w7912);
  FullAdder U2552 (w7912, w7811, IN54[47], w7913, w7914);
  FullAdder U2553 (w7914, w7813, IN55[46], w7915, w7916);
  FullAdder U2554 (w7916, w7815, IN56[45], w7917, w7918);
  FullAdder U2555 (w7918, w7817, IN57[44], w7919, w7920);
  FullAdder U2556 (w7920, w7819, IN58[43], w7921, w7922);
  FullAdder U2557 (w7922, w7821, IN59[42], w7923, w7924);
  FullAdder U2558 (w7924, w7823, IN60[41], w7925, w7926);
  FullAdder U2559 (w7926, w7825, IN61[40], w7927, w7928);
  FullAdder U2560 (w7928, w7827, IN62[39], w7929, w7930);
  FullAdder U2561 (w7930, w7829, IN63[38], w7931, w7932);
  FullAdder U2562 (w7932, w7831, IN64[37], w7933, w7934);
  FullAdder U2563 (w7934, w7833, IN65[36], w7935, w7936);
  FullAdder U2564 (w7936, w7835, IN66[35], w7937, w7938);
  FullAdder U2565 (w7938, w7837, IN67[34], w7939, w7940);
  FullAdder U2566 (w7940, w7839, IN68[33], w7941, w7942);
  FullAdder U2567 (w7942, w7841, IN69[32], w7943, w7944);
  FullAdder U2568 (w7944, w7843, IN70[31], w7945, w7946);
  FullAdder U2569 (w7946, w7845, IN71[30], w7947, w7948);
  FullAdder U2570 (w7948, w7847, IN72[29], w7949, w7950);
  FullAdder U2571 (w7950, w7849, IN73[28], w7951, w7952);
  FullAdder U2572 (w7952, w7851, IN74[27], w7953, w7954);
  FullAdder U2573 (w7954, w7853, IN75[26], w7955, w7956);
  FullAdder U2574 (w7956, w7855, IN76[25], w7957, w7958);
  FullAdder U2575 (w7958, w7857, IN77[24], w7959, w7960);
  FullAdder U2576 (w7960, w7859, IN78[23], w7961, w7962);
  FullAdder U2577 (w7962, w7861, IN79[22], w7963, w7964);
  FullAdder U2578 (w7964, w7863, IN80[21], w7965, w7966);
  FullAdder U2579 (w7966, w7865, IN81[20], w7967, w7968);
  FullAdder U2580 (w7968, w7867, IN82[19], w7969, w7970);
  FullAdder U2581 (w7970, w7869, IN83[18], w7971, w7972);
  FullAdder U2582 (w7972, w7871, IN84[17], w7973, w7974);
  FullAdder U2583 (w7974, w7873, IN85[16], w7975, w7976);
  FullAdder U2584 (w7976, w7875, IN86[15], w7977, w7978);
  FullAdder U2585 (w7978, w7877, IN87[14], w7979, w7980);
  FullAdder U2586 (w7980, w7879, IN88[13], w7981, w7982);
  FullAdder U2587 (w7982, w7881, IN89[12], w7983, w7984);
  FullAdder U2588 (w7984, w7883, IN90[11], w7985, w7986);
  FullAdder U2589 (w7986, w7885, IN91[10], w7987, w7988);
  FullAdder U2590 (w7988, w7887, IN92[9], w7989, w7990);
  FullAdder U2591 (w7990, w7889, IN93[8], w7991, w7992);
  FullAdder U2592 (w7992, w7891, IN94[7], w7993, w7994);
  FullAdder U2593 (w7994, w7893, IN95[6], w7995, w7996);
  FullAdder U2594 (w7996, w7895, IN96[5], w7997, w7998);
  FullAdder U2595 (w7998, w7897, IN97[4], w7999, w8000);
  FullAdder U2596 (w8000, w7899, IN98[3], w8001, w8002);
  FullAdder U2597 (w8002, w7901, IN99[2], w8003, w8004);
  FullAdder U2598 (w8004, w7903, IN100[1], w8005, w8006);
  FullAdder U2599 (w8006, w7904, IN101[0], w8007, w8008);
  HalfAdder U2600 (w7907, IN51[51], Out1[51], w8010);
  FullAdder U2601 (w8010, w7909, IN52[51], w8011, w8012);
  FullAdder U2602 (w8012, w7911, IN53[49], w8013, w8014);
  FullAdder U2603 (w8014, w7913, IN54[48], w8015, w8016);
  FullAdder U2604 (w8016, w7915, IN55[47], w8017, w8018);
  FullAdder U2605 (w8018, w7917, IN56[46], w8019, w8020);
  FullAdder U2606 (w8020, w7919, IN57[45], w8021, w8022);
  FullAdder U2607 (w8022, w7921, IN58[44], w8023, w8024);
  FullAdder U2608 (w8024, w7923, IN59[43], w8025, w8026);
  FullAdder U2609 (w8026, w7925, IN60[42], w8027, w8028);
  FullAdder U2610 (w8028, w7927, IN61[41], w8029, w8030);
  FullAdder U2611 (w8030, w7929, IN62[40], w8031, w8032);
  FullAdder U2612 (w8032, w7931, IN63[39], w8033, w8034);
  FullAdder U2613 (w8034, w7933, IN64[38], w8035, w8036);
  FullAdder U2614 (w8036, w7935, IN65[37], w8037, w8038);
  FullAdder U2615 (w8038, w7937, IN66[36], w8039, w8040);
  FullAdder U2616 (w8040, w7939, IN67[35], w8041, w8042);
  FullAdder U2617 (w8042, w7941, IN68[34], w8043, w8044);
  FullAdder U2618 (w8044, w7943, IN69[33], w8045, w8046);
  FullAdder U2619 (w8046, w7945, IN70[32], w8047, w8048);
  FullAdder U2620 (w8048, w7947, IN71[31], w8049, w8050);
  FullAdder U2621 (w8050, w7949, IN72[30], w8051, w8052);
  FullAdder U2622 (w8052, w7951, IN73[29], w8053, w8054);
  FullAdder U2623 (w8054, w7953, IN74[28], w8055, w8056);
  FullAdder U2624 (w8056, w7955, IN75[27], w8057, w8058);
  FullAdder U2625 (w8058, w7957, IN76[26], w8059, w8060);
  FullAdder U2626 (w8060, w7959, IN77[25], w8061, w8062);
  FullAdder U2627 (w8062, w7961, IN78[24], w8063, w8064);
  FullAdder U2628 (w8064, w7963, IN79[23], w8065, w8066);
  FullAdder U2629 (w8066, w7965, IN80[22], w8067, w8068);
  FullAdder U2630 (w8068, w7967, IN81[21], w8069, w8070);
  FullAdder U2631 (w8070, w7969, IN82[20], w8071, w8072);
  FullAdder U2632 (w8072, w7971, IN83[19], w8073, w8074);
  FullAdder U2633 (w8074, w7973, IN84[18], w8075, w8076);
  FullAdder U2634 (w8076, w7975, IN85[17], w8077, w8078);
  FullAdder U2635 (w8078, w7977, IN86[16], w8079, w8080);
  FullAdder U2636 (w8080, w7979, IN87[15], w8081, w8082);
  FullAdder U2637 (w8082, w7981, IN88[14], w8083, w8084);
  FullAdder U2638 (w8084, w7983, IN89[13], w8085, w8086);
  FullAdder U2639 (w8086, w7985, IN90[12], w8087, w8088);
  FullAdder U2640 (w8088, w7987, IN91[11], w8089, w8090);
  FullAdder U2641 (w8090, w7989, IN92[10], w8091, w8092);
  FullAdder U2642 (w8092, w7991, IN93[9], w8093, w8094);
  FullAdder U2643 (w8094, w7993, IN94[8], w8095, w8096);
  FullAdder U2644 (w8096, w7995, IN95[7], w8097, w8098);
  FullAdder U2645 (w8098, w7997, IN96[6], w8099, w8100);
  FullAdder U2646 (w8100, w7999, IN97[5], w8101, w8102);
  FullAdder U2647 (w8102, w8001, IN98[4], w8103, w8104);
  FullAdder U2648 (w8104, w8003, IN99[3], w8105, w8106);
  FullAdder U2649 (w8106, w8005, IN100[2], w8107, w8108);
  FullAdder U2650 (w8108, w8007, IN101[1], w8109, w8110);
  FullAdder U2651 (w8110, w8008, IN102[0], w8111, w8112);
  HalfAdder U2652 (w8011, IN52[52], Out1[52], w8114);
  FullAdder U2653 (w8114, w8013, IN53[50], Out1[53], w8116);
  FullAdder U2654 (w8116, w8015, IN54[49], Out1[54], w8118);
  FullAdder U2655 (w8118, w8017, IN55[48], Out1[55], w8120);
  FullAdder U2656 (w8120, w8019, IN56[47], Out1[56], w8122);
  FullAdder U2657 (w8122, w8021, IN57[46], Out1[57], w8124);
  FullAdder U2658 (w8124, w8023, IN58[45], Out1[58], w8126);
  FullAdder U2659 (w8126, w8025, IN59[44], Out1[59], w8128);
  FullAdder U2660 (w8128, w8027, IN60[43], Out1[60], w8130);
  FullAdder U2661 (w8130, w8029, IN61[42], Out1[61], w8132);
  FullAdder U2662 (w8132, w8031, IN62[41], Out1[62], w8134);
  FullAdder U2663 (w8134, w8033, IN63[40], Out1[63], w8136);
  FullAdder U2664 (w8136, w8035, IN64[39], Out1[64], w8138);
  FullAdder U2665 (w8138, w8037, IN65[38], Out1[65], w8140);
  FullAdder U2666 (w8140, w8039, IN66[37], Out1[66], w8142);
  FullAdder U2667 (w8142, w8041, IN67[36], Out1[67], w8144);
  FullAdder U2668 (w8144, w8043, IN68[35], Out1[68], w8146);
  FullAdder U2669 (w8146, w8045, IN69[34], Out1[69], w8148);
  FullAdder U2670 (w8148, w8047, IN70[33], Out1[70], w8150);
  FullAdder U2671 (w8150, w8049, IN71[32], Out1[71], w8152);
  FullAdder U2672 (w8152, w8051, IN72[31], Out1[72], w8154);
  FullAdder U2673 (w8154, w8053, IN73[30], Out1[73], w8156);
  FullAdder U2674 (w8156, w8055, IN74[29], Out1[74], w8158);
  FullAdder U2675 (w8158, w8057, IN75[28], Out1[75], w8160);
  FullAdder U2676 (w8160, w8059, IN76[27], Out1[76], w8162);
  FullAdder U2677 (w8162, w8061, IN77[26], Out1[77], w8164);
  FullAdder U2678 (w8164, w8063, IN78[25], Out1[78], w8166);
  FullAdder U2679 (w8166, w8065, IN79[24], Out1[79], w8168);
  FullAdder U2680 (w8168, w8067, IN80[23], Out1[80], w8170);
  FullAdder U2681 (w8170, w8069, IN81[22], Out1[81], w8172);
  FullAdder U2682 (w8172, w8071, IN82[21], Out1[82], w8174);
  FullAdder U2683 (w8174, w8073, IN83[20], Out1[83], w8176);
  FullAdder U2684 (w8176, w8075, IN84[19], Out1[84], w8178);
  FullAdder U2685 (w8178, w8077, IN85[18], Out1[85], w8180);
  FullAdder U2686 (w8180, w8079, IN86[17], Out1[86], w8182);
  FullAdder U2687 (w8182, w8081, IN87[16], Out1[87], w8184);
  FullAdder U2688 (w8184, w8083, IN88[15], Out1[88], w8186);
  FullAdder U2689 (w8186, w8085, IN89[14], Out1[89], w8188);
  FullAdder U2690 (w8188, w8087, IN90[13], Out1[90], w8190);
  FullAdder U2691 (w8190, w8089, IN91[12], Out1[91], w8192);
  FullAdder U2692 (w8192, w8091, IN92[11], Out1[92], w8194);
  FullAdder U2693 (w8194, w8093, IN93[10], Out1[93], w8196);
  FullAdder U2694 (w8196, w8095, IN94[9], Out1[94], w8198);
  FullAdder U2695 (w8198, w8097, IN95[8], Out1[95], w8200);
  FullAdder U2696 (w8200, w8099, IN96[7], Out1[96], w8202);
  FullAdder U2697 (w8202, w8101, IN97[6], Out1[97], w8204);
  FullAdder U2698 (w8204, w8103, IN98[5], Out1[98], w8206);
  FullAdder U2699 (w8206, w8105, IN99[4], Out1[99], w8208);
  FullAdder U2700 (w8208, w8107, IN100[3], Out1[100], w8210);
  FullAdder U2701 (w8210, w8109, IN101[2], Out1[101], w8212);
  FullAdder U2702 (w8212, w8111, IN102[1], Out1[102], w8214);
  FullAdder U2703 (w8214, w8112, IN103[0], Out1[103], Out1[104]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN53[51];
  assign Out2[1] = IN54[50];
  assign Out2[2] = IN55[49];
  assign Out2[3] = IN56[48];
  assign Out2[4] = IN57[47];
  assign Out2[5] = IN58[46];
  assign Out2[6] = IN59[45];
  assign Out2[7] = IN60[44];
  assign Out2[8] = IN61[43];
  assign Out2[9] = IN62[42];
  assign Out2[10] = IN63[41];
  assign Out2[11] = IN64[40];
  assign Out2[12] = IN65[39];
  assign Out2[13] = IN66[38];
  assign Out2[14] = IN67[37];
  assign Out2[15] = IN68[36];
  assign Out2[16] = IN69[35];
  assign Out2[17] = IN70[34];
  assign Out2[18] = IN71[33];
  assign Out2[19] = IN72[32];
  assign Out2[20] = IN73[31];
  assign Out2[21] = IN74[30];
  assign Out2[22] = IN75[29];
  assign Out2[23] = IN76[28];
  assign Out2[24] = IN77[27];
  assign Out2[25] = IN78[26];
  assign Out2[26] = IN79[25];
  assign Out2[27] = IN80[24];
  assign Out2[28] = IN81[23];
  assign Out2[29] = IN82[22];
  assign Out2[30] = IN83[21];
  assign Out2[31] = IN84[20];
  assign Out2[32] = IN85[19];
  assign Out2[33] = IN86[18];
  assign Out2[34] = IN87[17];
  assign Out2[35] = IN88[16];
  assign Out2[36] = IN89[15];
  assign Out2[37] = IN90[14];
  assign Out2[38] = IN91[13];
  assign Out2[39] = IN92[12];
  assign Out2[40] = IN93[11];
  assign Out2[41] = IN94[10];
  assign Out2[42] = IN95[9];
  assign Out2[43] = IN96[8];
  assign Out2[44] = IN97[7];
  assign Out2[45] = IN98[6];
  assign Out2[46] = IN99[5];
  assign Out2[47] = IN100[4];
  assign Out2[48] = IN101[3];
  assign Out2[49] = IN102[2];
  assign Out2[50] = IN103[1];
  assign Out2[51] = IN104[0];

endmodule
module RC_52_52(IN1, IN2, Out);
  input [51:0] IN1;
  input [51:0] IN2;
  output [52:0] Out;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w105);
  FullAdder U1 (IN1[1], IN2[1], w105, Out[1], w107);
  FullAdder U2 (IN1[2], IN2[2], w107, Out[2], w109);
  FullAdder U3 (IN1[3], IN2[3], w109, Out[3], w111);
  FullAdder U4 (IN1[4], IN2[4], w111, Out[4], w113);
  FullAdder U5 (IN1[5], IN2[5], w113, Out[5], w115);
  FullAdder U6 (IN1[6], IN2[6], w115, Out[6], w117);
  FullAdder U7 (IN1[7], IN2[7], w117, Out[7], w119);
  FullAdder U8 (IN1[8], IN2[8], w119, Out[8], w121);
  FullAdder U9 (IN1[9], IN2[9], w121, Out[9], w123);
  FullAdder U10 (IN1[10], IN2[10], w123, Out[10], w125);
  FullAdder U11 (IN1[11], IN2[11], w125, Out[11], w127);
  FullAdder U12 (IN1[12], IN2[12], w127, Out[12], w129);
  FullAdder U13 (IN1[13], IN2[13], w129, Out[13], w131);
  FullAdder U14 (IN1[14], IN2[14], w131, Out[14], w133);
  FullAdder U15 (IN1[15], IN2[15], w133, Out[15], w135);
  FullAdder U16 (IN1[16], IN2[16], w135, Out[16], w137);
  FullAdder U17 (IN1[17], IN2[17], w137, Out[17], w139);
  FullAdder U18 (IN1[18], IN2[18], w139, Out[18], w141);
  FullAdder U19 (IN1[19], IN2[19], w141, Out[19], w143);
  FullAdder U20 (IN1[20], IN2[20], w143, Out[20], w145);
  FullAdder U21 (IN1[21], IN2[21], w145, Out[21], w147);
  FullAdder U22 (IN1[22], IN2[22], w147, Out[22], w149);
  FullAdder U23 (IN1[23], IN2[23], w149, Out[23], w151);
  FullAdder U24 (IN1[24], IN2[24], w151, Out[24], w153);
  FullAdder U25 (IN1[25], IN2[25], w153, Out[25], w155);
  FullAdder U26 (IN1[26], IN2[26], w155, Out[26], w157);
  FullAdder U27 (IN1[27], IN2[27], w157, Out[27], w159);
  FullAdder U28 (IN1[28], IN2[28], w159, Out[28], w161);
  FullAdder U29 (IN1[29], IN2[29], w161, Out[29], w163);
  FullAdder U30 (IN1[30], IN2[30], w163, Out[30], w165);
  FullAdder U31 (IN1[31], IN2[31], w165, Out[31], w167);
  FullAdder U32 (IN1[32], IN2[32], w167, Out[32], w169);
  FullAdder U33 (IN1[33], IN2[33], w169, Out[33], w171);
  FullAdder U34 (IN1[34], IN2[34], w171, Out[34], w173);
  FullAdder U35 (IN1[35], IN2[35], w173, Out[35], w175);
  FullAdder U36 (IN1[36], IN2[36], w175, Out[36], w177);
  FullAdder U37 (IN1[37], IN2[37], w177, Out[37], w179);
  FullAdder U38 (IN1[38], IN2[38], w179, Out[38], w181);
  FullAdder U39 (IN1[39], IN2[39], w181, Out[39], w183);
  FullAdder U40 (IN1[40], IN2[40], w183, Out[40], w185);
  FullAdder U41 (IN1[41], IN2[41], w185, Out[41], w187);
  FullAdder U42 (IN1[42], IN2[42], w187, Out[42], w189);
  FullAdder U43 (IN1[43], IN2[43], w189, Out[43], w191);
  FullAdder U44 (IN1[44], IN2[44], w191, Out[44], w193);
  FullAdder U45 (IN1[45], IN2[45], w193, Out[45], w195);
  FullAdder U46 (IN1[46], IN2[46], w195, Out[46], w197);
  FullAdder U47 (IN1[47], IN2[47], w197, Out[47], w199);
  FullAdder U48 (IN1[48], IN2[48], w199, Out[48], w201);
  FullAdder U49 (IN1[49], IN2[49], w201, Out[49], w203);
  FullAdder U50 (IN1[50], IN2[50], w203, Out[50], w205);
  FullAdder U51 (IN1[51], IN2[51], w205, Out[51], Out[52]);

endmodule
module NR_53_53(IN1, IN2, Out);
  input [52:0] IN1;
  input [52:0] IN2;
  output [105:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [29:0] P29;
  wire [30:0] P30;
  wire [31:0] P31;
  wire [32:0] P32;
  wire [33:0] P33;
  wire [34:0] P34;
  wire [35:0] P35;
  wire [36:0] P36;
  wire [37:0] P37;
  wire [38:0] P38;
  wire [39:0] P39;
  wire [40:0] P40;
  wire [41:0] P41;
  wire [42:0] P42;
  wire [43:0] P43;
  wire [44:0] P44;
  wire [45:0] P45;
  wire [46:0] P46;
  wire [47:0] P47;
  wire [48:0] P48;
  wire [49:0] P49;
  wire [50:0] P50;
  wire [51:0] P51;
  wire [52:0] P52;
  wire [51:0] P53;
  wire [50:0] P54;
  wire [49:0] P55;
  wire [48:0] P56;
  wire [47:0] P57;
  wire [46:0] P58;
  wire [45:0] P59;
  wire [44:0] P60;
  wire [43:0] P61;
  wire [42:0] P62;
  wire [41:0] P63;
  wire [40:0] P64;
  wire [39:0] P65;
  wire [38:0] P66;
  wire [37:0] P67;
  wire [36:0] P68;
  wire [35:0] P69;
  wire [34:0] P70;
  wire [33:0] P71;
  wire [32:0] P72;
  wire [31:0] P73;
  wire [30:0] P74;
  wire [29:0] P75;
  wire [28:0] P76;
  wire [27:0] P77;
  wire [26:0] P78;
  wire [25:0] P79;
  wire [24:0] P80;
  wire [23:0] P81;
  wire [22:0] P82;
  wire [21:0] P83;
  wire [20:0] P84;
  wire [19:0] P85;
  wire [18:0] P86;
  wire [17:0] P87;
  wire [16:0] P88;
  wire [15:0] P89;
  wire [14:0] P90;
  wire [13:0] P91;
  wire [12:0] P92;
  wire [11:0] P93;
  wire [10:0] P94;
  wire [9:0] P95;
  wire [8:0] P96;
  wire [7:0] P97;
  wire [6:0] P98;
  wire [5:0] P99;
  wire [4:0] P100;
  wire [3:0] P101;
  wire [2:0] P102;
  wire [1:0] P103;
  wire [0:0] P104;
  wire [104:0] R1;
  wire [51:0] R2;
  wire [105:0] aOut;
  U_SP_53_53 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, R1, R2);
  RC_52_52 S2 (R1[104:53], R2, aOut[105:53]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign Out = aOut[105:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
