
module NR_58_1(
    input [57:0]IN1,
    input [0:0]IN2,
    output [57:0]Out
);
    assign Out = IN2;
endmodule
