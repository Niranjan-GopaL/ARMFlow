//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 12
  second input length: 36
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_12_36(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46);
  input [11:0] IN1;
  input [35:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [11:0] P12;
  output [11:0] P13;
  output [11:0] P14;
  output [11:0] P15;
  output [11:0] P16;
  output [11:0] P17;
  output [11:0] P18;
  output [11:0] P19;
  output [11:0] P20;
  output [11:0] P21;
  output [11:0] P22;
  output [11:0] P23;
  output [11:0] P24;
  output [11:0] P25;
  output [11:0] P26;
  output [11:0] P27;
  output [11:0] P28;
  output [11:0] P29;
  output [11:0] P30;
  output [11:0] P31;
  output [11:0] P32;
  output [11:0] P33;
  output [11:0] P34;
  output [11:0] P35;
  output [10:0] P36;
  output [9:0] P37;
  output [8:0] P38;
  output [7:0] P39;
  output [6:0] P40;
  output [5:0] P41;
  output [4:0] P42;
  output [3:0] P43;
  output [2:0] P44;
  output [1:0] P45;
  output [0:0] P46;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[0] = IN1[1]&IN2[35];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[1] = IN1[2]&IN2[34];
  assign P37[0] = IN1[2]&IN2[35];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[2] = IN1[3]&IN2[33];
  assign P37[1] = IN1[3]&IN2[34];
  assign P38[0] = IN1[3]&IN2[35];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[3] = IN1[4]&IN2[32];
  assign P37[2] = IN1[4]&IN2[33];
  assign P38[1] = IN1[4]&IN2[34];
  assign P39[0] = IN1[4]&IN2[35];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[4] = IN1[5]&IN2[31];
  assign P37[3] = IN1[5]&IN2[32];
  assign P38[2] = IN1[5]&IN2[33];
  assign P39[1] = IN1[5]&IN2[34];
  assign P40[0] = IN1[5]&IN2[35];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[5] = IN1[6]&IN2[30];
  assign P37[4] = IN1[6]&IN2[31];
  assign P38[3] = IN1[6]&IN2[32];
  assign P39[2] = IN1[6]&IN2[33];
  assign P40[1] = IN1[6]&IN2[34];
  assign P41[0] = IN1[6]&IN2[35];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[6] = IN1[7]&IN2[29];
  assign P37[5] = IN1[7]&IN2[30];
  assign P38[4] = IN1[7]&IN2[31];
  assign P39[3] = IN1[7]&IN2[32];
  assign P40[2] = IN1[7]&IN2[33];
  assign P41[1] = IN1[7]&IN2[34];
  assign P42[0] = IN1[7]&IN2[35];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[7] = IN1[8]&IN2[28];
  assign P37[6] = IN1[8]&IN2[29];
  assign P38[5] = IN1[8]&IN2[30];
  assign P39[4] = IN1[8]&IN2[31];
  assign P40[3] = IN1[8]&IN2[32];
  assign P41[2] = IN1[8]&IN2[33];
  assign P42[1] = IN1[8]&IN2[34];
  assign P43[0] = IN1[8]&IN2[35];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[8] = IN1[9]&IN2[27];
  assign P37[7] = IN1[9]&IN2[28];
  assign P38[6] = IN1[9]&IN2[29];
  assign P39[5] = IN1[9]&IN2[30];
  assign P40[4] = IN1[9]&IN2[31];
  assign P41[3] = IN1[9]&IN2[32];
  assign P42[2] = IN1[9]&IN2[33];
  assign P43[1] = IN1[9]&IN2[34];
  assign P44[0] = IN1[9]&IN2[35];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[9] = IN1[10]&IN2[26];
  assign P37[8] = IN1[10]&IN2[27];
  assign P38[7] = IN1[10]&IN2[28];
  assign P39[6] = IN1[10]&IN2[29];
  assign P40[5] = IN1[10]&IN2[30];
  assign P41[4] = IN1[10]&IN2[31];
  assign P42[3] = IN1[10]&IN2[32];
  assign P43[2] = IN1[10]&IN2[33];
  assign P44[1] = IN1[10]&IN2[34];
  assign P45[0] = IN1[10]&IN2[35];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[10] = IN1[11]&IN2[25];
  assign P37[9] = IN1[11]&IN2[26];
  assign P38[8] = IN1[11]&IN2[27];
  assign P39[7] = IN1[11]&IN2[28];
  assign P40[6] = IN1[11]&IN2[29];
  assign P41[5] = IN1[11]&IN2[30];
  assign P42[4] = IN1[11]&IN2[31];
  assign P43[3] = IN1[11]&IN2[32];
  assign P44[2] = IN1[11]&IN2[33];
  assign P45[1] = IN1[11]&IN2[34];
  assign P46[0] = IN1[11]&IN2[35];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [11:0] IN12;
  input [11:0] IN13;
  input [11:0] IN14;
  input [11:0] IN15;
  input [11:0] IN16;
  input [11:0] IN17;
  input [11:0] IN18;
  input [11:0] IN19;
  input [11:0] IN20;
  input [11:0] IN21;
  input [11:0] IN22;
  input [11:0] IN23;
  input [11:0] IN24;
  input [11:0] IN25;
  input [11:0] IN26;
  input [11:0] IN27;
  input [11:0] IN28;
  input [11:0] IN29;
  input [11:0] IN30;
  input [11:0] IN31;
  input [11:0] IN32;
  input [11:0] IN33;
  input [11:0] IN34;
  input [11:0] IN35;
  input [10:0] IN36;
  input [9:0] IN37;
  input [8:0] IN38;
  input [7:0] IN39;
  input [6:0] IN40;
  input [5:0] IN41;
  input [4:0] IN42;
  input [3:0] IN43;
  input [2:0] IN44;
  input [1:0] IN45;
  input [0:0] IN46;
  output [46:0] Out1;
  output [34:0] Out2;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1181;
  wire w1183;
  wire w1185;
  wire w1187;
  wire w1189;
  wire w1191;
  wire w1193;
  wire w1195;
  wire w1197;
  wire w1199;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w433);
  FullAdder U1 (w433, IN2[0], IN2[1], w434, w435);
  FullAdder U2 (w435, IN3[0], IN3[1], w436, w437);
  FullAdder U3 (w437, IN4[0], IN4[1], w438, w439);
  FullAdder U4 (w439, IN5[0], IN5[1], w440, w441);
  FullAdder U5 (w441, IN6[0], IN6[1], w442, w443);
  FullAdder U6 (w443, IN7[0], IN7[1], w444, w445);
  FullAdder U7 (w445, IN8[0], IN8[1], w446, w447);
  FullAdder U8 (w447, IN9[0], IN9[1], w448, w449);
  FullAdder U9 (w449, IN10[0], IN10[1], w450, w451);
  FullAdder U10 (w451, IN11[0], IN11[1], w452, w453);
  HalfAdder U11 (w434, IN2[2], Out1[2], w455);
  FullAdder U12 (w455, w436, IN3[2], w456, w457);
  FullAdder U13 (w457, w438, IN4[2], w458, w459);
  FullAdder U14 (w459, w440, IN5[2], w460, w461);
  FullAdder U15 (w461, w442, IN6[2], w462, w463);
  FullAdder U16 (w463, w444, IN7[2], w464, w465);
  FullAdder U17 (w465, w446, IN8[2], w466, w467);
  FullAdder U18 (w467, w448, IN9[2], w468, w469);
  FullAdder U19 (w469, w450, IN10[2], w470, w471);
  FullAdder U20 (w471, w452, IN11[2], w472, w473);
  FullAdder U21 (w473, w453, IN12[0], w474, w475);
  HalfAdder U22 (w456, IN3[3], Out1[3], w477);
  FullAdder U23 (w477, w458, IN4[3], w478, w479);
  FullAdder U24 (w479, w460, IN5[3], w480, w481);
  FullAdder U25 (w481, w462, IN6[3], w482, w483);
  FullAdder U26 (w483, w464, IN7[3], w484, w485);
  FullAdder U27 (w485, w466, IN8[3], w486, w487);
  FullAdder U28 (w487, w468, IN9[3], w488, w489);
  FullAdder U29 (w489, w470, IN10[3], w490, w491);
  FullAdder U30 (w491, w472, IN11[3], w492, w493);
  FullAdder U31 (w493, w474, IN12[1], w494, w495);
  FullAdder U32 (w495, w475, IN13[0], w496, w497);
  HalfAdder U33 (w478, IN4[4], Out1[4], w499);
  FullAdder U34 (w499, w480, IN5[4], w500, w501);
  FullAdder U35 (w501, w482, IN6[4], w502, w503);
  FullAdder U36 (w503, w484, IN7[4], w504, w505);
  FullAdder U37 (w505, w486, IN8[4], w506, w507);
  FullAdder U38 (w507, w488, IN9[4], w508, w509);
  FullAdder U39 (w509, w490, IN10[4], w510, w511);
  FullAdder U40 (w511, w492, IN11[4], w512, w513);
  FullAdder U41 (w513, w494, IN12[2], w514, w515);
  FullAdder U42 (w515, w496, IN13[1], w516, w517);
  FullAdder U43 (w517, w497, IN14[0], w518, w519);
  HalfAdder U44 (w500, IN5[5], Out1[5], w521);
  FullAdder U45 (w521, w502, IN6[5], w522, w523);
  FullAdder U46 (w523, w504, IN7[5], w524, w525);
  FullAdder U47 (w525, w506, IN8[5], w526, w527);
  FullAdder U48 (w527, w508, IN9[5], w528, w529);
  FullAdder U49 (w529, w510, IN10[5], w530, w531);
  FullAdder U50 (w531, w512, IN11[5], w532, w533);
  FullAdder U51 (w533, w514, IN12[3], w534, w535);
  FullAdder U52 (w535, w516, IN13[2], w536, w537);
  FullAdder U53 (w537, w518, IN14[1], w538, w539);
  FullAdder U54 (w539, w519, IN15[0], w540, w541);
  HalfAdder U55 (w522, IN6[6], Out1[6], w543);
  FullAdder U56 (w543, w524, IN7[6], w544, w545);
  FullAdder U57 (w545, w526, IN8[6], w546, w547);
  FullAdder U58 (w547, w528, IN9[6], w548, w549);
  FullAdder U59 (w549, w530, IN10[6], w550, w551);
  FullAdder U60 (w551, w532, IN11[6], w552, w553);
  FullAdder U61 (w553, w534, IN12[4], w554, w555);
  FullAdder U62 (w555, w536, IN13[3], w556, w557);
  FullAdder U63 (w557, w538, IN14[2], w558, w559);
  FullAdder U64 (w559, w540, IN15[1], w560, w561);
  FullAdder U65 (w561, w541, IN16[0], w562, w563);
  HalfAdder U66 (w544, IN7[7], Out1[7], w565);
  FullAdder U67 (w565, w546, IN8[7], w566, w567);
  FullAdder U68 (w567, w548, IN9[7], w568, w569);
  FullAdder U69 (w569, w550, IN10[7], w570, w571);
  FullAdder U70 (w571, w552, IN11[7], w572, w573);
  FullAdder U71 (w573, w554, IN12[5], w574, w575);
  FullAdder U72 (w575, w556, IN13[4], w576, w577);
  FullAdder U73 (w577, w558, IN14[3], w578, w579);
  FullAdder U74 (w579, w560, IN15[2], w580, w581);
  FullAdder U75 (w581, w562, IN16[1], w582, w583);
  FullAdder U76 (w583, w563, IN17[0], w584, w585);
  HalfAdder U77 (w566, IN8[8], Out1[8], w587);
  FullAdder U78 (w587, w568, IN9[8], w588, w589);
  FullAdder U79 (w589, w570, IN10[8], w590, w591);
  FullAdder U80 (w591, w572, IN11[8], w592, w593);
  FullAdder U81 (w593, w574, IN12[6], w594, w595);
  FullAdder U82 (w595, w576, IN13[5], w596, w597);
  FullAdder U83 (w597, w578, IN14[4], w598, w599);
  FullAdder U84 (w599, w580, IN15[3], w600, w601);
  FullAdder U85 (w601, w582, IN16[2], w602, w603);
  FullAdder U86 (w603, w584, IN17[1], w604, w605);
  FullAdder U87 (w605, w585, IN18[0], w606, w607);
  HalfAdder U88 (w588, IN9[9], Out1[9], w609);
  FullAdder U89 (w609, w590, IN10[9], w610, w611);
  FullAdder U90 (w611, w592, IN11[9], w612, w613);
  FullAdder U91 (w613, w594, IN12[7], w614, w615);
  FullAdder U92 (w615, w596, IN13[6], w616, w617);
  FullAdder U93 (w617, w598, IN14[5], w618, w619);
  FullAdder U94 (w619, w600, IN15[4], w620, w621);
  FullAdder U95 (w621, w602, IN16[3], w622, w623);
  FullAdder U96 (w623, w604, IN17[2], w624, w625);
  FullAdder U97 (w625, w606, IN18[1], w626, w627);
  FullAdder U98 (w627, w607, IN19[0], w628, w629);
  HalfAdder U99 (w610, IN10[10], Out1[10], w631);
  FullAdder U100 (w631, w612, IN11[10], w632, w633);
  FullAdder U101 (w633, w614, IN12[8], w634, w635);
  FullAdder U102 (w635, w616, IN13[7], w636, w637);
  FullAdder U103 (w637, w618, IN14[6], w638, w639);
  FullAdder U104 (w639, w620, IN15[5], w640, w641);
  FullAdder U105 (w641, w622, IN16[4], w642, w643);
  FullAdder U106 (w643, w624, IN17[3], w644, w645);
  FullAdder U107 (w645, w626, IN18[2], w646, w647);
  FullAdder U108 (w647, w628, IN19[1], w648, w649);
  FullAdder U109 (w649, w629, IN20[0], w650, w651);
  HalfAdder U110 (w632, IN11[11], Out1[11], w653);
  FullAdder U111 (w653, w634, IN12[9], w654, w655);
  FullAdder U112 (w655, w636, IN13[8], w656, w657);
  FullAdder U113 (w657, w638, IN14[7], w658, w659);
  FullAdder U114 (w659, w640, IN15[6], w660, w661);
  FullAdder U115 (w661, w642, IN16[5], w662, w663);
  FullAdder U116 (w663, w644, IN17[4], w664, w665);
  FullAdder U117 (w665, w646, IN18[3], w666, w667);
  FullAdder U118 (w667, w648, IN19[2], w668, w669);
  FullAdder U119 (w669, w650, IN20[1], w670, w671);
  FullAdder U120 (w671, w651, IN21[0], w672, w673);
  HalfAdder U121 (w654, IN12[10], Out1[12], w675);
  FullAdder U122 (w675, w656, IN13[9], w676, w677);
  FullAdder U123 (w677, w658, IN14[8], w678, w679);
  FullAdder U124 (w679, w660, IN15[7], w680, w681);
  FullAdder U125 (w681, w662, IN16[6], w682, w683);
  FullAdder U126 (w683, w664, IN17[5], w684, w685);
  FullAdder U127 (w685, w666, IN18[4], w686, w687);
  FullAdder U128 (w687, w668, IN19[3], w688, w689);
  FullAdder U129 (w689, w670, IN20[2], w690, w691);
  FullAdder U130 (w691, w672, IN21[1], w692, w693);
  FullAdder U131 (w693, w673, IN22[0], w694, w695);
  HalfAdder U132 (w676, IN13[10], Out1[13], w697);
  FullAdder U133 (w697, w678, IN14[9], w698, w699);
  FullAdder U134 (w699, w680, IN15[8], w700, w701);
  FullAdder U135 (w701, w682, IN16[7], w702, w703);
  FullAdder U136 (w703, w684, IN17[6], w704, w705);
  FullAdder U137 (w705, w686, IN18[5], w706, w707);
  FullAdder U138 (w707, w688, IN19[4], w708, w709);
  FullAdder U139 (w709, w690, IN20[3], w710, w711);
  FullAdder U140 (w711, w692, IN21[2], w712, w713);
  FullAdder U141 (w713, w694, IN22[1], w714, w715);
  FullAdder U142 (w715, w695, IN23[0], w716, w717);
  HalfAdder U143 (w698, IN14[10], Out1[14], w719);
  FullAdder U144 (w719, w700, IN15[9], w720, w721);
  FullAdder U145 (w721, w702, IN16[8], w722, w723);
  FullAdder U146 (w723, w704, IN17[7], w724, w725);
  FullAdder U147 (w725, w706, IN18[6], w726, w727);
  FullAdder U148 (w727, w708, IN19[5], w728, w729);
  FullAdder U149 (w729, w710, IN20[4], w730, w731);
  FullAdder U150 (w731, w712, IN21[3], w732, w733);
  FullAdder U151 (w733, w714, IN22[2], w734, w735);
  FullAdder U152 (w735, w716, IN23[1], w736, w737);
  FullAdder U153 (w737, w717, IN24[0], w738, w739);
  HalfAdder U154 (w720, IN15[10], Out1[15], w741);
  FullAdder U155 (w741, w722, IN16[9], w742, w743);
  FullAdder U156 (w743, w724, IN17[8], w744, w745);
  FullAdder U157 (w745, w726, IN18[7], w746, w747);
  FullAdder U158 (w747, w728, IN19[6], w748, w749);
  FullAdder U159 (w749, w730, IN20[5], w750, w751);
  FullAdder U160 (w751, w732, IN21[4], w752, w753);
  FullAdder U161 (w753, w734, IN22[3], w754, w755);
  FullAdder U162 (w755, w736, IN23[2], w756, w757);
  FullAdder U163 (w757, w738, IN24[1], w758, w759);
  FullAdder U164 (w759, w739, IN25[0], w760, w761);
  HalfAdder U165 (w742, IN16[10], Out1[16], w763);
  FullAdder U166 (w763, w744, IN17[9], w764, w765);
  FullAdder U167 (w765, w746, IN18[8], w766, w767);
  FullAdder U168 (w767, w748, IN19[7], w768, w769);
  FullAdder U169 (w769, w750, IN20[6], w770, w771);
  FullAdder U170 (w771, w752, IN21[5], w772, w773);
  FullAdder U171 (w773, w754, IN22[4], w774, w775);
  FullAdder U172 (w775, w756, IN23[3], w776, w777);
  FullAdder U173 (w777, w758, IN24[2], w778, w779);
  FullAdder U174 (w779, w760, IN25[1], w780, w781);
  FullAdder U175 (w781, w761, IN26[0], w782, w783);
  HalfAdder U176 (w764, IN17[10], Out1[17], w785);
  FullAdder U177 (w785, w766, IN18[9], w786, w787);
  FullAdder U178 (w787, w768, IN19[8], w788, w789);
  FullAdder U179 (w789, w770, IN20[7], w790, w791);
  FullAdder U180 (w791, w772, IN21[6], w792, w793);
  FullAdder U181 (w793, w774, IN22[5], w794, w795);
  FullAdder U182 (w795, w776, IN23[4], w796, w797);
  FullAdder U183 (w797, w778, IN24[3], w798, w799);
  FullAdder U184 (w799, w780, IN25[2], w800, w801);
  FullAdder U185 (w801, w782, IN26[1], w802, w803);
  FullAdder U186 (w803, w783, IN27[0], w804, w805);
  HalfAdder U187 (w786, IN18[10], Out1[18], w807);
  FullAdder U188 (w807, w788, IN19[9], w808, w809);
  FullAdder U189 (w809, w790, IN20[8], w810, w811);
  FullAdder U190 (w811, w792, IN21[7], w812, w813);
  FullAdder U191 (w813, w794, IN22[6], w814, w815);
  FullAdder U192 (w815, w796, IN23[5], w816, w817);
  FullAdder U193 (w817, w798, IN24[4], w818, w819);
  FullAdder U194 (w819, w800, IN25[3], w820, w821);
  FullAdder U195 (w821, w802, IN26[2], w822, w823);
  FullAdder U196 (w823, w804, IN27[1], w824, w825);
  FullAdder U197 (w825, w805, IN28[0], w826, w827);
  HalfAdder U198 (w808, IN19[10], Out1[19], w829);
  FullAdder U199 (w829, w810, IN20[9], w830, w831);
  FullAdder U200 (w831, w812, IN21[8], w832, w833);
  FullAdder U201 (w833, w814, IN22[7], w834, w835);
  FullAdder U202 (w835, w816, IN23[6], w836, w837);
  FullAdder U203 (w837, w818, IN24[5], w838, w839);
  FullAdder U204 (w839, w820, IN25[4], w840, w841);
  FullAdder U205 (w841, w822, IN26[3], w842, w843);
  FullAdder U206 (w843, w824, IN27[2], w844, w845);
  FullAdder U207 (w845, w826, IN28[1], w846, w847);
  FullAdder U208 (w847, w827, IN29[0], w848, w849);
  HalfAdder U209 (w830, IN20[10], Out1[20], w851);
  FullAdder U210 (w851, w832, IN21[9], w852, w853);
  FullAdder U211 (w853, w834, IN22[8], w854, w855);
  FullAdder U212 (w855, w836, IN23[7], w856, w857);
  FullAdder U213 (w857, w838, IN24[6], w858, w859);
  FullAdder U214 (w859, w840, IN25[5], w860, w861);
  FullAdder U215 (w861, w842, IN26[4], w862, w863);
  FullAdder U216 (w863, w844, IN27[3], w864, w865);
  FullAdder U217 (w865, w846, IN28[2], w866, w867);
  FullAdder U218 (w867, w848, IN29[1], w868, w869);
  FullAdder U219 (w869, w849, IN30[0], w870, w871);
  HalfAdder U220 (w852, IN21[10], Out1[21], w873);
  FullAdder U221 (w873, w854, IN22[9], w874, w875);
  FullAdder U222 (w875, w856, IN23[8], w876, w877);
  FullAdder U223 (w877, w858, IN24[7], w878, w879);
  FullAdder U224 (w879, w860, IN25[6], w880, w881);
  FullAdder U225 (w881, w862, IN26[5], w882, w883);
  FullAdder U226 (w883, w864, IN27[4], w884, w885);
  FullAdder U227 (w885, w866, IN28[3], w886, w887);
  FullAdder U228 (w887, w868, IN29[2], w888, w889);
  FullAdder U229 (w889, w870, IN30[1], w890, w891);
  FullAdder U230 (w891, w871, IN31[0], w892, w893);
  HalfAdder U231 (w874, IN22[10], Out1[22], w895);
  FullAdder U232 (w895, w876, IN23[9], w896, w897);
  FullAdder U233 (w897, w878, IN24[8], w898, w899);
  FullAdder U234 (w899, w880, IN25[7], w900, w901);
  FullAdder U235 (w901, w882, IN26[6], w902, w903);
  FullAdder U236 (w903, w884, IN27[5], w904, w905);
  FullAdder U237 (w905, w886, IN28[4], w906, w907);
  FullAdder U238 (w907, w888, IN29[3], w908, w909);
  FullAdder U239 (w909, w890, IN30[2], w910, w911);
  FullAdder U240 (w911, w892, IN31[1], w912, w913);
  FullAdder U241 (w913, w893, IN32[0], w914, w915);
  HalfAdder U242 (w896, IN23[10], Out1[23], w917);
  FullAdder U243 (w917, w898, IN24[9], w918, w919);
  FullAdder U244 (w919, w900, IN25[8], w920, w921);
  FullAdder U245 (w921, w902, IN26[7], w922, w923);
  FullAdder U246 (w923, w904, IN27[6], w924, w925);
  FullAdder U247 (w925, w906, IN28[5], w926, w927);
  FullAdder U248 (w927, w908, IN29[4], w928, w929);
  FullAdder U249 (w929, w910, IN30[3], w930, w931);
  FullAdder U250 (w931, w912, IN31[2], w932, w933);
  FullAdder U251 (w933, w914, IN32[1], w934, w935);
  FullAdder U252 (w935, w915, IN33[0], w936, w937);
  HalfAdder U253 (w918, IN24[10], Out1[24], w939);
  FullAdder U254 (w939, w920, IN25[9], w940, w941);
  FullAdder U255 (w941, w922, IN26[8], w942, w943);
  FullAdder U256 (w943, w924, IN27[7], w944, w945);
  FullAdder U257 (w945, w926, IN28[6], w946, w947);
  FullAdder U258 (w947, w928, IN29[5], w948, w949);
  FullAdder U259 (w949, w930, IN30[4], w950, w951);
  FullAdder U260 (w951, w932, IN31[3], w952, w953);
  FullAdder U261 (w953, w934, IN32[2], w954, w955);
  FullAdder U262 (w955, w936, IN33[1], w956, w957);
  FullAdder U263 (w957, w937, IN34[0], w958, w959);
  HalfAdder U264 (w940, IN25[10], Out1[25], w961);
  FullAdder U265 (w961, w942, IN26[9], w962, w963);
  FullAdder U266 (w963, w944, IN27[8], w964, w965);
  FullAdder U267 (w965, w946, IN28[7], w966, w967);
  FullAdder U268 (w967, w948, IN29[6], w968, w969);
  FullAdder U269 (w969, w950, IN30[5], w970, w971);
  FullAdder U270 (w971, w952, IN31[4], w972, w973);
  FullAdder U271 (w973, w954, IN32[3], w974, w975);
  FullAdder U272 (w975, w956, IN33[2], w976, w977);
  FullAdder U273 (w977, w958, IN34[1], w978, w979);
  FullAdder U274 (w979, w959, IN35[0], w980, w981);
  HalfAdder U275 (w962, IN26[10], Out1[26], w983);
  FullAdder U276 (w983, w964, IN27[9], w984, w985);
  FullAdder U277 (w985, w966, IN28[8], w986, w987);
  FullAdder U278 (w987, w968, IN29[7], w988, w989);
  FullAdder U279 (w989, w970, IN30[6], w990, w991);
  FullAdder U280 (w991, w972, IN31[5], w992, w993);
  FullAdder U281 (w993, w974, IN32[4], w994, w995);
  FullAdder U282 (w995, w976, IN33[3], w996, w997);
  FullAdder U283 (w997, w978, IN34[2], w998, w999);
  FullAdder U284 (w999, w980, IN35[1], w1000, w1001);
  FullAdder U285 (w1001, w981, IN36[0], w1002, w1003);
  HalfAdder U286 (w984, IN27[10], Out1[27], w1005);
  FullAdder U287 (w1005, w986, IN28[9], w1006, w1007);
  FullAdder U288 (w1007, w988, IN29[8], w1008, w1009);
  FullAdder U289 (w1009, w990, IN30[7], w1010, w1011);
  FullAdder U290 (w1011, w992, IN31[6], w1012, w1013);
  FullAdder U291 (w1013, w994, IN32[5], w1014, w1015);
  FullAdder U292 (w1015, w996, IN33[4], w1016, w1017);
  FullAdder U293 (w1017, w998, IN34[3], w1018, w1019);
  FullAdder U294 (w1019, w1000, IN35[2], w1020, w1021);
  FullAdder U295 (w1021, w1002, IN36[1], w1022, w1023);
  FullAdder U296 (w1023, w1003, IN37[0], w1024, w1025);
  HalfAdder U297 (w1006, IN28[10], Out1[28], w1027);
  FullAdder U298 (w1027, w1008, IN29[9], w1028, w1029);
  FullAdder U299 (w1029, w1010, IN30[8], w1030, w1031);
  FullAdder U300 (w1031, w1012, IN31[7], w1032, w1033);
  FullAdder U301 (w1033, w1014, IN32[6], w1034, w1035);
  FullAdder U302 (w1035, w1016, IN33[5], w1036, w1037);
  FullAdder U303 (w1037, w1018, IN34[4], w1038, w1039);
  FullAdder U304 (w1039, w1020, IN35[3], w1040, w1041);
  FullAdder U305 (w1041, w1022, IN36[2], w1042, w1043);
  FullAdder U306 (w1043, w1024, IN37[1], w1044, w1045);
  FullAdder U307 (w1045, w1025, IN38[0], w1046, w1047);
  HalfAdder U308 (w1028, IN29[10], Out1[29], w1049);
  FullAdder U309 (w1049, w1030, IN30[9], w1050, w1051);
  FullAdder U310 (w1051, w1032, IN31[8], w1052, w1053);
  FullAdder U311 (w1053, w1034, IN32[7], w1054, w1055);
  FullAdder U312 (w1055, w1036, IN33[6], w1056, w1057);
  FullAdder U313 (w1057, w1038, IN34[5], w1058, w1059);
  FullAdder U314 (w1059, w1040, IN35[4], w1060, w1061);
  FullAdder U315 (w1061, w1042, IN36[3], w1062, w1063);
  FullAdder U316 (w1063, w1044, IN37[2], w1064, w1065);
  FullAdder U317 (w1065, w1046, IN38[1], w1066, w1067);
  FullAdder U318 (w1067, w1047, IN39[0], w1068, w1069);
  HalfAdder U319 (w1050, IN30[10], Out1[30], w1071);
  FullAdder U320 (w1071, w1052, IN31[9], w1072, w1073);
  FullAdder U321 (w1073, w1054, IN32[8], w1074, w1075);
  FullAdder U322 (w1075, w1056, IN33[7], w1076, w1077);
  FullAdder U323 (w1077, w1058, IN34[6], w1078, w1079);
  FullAdder U324 (w1079, w1060, IN35[5], w1080, w1081);
  FullAdder U325 (w1081, w1062, IN36[4], w1082, w1083);
  FullAdder U326 (w1083, w1064, IN37[3], w1084, w1085);
  FullAdder U327 (w1085, w1066, IN38[2], w1086, w1087);
  FullAdder U328 (w1087, w1068, IN39[1], w1088, w1089);
  FullAdder U329 (w1089, w1069, IN40[0], w1090, w1091);
  HalfAdder U330 (w1072, IN31[10], Out1[31], w1093);
  FullAdder U331 (w1093, w1074, IN32[9], w1094, w1095);
  FullAdder U332 (w1095, w1076, IN33[8], w1096, w1097);
  FullAdder U333 (w1097, w1078, IN34[7], w1098, w1099);
  FullAdder U334 (w1099, w1080, IN35[6], w1100, w1101);
  FullAdder U335 (w1101, w1082, IN36[5], w1102, w1103);
  FullAdder U336 (w1103, w1084, IN37[4], w1104, w1105);
  FullAdder U337 (w1105, w1086, IN38[3], w1106, w1107);
  FullAdder U338 (w1107, w1088, IN39[2], w1108, w1109);
  FullAdder U339 (w1109, w1090, IN40[1], w1110, w1111);
  FullAdder U340 (w1111, w1091, IN41[0], w1112, w1113);
  HalfAdder U341 (w1094, IN32[10], Out1[32], w1115);
  FullAdder U342 (w1115, w1096, IN33[9], w1116, w1117);
  FullAdder U343 (w1117, w1098, IN34[8], w1118, w1119);
  FullAdder U344 (w1119, w1100, IN35[7], w1120, w1121);
  FullAdder U345 (w1121, w1102, IN36[6], w1122, w1123);
  FullAdder U346 (w1123, w1104, IN37[5], w1124, w1125);
  FullAdder U347 (w1125, w1106, IN38[4], w1126, w1127);
  FullAdder U348 (w1127, w1108, IN39[3], w1128, w1129);
  FullAdder U349 (w1129, w1110, IN40[2], w1130, w1131);
  FullAdder U350 (w1131, w1112, IN41[1], w1132, w1133);
  FullAdder U351 (w1133, w1113, IN42[0], w1134, w1135);
  HalfAdder U352 (w1116, IN33[10], Out1[33], w1137);
  FullAdder U353 (w1137, w1118, IN34[9], w1138, w1139);
  FullAdder U354 (w1139, w1120, IN35[8], w1140, w1141);
  FullAdder U355 (w1141, w1122, IN36[7], w1142, w1143);
  FullAdder U356 (w1143, w1124, IN37[6], w1144, w1145);
  FullAdder U357 (w1145, w1126, IN38[5], w1146, w1147);
  FullAdder U358 (w1147, w1128, IN39[4], w1148, w1149);
  FullAdder U359 (w1149, w1130, IN40[3], w1150, w1151);
  FullAdder U360 (w1151, w1132, IN41[2], w1152, w1153);
  FullAdder U361 (w1153, w1134, IN42[1], w1154, w1155);
  FullAdder U362 (w1155, w1135, IN43[0], w1156, w1157);
  HalfAdder U363 (w1138, IN34[10], Out1[34], w1159);
  FullAdder U364 (w1159, w1140, IN35[9], w1160, w1161);
  FullAdder U365 (w1161, w1142, IN36[8], w1162, w1163);
  FullAdder U366 (w1163, w1144, IN37[7], w1164, w1165);
  FullAdder U367 (w1165, w1146, IN38[6], w1166, w1167);
  FullAdder U368 (w1167, w1148, IN39[5], w1168, w1169);
  FullAdder U369 (w1169, w1150, IN40[4], w1170, w1171);
  FullAdder U370 (w1171, w1152, IN41[3], w1172, w1173);
  FullAdder U371 (w1173, w1154, IN42[2], w1174, w1175);
  FullAdder U372 (w1175, w1156, IN43[1], w1176, w1177);
  FullAdder U373 (w1177, w1157, IN44[0], w1178, w1179);
  HalfAdder U374 (w1160, IN35[10], Out1[35], w1181);
  FullAdder U375 (w1181, w1162, IN36[9], Out1[36], w1183);
  FullAdder U376 (w1183, w1164, IN37[8], Out1[37], w1185);
  FullAdder U377 (w1185, w1166, IN38[7], Out1[38], w1187);
  FullAdder U378 (w1187, w1168, IN39[6], Out1[39], w1189);
  FullAdder U379 (w1189, w1170, IN40[5], Out1[40], w1191);
  FullAdder U380 (w1191, w1172, IN41[4], Out1[41], w1193);
  FullAdder U381 (w1193, w1174, IN42[3], Out1[42], w1195);
  FullAdder U382 (w1195, w1176, IN43[2], Out1[43], w1197);
  FullAdder U383 (w1197, w1178, IN44[1], Out1[44], w1199);
  FullAdder U384 (w1199, w1179, IN45[0], Out1[45], Out1[46]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN12[11];
  assign Out2[1] = IN13[11];
  assign Out2[2] = IN14[11];
  assign Out2[3] = IN15[11];
  assign Out2[4] = IN16[11];
  assign Out2[5] = IN17[11];
  assign Out2[6] = IN18[11];
  assign Out2[7] = IN19[11];
  assign Out2[8] = IN20[11];
  assign Out2[9] = IN21[11];
  assign Out2[10] = IN22[11];
  assign Out2[11] = IN23[11];
  assign Out2[12] = IN24[11];
  assign Out2[13] = IN25[11];
  assign Out2[14] = IN26[11];
  assign Out2[15] = IN27[11];
  assign Out2[16] = IN28[11];
  assign Out2[17] = IN29[11];
  assign Out2[18] = IN30[11];
  assign Out2[19] = IN31[11];
  assign Out2[20] = IN32[11];
  assign Out2[21] = IN33[11];
  assign Out2[22] = IN34[11];
  assign Out2[23] = IN35[11];
  assign Out2[24] = IN36[10];
  assign Out2[25] = IN37[9];
  assign Out2[26] = IN38[8];
  assign Out2[27] = IN39[7];
  assign Out2[28] = IN40[6];
  assign Out2[29] = IN41[5];
  assign Out2[30] = IN42[4];
  assign Out2[31] = IN43[3];
  assign Out2[32] = IN44[2];
  assign Out2[33] = IN45[1];
  assign Out2[34] = IN46[0];

endmodule
module RC_35_35(IN1, IN2, Out);
  input [34:0] IN1;
  input [34:0] IN2;
  output [35:0] Out;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w71);
  FullAdder U1 (IN1[1], IN2[1], w71, Out[1], w73);
  FullAdder U2 (IN1[2], IN2[2], w73, Out[2], w75);
  FullAdder U3 (IN1[3], IN2[3], w75, Out[3], w77);
  FullAdder U4 (IN1[4], IN2[4], w77, Out[4], w79);
  FullAdder U5 (IN1[5], IN2[5], w79, Out[5], w81);
  FullAdder U6 (IN1[6], IN2[6], w81, Out[6], w83);
  FullAdder U7 (IN1[7], IN2[7], w83, Out[7], w85);
  FullAdder U8 (IN1[8], IN2[8], w85, Out[8], w87);
  FullAdder U9 (IN1[9], IN2[9], w87, Out[9], w89);
  FullAdder U10 (IN1[10], IN2[10], w89, Out[10], w91);
  FullAdder U11 (IN1[11], IN2[11], w91, Out[11], w93);
  FullAdder U12 (IN1[12], IN2[12], w93, Out[12], w95);
  FullAdder U13 (IN1[13], IN2[13], w95, Out[13], w97);
  FullAdder U14 (IN1[14], IN2[14], w97, Out[14], w99);
  FullAdder U15 (IN1[15], IN2[15], w99, Out[15], w101);
  FullAdder U16 (IN1[16], IN2[16], w101, Out[16], w103);
  FullAdder U17 (IN1[17], IN2[17], w103, Out[17], w105);
  FullAdder U18 (IN1[18], IN2[18], w105, Out[18], w107);
  FullAdder U19 (IN1[19], IN2[19], w107, Out[19], w109);
  FullAdder U20 (IN1[20], IN2[20], w109, Out[20], w111);
  FullAdder U21 (IN1[21], IN2[21], w111, Out[21], w113);
  FullAdder U22 (IN1[22], IN2[22], w113, Out[22], w115);
  FullAdder U23 (IN1[23], IN2[23], w115, Out[23], w117);
  FullAdder U24 (IN1[24], IN2[24], w117, Out[24], w119);
  FullAdder U25 (IN1[25], IN2[25], w119, Out[25], w121);
  FullAdder U26 (IN1[26], IN2[26], w121, Out[26], w123);
  FullAdder U27 (IN1[27], IN2[27], w123, Out[27], w125);
  FullAdder U28 (IN1[28], IN2[28], w125, Out[28], w127);
  FullAdder U29 (IN1[29], IN2[29], w127, Out[29], w129);
  FullAdder U30 (IN1[30], IN2[30], w129, Out[30], w131);
  FullAdder U31 (IN1[31], IN2[31], w131, Out[31], w133);
  FullAdder U32 (IN1[32], IN2[32], w133, Out[32], w135);
  FullAdder U33 (IN1[33], IN2[33], w135, Out[33], w137);
  FullAdder U34 (IN1[34], IN2[34], w137, Out[34], Out[35]);

endmodule
module NR_12_36(IN1, IN2, Out);
  input [11:0] IN1;
  input [35:0] IN2;
  output [47:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [11:0] P12;
  wire [11:0] P13;
  wire [11:0] P14;
  wire [11:0] P15;
  wire [11:0] P16;
  wire [11:0] P17;
  wire [11:0] P18;
  wire [11:0] P19;
  wire [11:0] P20;
  wire [11:0] P21;
  wire [11:0] P22;
  wire [11:0] P23;
  wire [11:0] P24;
  wire [11:0] P25;
  wire [11:0] P26;
  wire [11:0] P27;
  wire [11:0] P28;
  wire [11:0] P29;
  wire [11:0] P30;
  wire [11:0] P31;
  wire [11:0] P32;
  wire [11:0] P33;
  wire [11:0] P34;
  wire [11:0] P35;
  wire [10:0] P36;
  wire [9:0] P37;
  wire [8:0] P38;
  wire [7:0] P39;
  wire [6:0] P40;
  wire [5:0] P41;
  wire [4:0] P42;
  wire [3:0] P43;
  wire [2:0] P44;
  wire [1:0] P45;
  wire [0:0] P46;
  wire [46:0] R1;
  wire [34:0] R2;
  wire [47:0] aOut;
  U_SP_12_36 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, R1, R2);
  RC_35_35 S2 (R1[46:12], R2, aOut[47:12]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign Out = aOut[47:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
