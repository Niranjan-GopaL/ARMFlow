
module customAdder33_0(
    input [32 : 0] A,
    input [32 : 0] B,
    output [33 : 0] Sum
);

    assign Sum = A+B;

endmodule
