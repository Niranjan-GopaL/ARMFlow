//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 61
  second input length: 4
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_61_4(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63);
  input [60:0] IN1;
  input [3:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [3:0] P4;
  output [3:0] P5;
  output [3:0] P6;
  output [3:0] P7;
  output [3:0] P8;
  output [3:0] P9;
  output [3:0] P10;
  output [3:0] P11;
  output [3:0] P12;
  output [3:0] P13;
  output [3:0] P14;
  output [3:0] P15;
  output [3:0] P16;
  output [3:0] P17;
  output [3:0] P18;
  output [3:0] P19;
  output [3:0] P20;
  output [3:0] P21;
  output [3:0] P22;
  output [3:0] P23;
  output [3:0] P24;
  output [3:0] P25;
  output [3:0] P26;
  output [3:0] P27;
  output [3:0] P28;
  output [3:0] P29;
  output [3:0] P30;
  output [3:0] P31;
  output [3:0] P32;
  output [3:0] P33;
  output [3:0] P34;
  output [3:0] P35;
  output [3:0] P36;
  output [3:0] P37;
  output [3:0] P38;
  output [3:0] P39;
  output [3:0] P40;
  output [3:0] P41;
  output [3:0] P42;
  output [3:0] P43;
  output [3:0] P44;
  output [3:0] P45;
  output [3:0] P46;
  output [3:0] P47;
  output [3:0] P48;
  output [3:0] P49;
  output [3:0] P50;
  output [3:0] P51;
  output [3:0] P52;
  output [3:0] P53;
  output [3:0] P54;
  output [3:0] P55;
  output [3:0] P56;
  output [3:0] P57;
  output [3:0] P58;
  output [3:0] P59;
  output [3:0] P60;
  output [2:0] P61;
  output [1:0] P62;
  output [0:0] P63;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[0] = IN1[1]&IN2[3];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[1] = IN1[2]&IN2[2];
  assign P5[0] = IN1[2]&IN2[3];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[2] = IN1[3]&IN2[1];
  assign P5[1] = IN1[3]&IN2[2];
  assign P6[0] = IN1[3]&IN2[3];
  assign P4[3] = IN1[4]&IN2[0];
  assign P5[2] = IN1[4]&IN2[1];
  assign P6[1] = IN1[4]&IN2[2];
  assign P7[0] = IN1[4]&IN2[3];
  assign P5[3] = IN1[5]&IN2[0];
  assign P6[2] = IN1[5]&IN2[1];
  assign P7[1] = IN1[5]&IN2[2];
  assign P8[0] = IN1[5]&IN2[3];
  assign P6[3] = IN1[6]&IN2[0];
  assign P7[2] = IN1[6]&IN2[1];
  assign P8[1] = IN1[6]&IN2[2];
  assign P9[0] = IN1[6]&IN2[3];
  assign P7[3] = IN1[7]&IN2[0];
  assign P8[2] = IN1[7]&IN2[1];
  assign P9[1] = IN1[7]&IN2[2];
  assign P10[0] = IN1[7]&IN2[3];
  assign P8[3] = IN1[8]&IN2[0];
  assign P9[2] = IN1[8]&IN2[1];
  assign P10[1] = IN1[8]&IN2[2];
  assign P11[0] = IN1[8]&IN2[3];
  assign P9[3] = IN1[9]&IN2[0];
  assign P10[2] = IN1[9]&IN2[1];
  assign P11[1] = IN1[9]&IN2[2];
  assign P12[0] = IN1[9]&IN2[3];
  assign P10[3] = IN1[10]&IN2[0];
  assign P11[2] = IN1[10]&IN2[1];
  assign P12[1] = IN1[10]&IN2[2];
  assign P13[0] = IN1[10]&IN2[3];
  assign P11[3] = IN1[11]&IN2[0];
  assign P12[2] = IN1[11]&IN2[1];
  assign P13[1] = IN1[11]&IN2[2];
  assign P14[0] = IN1[11]&IN2[3];
  assign P12[3] = IN1[12]&IN2[0];
  assign P13[2] = IN1[12]&IN2[1];
  assign P14[1] = IN1[12]&IN2[2];
  assign P15[0] = IN1[12]&IN2[3];
  assign P13[3] = IN1[13]&IN2[0];
  assign P14[2] = IN1[13]&IN2[1];
  assign P15[1] = IN1[13]&IN2[2];
  assign P16[0] = IN1[13]&IN2[3];
  assign P14[3] = IN1[14]&IN2[0];
  assign P15[2] = IN1[14]&IN2[1];
  assign P16[1] = IN1[14]&IN2[2];
  assign P17[0] = IN1[14]&IN2[3];
  assign P15[3] = IN1[15]&IN2[0];
  assign P16[2] = IN1[15]&IN2[1];
  assign P17[1] = IN1[15]&IN2[2];
  assign P18[0] = IN1[15]&IN2[3];
  assign P16[3] = IN1[16]&IN2[0];
  assign P17[2] = IN1[16]&IN2[1];
  assign P18[1] = IN1[16]&IN2[2];
  assign P19[0] = IN1[16]&IN2[3];
  assign P17[3] = IN1[17]&IN2[0];
  assign P18[2] = IN1[17]&IN2[1];
  assign P19[1] = IN1[17]&IN2[2];
  assign P20[0] = IN1[17]&IN2[3];
  assign P18[3] = IN1[18]&IN2[0];
  assign P19[2] = IN1[18]&IN2[1];
  assign P20[1] = IN1[18]&IN2[2];
  assign P21[0] = IN1[18]&IN2[3];
  assign P19[3] = IN1[19]&IN2[0];
  assign P20[2] = IN1[19]&IN2[1];
  assign P21[1] = IN1[19]&IN2[2];
  assign P22[0] = IN1[19]&IN2[3];
  assign P20[3] = IN1[20]&IN2[0];
  assign P21[2] = IN1[20]&IN2[1];
  assign P22[1] = IN1[20]&IN2[2];
  assign P23[0] = IN1[20]&IN2[3];
  assign P21[3] = IN1[21]&IN2[0];
  assign P22[2] = IN1[21]&IN2[1];
  assign P23[1] = IN1[21]&IN2[2];
  assign P24[0] = IN1[21]&IN2[3];
  assign P22[3] = IN1[22]&IN2[0];
  assign P23[2] = IN1[22]&IN2[1];
  assign P24[1] = IN1[22]&IN2[2];
  assign P25[0] = IN1[22]&IN2[3];
  assign P23[3] = IN1[23]&IN2[0];
  assign P24[2] = IN1[23]&IN2[1];
  assign P25[1] = IN1[23]&IN2[2];
  assign P26[0] = IN1[23]&IN2[3];
  assign P24[3] = IN1[24]&IN2[0];
  assign P25[2] = IN1[24]&IN2[1];
  assign P26[1] = IN1[24]&IN2[2];
  assign P27[0] = IN1[24]&IN2[3];
  assign P25[3] = IN1[25]&IN2[0];
  assign P26[2] = IN1[25]&IN2[1];
  assign P27[1] = IN1[25]&IN2[2];
  assign P28[0] = IN1[25]&IN2[3];
  assign P26[3] = IN1[26]&IN2[0];
  assign P27[2] = IN1[26]&IN2[1];
  assign P28[1] = IN1[26]&IN2[2];
  assign P29[0] = IN1[26]&IN2[3];
  assign P27[3] = IN1[27]&IN2[0];
  assign P28[2] = IN1[27]&IN2[1];
  assign P29[1] = IN1[27]&IN2[2];
  assign P30[0] = IN1[27]&IN2[3];
  assign P28[3] = IN1[28]&IN2[0];
  assign P29[2] = IN1[28]&IN2[1];
  assign P30[1] = IN1[28]&IN2[2];
  assign P31[0] = IN1[28]&IN2[3];
  assign P29[3] = IN1[29]&IN2[0];
  assign P30[2] = IN1[29]&IN2[1];
  assign P31[1] = IN1[29]&IN2[2];
  assign P32[0] = IN1[29]&IN2[3];
  assign P30[3] = IN1[30]&IN2[0];
  assign P31[2] = IN1[30]&IN2[1];
  assign P32[1] = IN1[30]&IN2[2];
  assign P33[0] = IN1[30]&IN2[3];
  assign P31[3] = IN1[31]&IN2[0];
  assign P32[2] = IN1[31]&IN2[1];
  assign P33[1] = IN1[31]&IN2[2];
  assign P34[0] = IN1[31]&IN2[3];
  assign P32[3] = IN1[32]&IN2[0];
  assign P33[2] = IN1[32]&IN2[1];
  assign P34[1] = IN1[32]&IN2[2];
  assign P35[0] = IN1[32]&IN2[3];
  assign P33[3] = IN1[33]&IN2[0];
  assign P34[2] = IN1[33]&IN2[1];
  assign P35[1] = IN1[33]&IN2[2];
  assign P36[0] = IN1[33]&IN2[3];
  assign P34[3] = IN1[34]&IN2[0];
  assign P35[2] = IN1[34]&IN2[1];
  assign P36[1] = IN1[34]&IN2[2];
  assign P37[0] = IN1[34]&IN2[3];
  assign P35[3] = IN1[35]&IN2[0];
  assign P36[2] = IN1[35]&IN2[1];
  assign P37[1] = IN1[35]&IN2[2];
  assign P38[0] = IN1[35]&IN2[3];
  assign P36[3] = IN1[36]&IN2[0];
  assign P37[2] = IN1[36]&IN2[1];
  assign P38[1] = IN1[36]&IN2[2];
  assign P39[0] = IN1[36]&IN2[3];
  assign P37[3] = IN1[37]&IN2[0];
  assign P38[2] = IN1[37]&IN2[1];
  assign P39[1] = IN1[37]&IN2[2];
  assign P40[0] = IN1[37]&IN2[3];
  assign P38[3] = IN1[38]&IN2[0];
  assign P39[2] = IN1[38]&IN2[1];
  assign P40[1] = IN1[38]&IN2[2];
  assign P41[0] = IN1[38]&IN2[3];
  assign P39[3] = IN1[39]&IN2[0];
  assign P40[2] = IN1[39]&IN2[1];
  assign P41[1] = IN1[39]&IN2[2];
  assign P42[0] = IN1[39]&IN2[3];
  assign P40[3] = IN1[40]&IN2[0];
  assign P41[2] = IN1[40]&IN2[1];
  assign P42[1] = IN1[40]&IN2[2];
  assign P43[0] = IN1[40]&IN2[3];
  assign P41[3] = IN1[41]&IN2[0];
  assign P42[2] = IN1[41]&IN2[1];
  assign P43[1] = IN1[41]&IN2[2];
  assign P44[0] = IN1[41]&IN2[3];
  assign P42[3] = IN1[42]&IN2[0];
  assign P43[2] = IN1[42]&IN2[1];
  assign P44[1] = IN1[42]&IN2[2];
  assign P45[0] = IN1[42]&IN2[3];
  assign P43[3] = IN1[43]&IN2[0];
  assign P44[2] = IN1[43]&IN2[1];
  assign P45[1] = IN1[43]&IN2[2];
  assign P46[0] = IN1[43]&IN2[3];
  assign P44[3] = IN1[44]&IN2[0];
  assign P45[2] = IN1[44]&IN2[1];
  assign P46[1] = IN1[44]&IN2[2];
  assign P47[0] = IN1[44]&IN2[3];
  assign P45[3] = IN1[45]&IN2[0];
  assign P46[2] = IN1[45]&IN2[1];
  assign P47[1] = IN1[45]&IN2[2];
  assign P48[0] = IN1[45]&IN2[3];
  assign P46[3] = IN1[46]&IN2[0];
  assign P47[2] = IN1[46]&IN2[1];
  assign P48[1] = IN1[46]&IN2[2];
  assign P49[0] = IN1[46]&IN2[3];
  assign P47[3] = IN1[47]&IN2[0];
  assign P48[2] = IN1[47]&IN2[1];
  assign P49[1] = IN1[47]&IN2[2];
  assign P50[0] = IN1[47]&IN2[3];
  assign P48[3] = IN1[48]&IN2[0];
  assign P49[2] = IN1[48]&IN2[1];
  assign P50[1] = IN1[48]&IN2[2];
  assign P51[0] = IN1[48]&IN2[3];
  assign P49[3] = IN1[49]&IN2[0];
  assign P50[2] = IN1[49]&IN2[1];
  assign P51[1] = IN1[49]&IN2[2];
  assign P52[0] = IN1[49]&IN2[3];
  assign P50[3] = IN1[50]&IN2[0];
  assign P51[2] = IN1[50]&IN2[1];
  assign P52[1] = IN1[50]&IN2[2];
  assign P53[0] = IN1[50]&IN2[3];
  assign P51[3] = IN1[51]&IN2[0];
  assign P52[2] = IN1[51]&IN2[1];
  assign P53[1] = IN1[51]&IN2[2];
  assign P54[0] = IN1[51]&IN2[3];
  assign P52[3] = IN1[52]&IN2[0];
  assign P53[2] = IN1[52]&IN2[1];
  assign P54[1] = IN1[52]&IN2[2];
  assign P55[0] = IN1[52]&IN2[3];
  assign P53[3] = IN1[53]&IN2[0];
  assign P54[2] = IN1[53]&IN2[1];
  assign P55[1] = IN1[53]&IN2[2];
  assign P56[0] = IN1[53]&IN2[3];
  assign P54[3] = IN1[54]&IN2[0];
  assign P55[2] = IN1[54]&IN2[1];
  assign P56[1] = IN1[54]&IN2[2];
  assign P57[0] = IN1[54]&IN2[3];
  assign P55[3] = IN1[55]&IN2[0];
  assign P56[2] = IN1[55]&IN2[1];
  assign P57[1] = IN1[55]&IN2[2];
  assign P58[0] = IN1[55]&IN2[3];
  assign P56[3] = IN1[56]&IN2[0];
  assign P57[2] = IN1[56]&IN2[1];
  assign P58[1] = IN1[56]&IN2[2];
  assign P59[0] = IN1[56]&IN2[3];
  assign P57[3] = IN1[57]&IN2[0];
  assign P58[2] = IN1[57]&IN2[1];
  assign P59[1] = IN1[57]&IN2[2];
  assign P60[0] = IN1[57]&IN2[3];
  assign P58[3] = IN1[58]&IN2[0];
  assign P59[2] = IN1[58]&IN2[1];
  assign P60[1] = IN1[58]&IN2[2];
  assign P61[0] = IN1[58]&IN2[3];
  assign P59[3] = IN1[59]&IN2[0];
  assign P60[2] = IN1[59]&IN2[1];
  assign P61[1] = IN1[59]&IN2[2];
  assign P62[0] = IN1[59]&IN2[3];
  assign P60[3] = IN1[60]&IN2[0];
  assign P61[2] = IN1[60]&IN2[1];
  assign P62[1] = IN1[60]&IN2[2];
  assign P63[0] = IN1[60]&IN2[3];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [3:0] IN4;
  input [3:0] IN5;
  input [3:0] IN6;
  input [3:0] IN7;
  input [3:0] IN8;
  input [3:0] IN9;
  input [3:0] IN10;
  input [3:0] IN11;
  input [3:0] IN12;
  input [3:0] IN13;
  input [3:0] IN14;
  input [3:0] IN15;
  input [3:0] IN16;
  input [3:0] IN17;
  input [3:0] IN18;
  input [3:0] IN19;
  input [3:0] IN20;
  input [3:0] IN21;
  input [3:0] IN22;
  input [3:0] IN23;
  input [3:0] IN24;
  input [3:0] IN25;
  input [3:0] IN26;
  input [3:0] IN27;
  input [3:0] IN28;
  input [3:0] IN29;
  input [3:0] IN30;
  input [3:0] IN31;
  input [3:0] IN32;
  input [3:0] IN33;
  input [3:0] IN34;
  input [3:0] IN35;
  input [3:0] IN36;
  input [3:0] IN37;
  input [3:0] IN38;
  input [3:0] IN39;
  input [3:0] IN40;
  input [3:0] IN41;
  input [3:0] IN42;
  input [3:0] IN43;
  input [3:0] IN44;
  input [3:0] IN45;
  input [3:0] IN46;
  input [3:0] IN47;
  input [3:0] IN48;
  input [3:0] IN49;
  input [3:0] IN50;
  input [3:0] IN51;
  input [3:0] IN52;
  input [3:0] IN53;
  input [3:0] IN54;
  input [3:0] IN55;
  input [3:0] IN56;
  input [3:0] IN57;
  input [3:0] IN58;
  input [3:0] IN59;
  input [3:0] IN60;
  input [2:0] IN61;
  input [1:0] IN62;
  input [0:0] IN63;
  output [63:0] Out1;
  output [2:0] Out2;
  wire w245;
  wire w246;
  wire w247;
  wire w248;
  wire w249;
  wire w250;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w485;
  wire w487;
  wire w489;
  wire w491;
  wire w493;
  wire w495;
  wire w497;
  wire w499;
  wire w501;
  wire w503;
  wire w505;
  wire w507;
  wire w509;
  wire w511;
  wire w513;
  wire w515;
  wire w517;
  wire w519;
  wire w521;
  wire w523;
  wire w525;
  wire w527;
  wire w529;
  wire w531;
  wire w533;
  wire w535;
  wire w537;
  wire w539;
  wire w541;
  wire w543;
  wire w545;
  wire w547;
  wire w549;
  wire w551;
  wire w553;
  wire w555;
  wire w557;
  wire w559;
  wire w561;
  wire w563;
  wire w565;
  wire w567;
  wire w569;
  wire w571;
  wire w573;
  wire w575;
  wire w577;
  wire w579;
  wire w581;
  wire w583;
  wire w585;
  wire w587;
  wire w589;
  wire w591;
  wire w593;
  wire w595;
  wire w597;
  wire w599;
  wire w601;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w245);
  FullAdder U1 (w245, IN2[0], IN2[1], w246, w247);
  FullAdder U2 (w247, IN3[0], IN3[1], w248, w249);
  FullAdder U3 (w249, IN4[0], IN4[1], w250, w251);
  FullAdder U4 (w251, IN5[0], IN5[1], w252, w253);
  FullAdder U5 (w253, IN6[0], IN6[1], w254, w255);
  FullAdder U6 (w255, IN7[0], IN7[1], w256, w257);
  FullAdder U7 (w257, IN8[0], IN8[1], w258, w259);
  FullAdder U8 (w259, IN9[0], IN9[1], w260, w261);
  FullAdder U9 (w261, IN10[0], IN10[1], w262, w263);
  FullAdder U10 (w263, IN11[0], IN11[1], w264, w265);
  FullAdder U11 (w265, IN12[0], IN12[1], w266, w267);
  FullAdder U12 (w267, IN13[0], IN13[1], w268, w269);
  FullAdder U13 (w269, IN14[0], IN14[1], w270, w271);
  FullAdder U14 (w271, IN15[0], IN15[1], w272, w273);
  FullAdder U15 (w273, IN16[0], IN16[1], w274, w275);
  FullAdder U16 (w275, IN17[0], IN17[1], w276, w277);
  FullAdder U17 (w277, IN18[0], IN18[1], w278, w279);
  FullAdder U18 (w279, IN19[0], IN19[1], w280, w281);
  FullAdder U19 (w281, IN20[0], IN20[1], w282, w283);
  FullAdder U20 (w283, IN21[0], IN21[1], w284, w285);
  FullAdder U21 (w285, IN22[0], IN22[1], w286, w287);
  FullAdder U22 (w287, IN23[0], IN23[1], w288, w289);
  FullAdder U23 (w289, IN24[0], IN24[1], w290, w291);
  FullAdder U24 (w291, IN25[0], IN25[1], w292, w293);
  FullAdder U25 (w293, IN26[0], IN26[1], w294, w295);
  FullAdder U26 (w295, IN27[0], IN27[1], w296, w297);
  FullAdder U27 (w297, IN28[0], IN28[1], w298, w299);
  FullAdder U28 (w299, IN29[0], IN29[1], w300, w301);
  FullAdder U29 (w301, IN30[0], IN30[1], w302, w303);
  FullAdder U30 (w303, IN31[0], IN31[1], w304, w305);
  FullAdder U31 (w305, IN32[0], IN32[1], w306, w307);
  FullAdder U32 (w307, IN33[0], IN33[1], w308, w309);
  FullAdder U33 (w309, IN34[0], IN34[1], w310, w311);
  FullAdder U34 (w311, IN35[0], IN35[1], w312, w313);
  FullAdder U35 (w313, IN36[0], IN36[1], w314, w315);
  FullAdder U36 (w315, IN37[0], IN37[1], w316, w317);
  FullAdder U37 (w317, IN38[0], IN38[1], w318, w319);
  FullAdder U38 (w319, IN39[0], IN39[1], w320, w321);
  FullAdder U39 (w321, IN40[0], IN40[1], w322, w323);
  FullAdder U40 (w323, IN41[0], IN41[1], w324, w325);
  FullAdder U41 (w325, IN42[0], IN42[1], w326, w327);
  FullAdder U42 (w327, IN43[0], IN43[1], w328, w329);
  FullAdder U43 (w329, IN44[0], IN44[1], w330, w331);
  FullAdder U44 (w331, IN45[0], IN45[1], w332, w333);
  FullAdder U45 (w333, IN46[0], IN46[1], w334, w335);
  FullAdder U46 (w335, IN47[0], IN47[1], w336, w337);
  FullAdder U47 (w337, IN48[0], IN48[1], w338, w339);
  FullAdder U48 (w339, IN49[0], IN49[1], w340, w341);
  FullAdder U49 (w341, IN50[0], IN50[1], w342, w343);
  FullAdder U50 (w343, IN51[0], IN51[1], w344, w345);
  FullAdder U51 (w345, IN52[0], IN52[1], w346, w347);
  FullAdder U52 (w347, IN53[0], IN53[1], w348, w349);
  FullAdder U53 (w349, IN54[0], IN54[1], w350, w351);
  FullAdder U54 (w351, IN55[0], IN55[1], w352, w353);
  FullAdder U55 (w353, IN56[0], IN56[1], w354, w355);
  FullAdder U56 (w355, IN57[0], IN57[1], w356, w357);
  FullAdder U57 (w357, IN58[0], IN58[1], w358, w359);
  FullAdder U58 (w359, IN59[0], IN59[1], w360, w361);
  FullAdder U59 (w361, IN60[0], IN60[1], w362, w363);
  HalfAdder U60 (w246, IN2[2], Out1[2], w365);
  FullAdder U61 (w365, w248, IN3[2], w366, w367);
  FullAdder U62 (w367, w250, IN4[2], w368, w369);
  FullAdder U63 (w369, w252, IN5[2], w370, w371);
  FullAdder U64 (w371, w254, IN6[2], w372, w373);
  FullAdder U65 (w373, w256, IN7[2], w374, w375);
  FullAdder U66 (w375, w258, IN8[2], w376, w377);
  FullAdder U67 (w377, w260, IN9[2], w378, w379);
  FullAdder U68 (w379, w262, IN10[2], w380, w381);
  FullAdder U69 (w381, w264, IN11[2], w382, w383);
  FullAdder U70 (w383, w266, IN12[2], w384, w385);
  FullAdder U71 (w385, w268, IN13[2], w386, w387);
  FullAdder U72 (w387, w270, IN14[2], w388, w389);
  FullAdder U73 (w389, w272, IN15[2], w390, w391);
  FullAdder U74 (w391, w274, IN16[2], w392, w393);
  FullAdder U75 (w393, w276, IN17[2], w394, w395);
  FullAdder U76 (w395, w278, IN18[2], w396, w397);
  FullAdder U77 (w397, w280, IN19[2], w398, w399);
  FullAdder U78 (w399, w282, IN20[2], w400, w401);
  FullAdder U79 (w401, w284, IN21[2], w402, w403);
  FullAdder U80 (w403, w286, IN22[2], w404, w405);
  FullAdder U81 (w405, w288, IN23[2], w406, w407);
  FullAdder U82 (w407, w290, IN24[2], w408, w409);
  FullAdder U83 (w409, w292, IN25[2], w410, w411);
  FullAdder U84 (w411, w294, IN26[2], w412, w413);
  FullAdder U85 (w413, w296, IN27[2], w414, w415);
  FullAdder U86 (w415, w298, IN28[2], w416, w417);
  FullAdder U87 (w417, w300, IN29[2], w418, w419);
  FullAdder U88 (w419, w302, IN30[2], w420, w421);
  FullAdder U89 (w421, w304, IN31[2], w422, w423);
  FullAdder U90 (w423, w306, IN32[2], w424, w425);
  FullAdder U91 (w425, w308, IN33[2], w426, w427);
  FullAdder U92 (w427, w310, IN34[2], w428, w429);
  FullAdder U93 (w429, w312, IN35[2], w430, w431);
  FullAdder U94 (w431, w314, IN36[2], w432, w433);
  FullAdder U95 (w433, w316, IN37[2], w434, w435);
  FullAdder U96 (w435, w318, IN38[2], w436, w437);
  FullAdder U97 (w437, w320, IN39[2], w438, w439);
  FullAdder U98 (w439, w322, IN40[2], w440, w441);
  FullAdder U99 (w441, w324, IN41[2], w442, w443);
  FullAdder U100 (w443, w326, IN42[2], w444, w445);
  FullAdder U101 (w445, w328, IN43[2], w446, w447);
  FullAdder U102 (w447, w330, IN44[2], w448, w449);
  FullAdder U103 (w449, w332, IN45[2], w450, w451);
  FullAdder U104 (w451, w334, IN46[2], w452, w453);
  FullAdder U105 (w453, w336, IN47[2], w454, w455);
  FullAdder U106 (w455, w338, IN48[2], w456, w457);
  FullAdder U107 (w457, w340, IN49[2], w458, w459);
  FullAdder U108 (w459, w342, IN50[2], w460, w461);
  FullAdder U109 (w461, w344, IN51[2], w462, w463);
  FullAdder U110 (w463, w346, IN52[2], w464, w465);
  FullAdder U111 (w465, w348, IN53[2], w466, w467);
  FullAdder U112 (w467, w350, IN54[2], w468, w469);
  FullAdder U113 (w469, w352, IN55[2], w470, w471);
  FullAdder U114 (w471, w354, IN56[2], w472, w473);
  FullAdder U115 (w473, w356, IN57[2], w474, w475);
  FullAdder U116 (w475, w358, IN58[2], w476, w477);
  FullAdder U117 (w477, w360, IN59[2], w478, w479);
  FullAdder U118 (w479, w362, IN60[2], w480, w481);
  FullAdder U119 (w481, w363, IN61[0], w482, w483);
  HalfAdder U120 (w366, IN3[3], Out1[3], w485);
  FullAdder U121 (w485, w368, IN4[3], Out1[4], w487);
  FullAdder U122 (w487, w370, IN5[3], Out1[5], w489);
  FullAdder U123 (w489, w372, IN6[3], Out1[6], w491);
  FullAdder U124 (w491, w374, IN7[3], Out1[7], w493);
  FullAdder U125 (w493, w376, IN8[3], Out1[8], w495);
  FullAdder U126 (w495, w378, IN9[3], Out1[9], w497);
  FullAdder U127 (w497, w380, IN10[3], Out1[10], w499);
  FullAdder U128 (w499, w382, IN11[3], Out1[11], w501);
  FullAdder U129 (w501, w384, IN12[3], Out1[12], w503);
  FullAdder U130 (w503, w386, IN13[3], Out1[13], w505);
  FullAdder U131 (w505, w388, IN14[3], Out1[14], w507);
  FullAdder U132 (w507, w390, IN15[3], Out1[15], w509);
  FullAdder U133 (w509, w392, IN16[3], Out1[16], w511);
  FullAdder U134 (w511, w394, IN17[3], Out1[17], w513);
  FullAdder U135 (w513, w396, IN18[3], Out1[18], w515);
  FullAdder U136 (w515, w398, IN19[3], Out1[19], w517);
  FullAdder U137 (w517, w400, IN20[3], Out1[20], w519);
  FullAdder U138 (w519, w402, IN21[3], Out1[21], w521);
  FullAdder U139 (w521, w404, IN22[3], Out1[22], w523);
  FullAdder U140 (w523, w406, IN23[3], Out1[23], w525);
  FullAdder U141 (w525, w408, IN24[3], Out1[24], w527);
  FullAdder U142 (w527, w410, IN25[3], Out1[25], w529);
  FullAdder U143 (w529, w412, IN26[3], Out1[26], w531);
  FullAdder U144 (w531, w414, IN27[3], Out1[27], w533);
  FullAdder U145 (w533, w416, IN28[3], Out1[28], w535);
  FullAdder U146 (w535, w418, IN29[3], Out1[29], w537);
  FullAdder U147 (w537, w420, IN30[3], Out1[30], w539);
  FullAdder U148 (w539, w422, IN31[3], Out1[31], w541);
  FullAdder U149 (w541, w424, IN32[3], Out1[32], w543);
  FullAdder U150 (w543, w426, IN33[3], Out1[33], w545);
  FullAdder U151 (w545, w428, IN34[3], Out1[34], w547);
  FullAdder U152 (w547, w430, IN35[3], Out1[35], w549);
  FullAdder U153 (w549, w432, IN36[3], Out1[36], w551);
  FullAdder U154 (w551, w434, IN37[3], Out1[37], w553);
  FullAdder U155 (w553, w436, IN38[3], Out1[38], w555);
  FullAdder U156 (w555, w438, IN39[3], Out1[39], w557);
  FullAdder U157 (w557, w440, IN40[3], Out1[40], w559);
  FullAdder U158 (w559, w442, IN41[3], Out1[41], w561);
  FullAdder U159 (w561, w444, IN42[3], Out1[42], w563);
  FullAdder U160 (w563, w446, IN43[3], Out1[43], w565);
  FullAdder U161 (w565, w448, IN44[3], Out1[44], w567);
  FullAdder U162 (w567, w450, IN45[3], Out1[45], w569);
  FullAdder U163 (w569, w452, IN46[3], Out1[46], w571);
  FullAdder U164 (w571, w454, IN47[3], Out1[47], w573);
  FullAdder U165 (w573, w456, IN48[3], Out1[48], w575);
  FullAdder U166 (w575, w458, IN49[3], Out1[49], w577);
  FullAdder U167 (w577, w460, IN50[3], Out1[50], w579);
  FullAdder U168 (w579, w462, IN51[3], Out1[51], w581);
  FullAdder U169 (w581, w464, IN52[3], Out1[52], w583);
  FullAdder U170 (w583, w466, IN53[3], Out1[53], w585);
  FullAdder U171 (w585, w468, IN54[3], Out1[54], w587);
  FullAdder U172 (w587, w470, IN55[3], Out1[55], w589);
  FullAdder U173 (w589, w472, IN56[3], Out1[56], w591);
  FullAdder U174 (w591, w474, IN57[3], Out1[57], w593);
  FullAdder U175 (w593, w476, IN58[3], Out1[58], w595);
  FullAdder U176 (w595, w478, IN59[3], Out1[59], w597);
  FullAdder U177 (w597, w480, IN60[3], Out1[60], w599);
  FullAdder U178 (w599, w482, IN61[1], Out1[61], w601);
  FullAdder U179 (w601, w483, IN62[0], Out1[62], Out1[63]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN61[2];
  assign Out2[1] = IN62[1];
  assign Out2[2] = IN63[0];

endmodule
module RC_3_3(IN1, IN2, Out);
  input [2:0] IN1;
  input [2:0] IN2;
  output [3:0] Out;
  wire w7;
  wire w9;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w7);
  FullAdder U1 (IN1[1], IN2[1], w7, Out[1], w9);
  FullAdder U2 (IN1[2], IN2[2], w9, Out[2], Out[3]);

endmodule
module NR_61_4(IN1, IN2, Out);
  input [60:0] IN1;
  input [3:0] IN2;
  output [64:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [3:0] P4;
  wire [3:0] P5;
  wire [3:0] P6;
  wire [3:0] P7;
  wire [3:0] P8;
  wire [3:0] P9;
  wire [3:0] P10;
  wire [3:0] P11;
  wire [3:0] P12;
  wire [3:0] P13;
  wire [3:0] P14;
  wire [3:0] P15;
  wire [3:0] P16;
  wire [3:0] P17;
  wire [3:0] P18;
  wire [3:0] P19;
  wire [3:0] P20;
  wire [3:0] P21;
  wire [3:0] P22;
  wire [3:0] P23;
  wire [3:0] P24;
  wire [3:0] P25;
  wire [3:0] P26;
  wire [3:0] P27;
  wire [3:0] P28;
  wire [3:0] P29;
  wire [3:0] P30;
  wire [3:0] P31;
  wire [3:0] P32;
  wire [3:0] P33;
  wire [3:0] P34;
  wire [3:0] P35;
  wire [3:0] P36;
  wire [3:0] P37;
  wire [3:0] P38;
  wire [3:0] P39;
  wire [3:0] P40;
  wire [3:0] P41;
  wire [3:0] P42;
  wire [3:0] P43;
  wire [3:0] P44;
  wire [3:0] P45;
  wire [3:0] P46;
  wire [3:0] P47;
  wire [3:0] P48;
  wire [3:0] P49;
  wire [3:0] P50;
  wire [3:0] P51;
  wire [3:0] P52;
  wire [3:0] P53;
  wire [3:0] P54;
  wire [3:0] P55;
  wire [3:0] P56;
  wire [3:0] P57;
  wire [3:0] P58;
  wire [3:0] P59;
  wire [3:0] P60;
  wire [2:0] P61;
  wire [1:0] P62;
  wire [0:0] P63;
  wire [63:0] R1;
  wire [2:0] R2;
  wire [64:0] aOut;
  U_SP_61_4 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, R1, R2);
  RC_3_3 S2 (R1[63:61], R2, aOut[64:61]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign aOut[57] = R1[57];
  assign aOut[58] = R1[58];
  assign aOut[59] = R1[59];
  assign aOut[60] = R1[60];
  assign Out = aOut[64:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
