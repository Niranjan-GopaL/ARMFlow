
module customAdder62_0(
    input [61 : 0] A,
    input [61 : 0] B,
    output [62 : 0] Sum
);

    assign Sum = A+B;

endmodule
