
module customAdder63_0(
    input [62 : 0] A,
    input [62 : 0] B,
    output [63 : 0] Sum
);

    assign Sum = A+B;

endmodule
