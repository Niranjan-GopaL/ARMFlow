//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 26
  second input length: 38
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_26_38(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  input [25:0] IN1;
  input [37:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [25:0] P26;
  output [25:0] P27;
  output [25:0] P28;
  output [25:0] P29;
  output [25:0] P30;
  output [25:0] P31;
  output [25:0] P32;
  output [25:0] P33;
  output [25:0] P34;
  output [25:0] P35;
  output [25:0] P36;
  output [25:0] P37;
  output [24:0] P38;
  output [23:0] P39;
  output [22:0] P40;
  output [21:0] P41;
  output [20:0] P42;
  output [19:0] P43;
  output [18:0] P44;
  output [17:0] P45;
  output [16:0] P46;
  output [15:0] P47;
  output [14:0] P48;
  output [13:0] P49;
  output [12:0] P50;
  output [11:0] P51;
  output [10:0] P52;
  output [9:0] P53;
  output [8:0] P54;
  output [7:0] P55;
  output [6:0] P56;
  output [5:0] P57;
  output [4:0] P58;
  output [3:0] P59;
  output [2:0] P60;
  output [1:0] P61;
  output [0:0] P62;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[0] = IN1[1]&IN2[37];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[1] = IN1[2]&IN2[36];
  assign P39[0] = IN1[2]&IN2[37];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[2] = IN1[3]&IN2[35];
  assign P39[1] = IN1[3]&IN2[36];
  assign P40[0] = IN1[3]&IN2[37];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[3] = IN1[4]&IN2[34];
  assign P39[2] = IN1[4]&IN2[35];
  assign P40[1] = IN1[4]&IN2[36];
  assign P41[0] = IN1[4]&IN2[37];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[4] = IN1[5]&IN2[33];
  assign P39[3] = IN1[5]&IN2[34];
  assign P40[2] = IN1[5]&IN2[35];
  assign P41[1] = IN1[5]&IN2[36];
  assign P42[0] = IN1[5]&IN2[37];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[5] = IN1[6]&IN2[32];
  assign P39[4] = IN1[6]&IN2[33];
  assign P40[3] = IN1[6]&IN2[34];
  assign P41[2] = IN1[6]&IN2[35];
  assign P42[1] = IN1[6]&IN2[36];
  assign P43[0] = IN1[6]&IN2[37];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[6] = IN1[7]&IN2[31];
  assign P39[5] = IN1[7]&IN2[32];
  assign P40[4] = IN1[7]&IN2[33];
  assign P41[3] = IN1[7]&IN2[34];
  assign P42[2] = IN1[7]&IN2[35];
  assign P43[1] = IN1[7]&IN2[36];
  assign P44[0] = IN1[7]&IN2[37];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[7] = IN1[8]&IN2[30];
  assign P39[6] = IN1[8]&IN2[31];
  assign P40[5] = IN1[8]&IN2[32];
  assign P41[4] = IN1[8]&IN2[33];
  assign P42[3] = IN1[8]&IN2[34];
  assign P43[2] = IN1[8]&IN2[35];
  assign P44[1] = IN1[8]&IN2[36];
  assign P45[0] = IN1[8]&IN2[37];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[8] = IN1[9]&IN2[29];
  assign P39[7] = IN1[9]&IN2[30];
  assign P40[6] = IN1[9]&IN2[31];
  assign P41[5] = IN1[9]&IN2[32];
  assign P42[4] = IN1[9]&IN2[33];
  assign P43[3] = IN1[9]&IN2[34];
  assign P44[2] = IN1[9]&IN2[35];
  assign P45[1] = IN1[9]&IN2[36];
  assign P46[0] = IN1[9]&IN2[37];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[9] = IN1[10]&IN2[28];
  assign P39[8] = IN1[10]&IN2[29];
  assign P40[7] = IN1[10]&IN2[30];
  assign P41[6] = IN1[10]&IN2[31];
  assign P42[5] = IN1[10]&IN2[32];
  assign P43[4] = IN1[10]&IN2[33];
  assign P44[3] = IN1[10]&IN2[34];
  assign P45[2] = IN1[10]&IN2[35];
  assign P46[1] = IN1[10]&IN2[36];
  assign P47[0] = IN1[10]&IN2[37];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[10] = IN1[11]&IN2[27];
  assign P39[9] = IN1[11]&IN2[28];
  assign P40[8] = IN1[11]&IN2[29];
  assign P41[7] = IN1[11]&IN2[30];
  assign P42[6] = IN1[11]&IN2[31];
  assign P43[5] = IN1[11]&IN2[32];
  assign P44[4] = IN1[11]&IN2[33];
  assign P45[3] = IN1[11]&IN2[34];
  assign P46[2] = IN1[11]&IN2[35];
  assign P47[1] = IN1[11]&IN2[36];
  assign P48[0] = IN1[11]&IN2[37];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[11] = IN1[12]&IN2[26];
  assign P39[10] = IN1[12]&IN2[27];
  assign P40[9] = IN1[12]&IN2[28];
  assign P41[8] = IN1[12]&IN2[29];
  assign P42[7] = IN1[12]&IN2[30];
  assign P43[6] = IN1[12]&IN2[31];
  assign P44[5] = IN1[12]&IN2[32];
  assign P45[4] = IN1[12]&IN2[33];
  assign P46[3] = IN1[12]&IN2[34];
  assign P47[2] = IN1[12]&IN2[35];
  assign P48[1] = IN1[12]&IN2[36];
  assign P49[0] = IN1[12]&IN2[37];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[12] = IN1[13]&IN2[25];
  assign P39[11] = IN1[13]&IN2[26];
  assign P40[10] = IN1[13]&IN2[27];
  assign P41[9] = IN1[13]&IN2[28];
  assign P42[8] = IN1[13]&IN2[29];
  assign P43[7] = IN1[13]&IN2[30];
  assign P44[6] = IN1[13]&IN2[31];
  assign P45[5] = IN1[13]&IN2[32];
  assign P46[4] = IN1[13]&IN2[33];
  assign P47[3] = IN1[13]&IN2[34];
  assign P48[2] = IN1[13]&IN2[35];
  assign P49[1] = IN1[13]&IN2[36];
  assign P50[0] = IN1[13]&IN2[37];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[13] = IN1[14]&IN2[24];
  assign P39[12] = IN1[14]&IN2[25];
  assign P40[11] = IN1[14]&IN2[26];
  assign P41[10] = IN1[14]&IN2[27];
  assign P42[9] = IN1[14]&IN2[28];
  assign P43[8] = IN1[14]&IN2[29];
  assign P44[7] = IN1[14]&IN2[30];
  assign P45[6] = IN1[14]&IN2[31];
  assign P46[5] = IN1[14]&IN2[32];
  assign P47[4] = IN1[14]&IN2[33];
  assign P48[3] = IN1[14]&IN2[34];
  assign P49[2] = IN1[14]&IN2[35];
  assign P50[1] = IN1[14]&IN2[36];
  assign P51[0] = IN1[14]&IN2[37];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[14] = IN1[15]&IN2[23];
  assign P39[13] = IN1[15]&IN2[24];
  assign P40[12] = IN1[15]&IN2[25];
  assign P41[11] = IN1[15]&IN2[26];
  assign P42[10] = IN1[15]&IN2[27];
  assign P43[9] = IN1[15]&IN2[28];
  assign P44[8] = IN1[15]&IN2[29];
  assign P45[7] = IN1[15]&IN2[30];
  assign P46[6] = IN1[15]&IN2[31];
  assign P47[5] = IN1[15]&IN2[32];
  assign P48[4] = IN1[15]&IN2[33];
  assign P49[3] = IN1[15]&IN2[34];
  assign P50[2] = IN1[15]&IN2[35];
  assign P51[1] = IN1[15]&IN2[36];
  assign P52[0] = IN1[15]&IN2[37];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[15] = IN1[16]&IN2[22];
  assign P39[14] = IN1[16]&IN2[23];
  assign P40[13] = IN1[16]&IN2[24];
  assign P41[12] = IN1[16]&IN2[25];
  assign P42[11] = IN1[16]&IN2[26];
  assign P43[10] = IN1[16]&IN2[27];
  assign P44[9] = IN1[16]&IN2[28];
  assign P45[8] = IN1[16]&IN2[29];
  assign P46[7] = IN1[16]&IN2[30];
  assign P47[6] = IN1[16]&IN2[31];
  assign P48[5] = IN1[16]&IN2[32];
  assign P49[4] = IN1[16]&IN2[33];
  assign P50[3] = IN1[16]&IN2[34];
  assign P51[2] = IN1[16]&IN2[35];
  assign P52[1] = IN1[16]&IN2[36];
  assign P53[0] = IN1[16]&IN2[37];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[16] = IN1[17]&IN2[21];
  assign P39[15] = IN1[17]&IN2[22];
  assign P40[14] = IN1[17]&IN2[23];
  assign P41[13] = IN1[17]&IN2[24];
  assign P42[12] = IN1[17]&IN2[25];
  assign P43[11] = IN1[17]&IN2[26];
  assign P44[10] = IN1[17]&IN2[27];
  assign P45[9] = IN1[17]&IN2[28];
  assign P46[8] = IN1[17]&IN2[29];
  assign P47[7] = IN1[17]&IN2[30];
  assign P48[6] = IN1[17]&IN2[31];
  assign P49[5] = IN1[17]&IN2[32];
  assign P50[4] = IN1[17]&IN2[33];
  assign P51[3] = IN1[17]&IN2[34];
  assign P52[2] = IN1[17]&IN2[35];
  assign P53[1] = IN1[17]&IN2[36];
  assign P54[0] = IN1[17]&IN2[37];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[17] = IN1[18]&IN2[20];
  assign P39[16] = IN1[18]&IN2[21];
  assign P40[15] = IN1[18]&IN2[22];
  assign P41[14] = IN1[18]&IN2[23];
  assign P42[13] = IN1[18]&IN2[24];
  assign P43[12] = IN1[18]&IN2[25];
  assign P44[11] = IN1[18]&IN2[26];
  assign P45[10] = IN1[18]&IN2[27];
  assign P46[9] = IN1[18]&IN2[28];
  assign P47[8] = IN1[18]&IN2[29];
  assign P48[7] = IN1[18]&IN2[30];
  assign P49[6] = IN1[18]&IN2[31];
  assign P50[5] = IN1[18]&IN2[32];
  assign P51[4] = IN1[18]&IN2[33];
  assign P52[3] = IN1[18]&IN2[34];
  assign P53[2] = IN1[18]&IN2[35];
  assign P54[1] = IN1[18]&IN2[36];
  assign P55[0] = IN1[18]&IN2[37];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[18] = IN1[19]&IN2[19];
  assign P39[17] = IN1[19]&IN2[20];
  assign P40[16] = IN1[19]&IN2[21];
  assign P41[15] = IN1[19]&IN2[22];
  assign P42[14] = IN1[19]&IN2[23];
  assign P43[13] = IN1[19]&IN2[24];
  assign P44[12] = IN1[19]&IN2[25];
  assign P45[11] = IN1[19]&IN2[26];
  assign P46[10] = IN1[19]&IN2[27];
  assign P47[9] = IN1[19]&IN2[28];
  assign P48[8] = IN1[19]&IN2[29];
  assign P49[7] = IN1[19]&IN2[30];
  assign P50[6] = IN1[19]&IN2[31];
  assign P51[5] = IN1[19]&IN2[32];
  assign P52[4] = IN1[19]&IN2[33];
  assign P53[3] = IN1[19]&IN2[34];
  assign P54[2] = IN1[19]&IN2[35];
  assign P55[1] = IN1[19]&IN2[36];
  assign P56[0] = IN1[19]&IN2[37];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[19] = IN1[20]&IN2[18];
  assign P39[18] = IN1[20]&IN2[19];
  assign P40[17] = IN1[20]&IN2[20];
  assign P41[16] = IN1[20]&IN2[21];
  assign P42[15] = IN1[20]&IN2[22];
  assign P43[14] = IN1[20]&IN2[23];
  assign P44[13] = IN1[20]&IN2[24];
  assign P45[12] = IN1[20]&IN2[25];
  assign P46[11] = IN1[20]&IN2[26];
  assign P47[10] = IN1[20]&IN2[27];
  assign P48[9] = IN1[20]&IN2[28];
  assign P49[8] = IN1[20]&IN2[29];
  assign P50[7] = IN1[20]&IN2[30];
  assign P51[6] = IN1[20]&IN2[31];
  assign P52[5] = IN1[20]&IN2[32];
  assign P53[4] = IN1[20]&IN2[33];
  assign P54[3] = IN1[20]&IN2[34];
  assign P55[2] = IN1[20]&IN2[35];
  assign P56[1] = IN1[20]&IN2[36];
  assign P57[0] = IN1[20]&IN2[37];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[21] = IN1[21]&IN2[14];
  assign P36[21] = IN1[21]&IN2[15];
  assign P37[21] = IN1[21]&IN2[16];
  assign P38[20] = IN1[21]&IN2[17];
  assign P39[19] = IN1[21]&IN2[18];
  assign P40[18] = IN1[21]&IN2[19];
  assign P41[17] = IN1[21]&IN2[20];
  assign P42[16] = IN1[21]&IN2[21];
  assign P43[15] = IN1[21]&IN2[22];
  assign P44[14] = IN1[21]&IN2[23];
  assign P45[13] = IN1[21]&IN2[24];
  assign P46[12] = IN1[21]&IN2[25];
  assign P47[11] = IN1[21]&IN2[26];
  assign P48[10] = IN1[21]&IN2[27];
  assign P49[9] = IN1[21]&IN2[28];
  assign P50[8] = IN1[21]&IN2[29];
  assign P51[7] = IN1[21]&IN2[30];
  assign P52[6] = IN1[21]&IN2[31];
  assign P53[5] = IN1[21]&IN2[32];
  assign P54[4] = IN1[21]&IN2[33];
  assign P55[3] = IN1[21]&IN2[34];
  assign P56[2] = IN1[21]&IN2[35];
  assign P57[1] = IN1[21]&IN2[36];
  assign P58[0] = IN1[21]&IN2[37];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[22] = IN1[22]&IN2[13];
  assign P36[22] = IN1[22]&IN2[14];
  assign P37[22] = IN1[22]&IN2[15];
  assign P38[21] = IN1[22]&IN2[16];
  assign P39[20] = IN1[22]&IN2[17];
  assign P40[19] = IN1[22]&IN2[18];
  assign P41[18] = IN1[22]&IN2[19];
  assign P42[17] = IN1[22]&IN2[20];
  assign P43[16] = IN1[22]&IN2[21];
  assign P44[15] = IN1[22]&IN2[22];
  assign P45[14] = IN1[22]&IN2[23];
  assign P46[13] = IN1[22]&IN2[24];
  assign P47[12] = IN1[22]&IN2[25];
  assign P48[11] = IN1[22]&IN2[26];
  assign P49[10] = IN1[22]&IN2[27];
  assign P50[9] = IN1[22]&IN2[28];
  assign P51[8] = IN1[22]&IN2[29];
  assign P52[7] = IN1[22]&IN2[30];
  assign P53[6] = IN1[22]&IN2[31];
  assign P54[5] = IN1[22]&IN2[32];
  assign P55[4] = IN1[22]&IN2[33];
  assign P56[3] = IN1[22]&IN2[34];
  assign P57[2] = IN1[22]&IN2[35];
  assign P58[1] = IN1[22]&IN2[36];
  assign P59[0] = IN1[22]&IN2[37];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[23] = IN1[23]&IN2[12];
  assign P36[23] = IN1[23]&IN2[13];
  assign P37[23] = IN1[23]&IN2[14];
  assign P38[22] = IN1[23]&IN2[15];
  assign P39[21] = IN1[23]&IN2[16];
  assign P40[20] = IN1[23]&IN2[17];
  assign P41[19] = IN1[23]&IN2[18];
  assign P42[18] = IN1[23]&IN2[19];
  assign P43[17] = IN1[23]&IN2[20];
  assign P44[16] = IN1[23]&IN2[21];
  assign P45[15] = IN1[23]&IN2[22];
  assign P46[14] = IN1[23]&IN2[23];
  assign P47[13] = IN1[23]&IN2[24];
  assign P48[12] = IN1[23]&IN2[25];
  assign P49[11] = IN1[23]&IN2[26];
  assign P50[10] = IN1[23]&IN2[27];
  assign P51[9] = IN1[23]&IN2[28];
  assign P52[8] = IN1[23]&IN2[29];
  assign P53[7] = IN1[23]&IN2[30];
  assign P54[6] = IN1[23]&IN2[31];
  assign P55[5] = IN1[23]&IN2[32];
  assign P56[4] = IN1[23]&IN2[33];
  assign P57[3] = IN1[23]&IN2[34];
  assign P58[2] = IN1[23]&IN2[35];
  assign P59[1] = IN1[23]&IN2[36];
  assign P60[0] = IN1[23]&IN2[37];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[24] = IN1[24]&IN2[11];
  assign P36[24] = IN1[24]&IN2[12];
  assign P37[24] = IN1[24]&IN2[13];
  assign P38[23] = IN1[24]&IN2[14];
  assign P39[22] = IN1[24]&IN2[15];
  assign P40[21] = IN1[24]&IN2[16];
  assign P41[20] = IN1[24]&IN2[17];
  assign P42[19] = IN1[24]&IN2[18];
  assign P43[18] = IN1[24]&IN2[19];
  assign P44[17] = IN1[24]&IN2[20];
  assign P45[16] = IN1[24]&IN2[21];
  assign P46[15] = IN1[24]&IN2[22];
  assign P47[14] = IN1[24]&IN2[23];
  assign P48[13] = IN1[24]&IN2[24];
  assign P49[12] = IN1[24]&IN2[25];
  assign P50[11] = IN1[24]&IN2[26];
  assign P51[10] = IN1[24]&IN2[27];
  assign P52[9] = IN1[24]&IN2[28];
  assign P53[8] = IN1[24]&IN2[29];
  assign P54[7] = IN1[24]&IN2[30];
  assign P55[6] = IN1[24]&IN2[31];
  assign P56[5] = IN1[24]&IN2[32];
  assign P57[4] = IN1[24]&IN2[33];
  assign P58[3] = IN1[24]&IN2[34];
  assign P59[2] = IN1[24]&IN2[35];
  assign P60[1] = IN1[24]&IN2[36];
  assign P61[0] = IN1[24]&IN2[37];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[25] = IN1[25]&IN2[10];
  assign P36[25] = IN1[25]&IN2[11];
  assign P37[25] = IN1[25]&IN2[12];
  assign P38[24] = IN1[25]&IN2[13];
  assign P39[23] = IN1[25]&IN2[14];
  assign P40[22] = IN1[25]&IN2[15];
  assign P41[21] = IN1[25]&IN2[16];
  assign P42[20] = IN1[25]&IN2[17];
  assign P43[19] = IN1[25]&IN2[18];
  assign P44[18] = IN1[25]&IN2[19];
  assign P45[17] = IN1[25]&IN2[20];
  assign P46[16] = IN1[25]&IN2[21];
  assign P47[15] = IN1[25]&IN2[22];
  assign P48[14] = IN1[25]&IN2[23];
  assign P49[13] = IN1[25]&IN2[24];
  assign P50[12] = IN1[25]&IN2[25];
  assign P51[11] = IN1[25]&IN2[26];
  assign P52[10] = IN1[25]&IN2[27];
  assign P53[9] = IN1[25]&IN2[28];
  assign P54[8] = IN1[25]&IN2[29];
  assign P55[7] = IN1[25]&IN2[30];
  assign P56[6] = IN1[25]&IN2[31];
  assign P57[5] = IN1[25]&IN2[32];
  assign P58[4] = IN1[25]&IN2[33];
  assign P59[3] = IN1[25]&IN2[34];
  assign P60[2] = IN1[25]&IN2[35];
  assign P61[1] = IN1[25]&IN2[36];
  assign P62[0] = IN1[25]&IN2[37];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [25:0] IN26;
  input [25:0] IN27;
  input [25:0] IN28;
  input [25:0] IN29;
  input [25:0] IN30;
  input [25:0] IN31;
  input [25:0] IN32;
  input [25:0] IN33;
  input [25:0] IN34;
  input [25:0] IN35;
  input [25:0] IN36;
  input [25:0] IN37;
  input [24:0] IN38;
  input [23:0] IN39;
  input [22:0] IN40;
  input [21:0] IN41;
  input [20:0] IN42;
  input [19:0] IN43;
  input [18:0] IN44;
  input [17:0] IN45;
  input [16:0] IN46;
  input [15:0] IN47;
  input [14:0] IN48;
  input [13:0] IN49;
  input [12:0] IN50;
  input [11:0] IN51;
  input [10:0] IN52;
  input [9:0] IN53;
  input [8:0] IN54;
  input [7:0] IN55;
  input [6:0] IN56;
  input [5:0] IN57;
  input [4:0] IN58;
  input [3:0] IN59;
  input [2:0] IN60;
  input [1:0] IN61;
  input [0:0] IN62;
  output [62:0] Out1;
  output [36:0] Out2;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1984;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2050;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2139;
  wire w2140;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2585;
  wire w2586;
  wire w2587;
  wire w2589;
  wire w2590;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2614;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2631;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2680;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2685;
  wire w2686;
  wire w2687;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2694;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2708;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2747;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2770;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2774;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2785;
  wire w2786;
  wire w2787;
  wire w2789;
  wire w2791;
  wire w2793;
  wire w2795;
  wire w2797;
  wire w2799;
  wire w2801;
  wire w2803;
  wire w2805;
  wire w2807;
  wire w2809;
  wire w2811;
  wire w2813;
  wire w2815;
  wire w2817;
  wire w2819;
  wire w2821;
  wire w2823;
  wire w2825;
  wire w2827;
  wire w2829;
  wire w2831;
  wire w2833;
  wire w2835;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w989);
  FullAdder U1 (w989, IN2[0], IN2[1], w990, w991);
  FullAdder U2 (w991, IN3[0], IN3[1], w992, w993);
  FullAdder U3 (w993, IN4[0], IN4[1], w994, w995);
  FullAdder U4 (w995, IN5[0], IN5[1], w996, w997);
  FullAdder U5 (w997, IN6[0], IN6[1], w998, w999);
  FullAdder U6 (w999, IN7[0], IN7[1], w1000, w1001);
  FullAdder U7 (w1001, IN8[0], IN8[1], w1002, w1003);
  FullAdder U8 (w1003, IN9[0], IN9[1], w1004, w1005);
  FullAdder U9 (w1005, IN10[0], IN10[1], w1006, w1007);
  FullAdder U10 (w1007, IN11[0], IN11[1], w1008, w1009);
  FullAdder U11 (w1009, IN12[0], IN12[1], w1010, w1011);
  FullAdder U12 (w1011, IN13[0], IN13[1], w1012, w1013);
  FullAdder U13 (w1013, IN14[0], IN14[1], w1014, w1015);
  FullAdder U14 (w1015, IN15[0], IN15[1], w1016, w1017);
  FullAdder U15 (w1017, IN16[0], IN16[1], w1018, w1019);
  FullAdder U16 (w1019, IN17[0], IN17[1], w1020, w1021);
  FullAdder U17 (w1021, IN18[0], IN18[1], w1022, w1023);
  FullAdder U18 (w1023, IN19[0], IN19[1], w1024, w1025);
  FullAdder U19 (w1025, IN20[0], IN20[1], w1026, w1027);
  FullAdder U20 (w1027, IN21[0], IN21[1], w1028, w1029);
  FullAdder U21 (w1029, IN22[0], IN22[1], w1030, w1031);
  FullAdder U22 (w1031, IN23[0], IN23[1], w1032, w1033);
  FullAdder U23 (w1033, IN24[0], IN24[1], w1034, w1035);
  FullAdder U24 (w1035, IN25[0], IN25[1], w1036, w1037);
  HalfAdder U25 (w990, IN2[2], Out1[2], w1039);
  FullAdder U26 (w1039, w992, IN3[2], w1040, w1041);
  FullAdder U27 (w1041, w994, IN4[2], w1042, w1043);
  FullAdder U28 (w1043, w996, IN5[2], w1044, w1045);
  FullAdder U29 (w1045, w998, IN6[2], w1046, w1047);
  FullAdder U30 (w1047, w1000, IN7[2], w1048, w1049);
  FullAdder U31 (w1049, w1002, IN8[2], w1050, w1051);
  FullAdder U32 (w1051, w1004, IN9[2], w1052, w1053);
  FullAdder U33 (w1053, w1006, IN10[2], w1054, w1055);
  FullAdder U34 (w1055, w1008, IN11[2], w1056, w1057);
  FullAdder U35 (w1057, w1010, IN12[2], w1058, w1059);
  FullAdder U36 (w1059, w1012, IN13[2], w1060, w1061);
  FullAdder U37 (w1061, w1014, IN14[2], w1062, w1063);
  FullAdder U38 (w1063, w1016, IN15[2], w1064, w1065);
  FullAdder U39 (w1065, w1018, IN16[2], w1066, w1067);
  FullAdder U40 (w1067, w1020, IN17[2], w1068, w1069);
  FullAdder U41 (w1069, w1022, IN18[2], w1070, w1071);
  FullAdder U42 (w1071, w1024, IN19[2], w1072, w1073);
  FullAdder U43 (w1073, w1026, IN20[2], w1074, w1075);
  FullAdder U44 (w1075, w1028, IN21[2], w1076, w1077);
  FullAdder U45 (w1077, w1030, IN22[2], w1078, w1079);
  FullAdder U46 (w1079, w1032, IN23[2], w1080, w1081);
  FullAdder U47 (w1081, w1034, IN24[2], w1082, w1083);
  FullAdder U48 (w1083, w1036, IN25[2], w1084, w1085);
  FullAdder U49 (w1085, w1037, IN26[0], w1086, w1087);
  HalfAdder U50 (w1040, IN3[3], Out1[3], w1089);
  FullAdder U51 (w1089, w1042, IN4[3], w1090, w1091);
  FullAdder U52 (w1091, w1044, IN5[3], w1092, w1093);
  FullAdder U53 (w1093, w1046, IN6[3], w1094, w1095);
  FullAdder U54 (w1095, w1048, IN7[3], w1096, w1097);
  FullAdder U55 (w1097, w1050, IN8[3], w1098, w1099);
  FullAdder U56 (w1099, w1052, IN9[3], w1100, w1101);
  FullAdder U57 (w1101, w1054, IN10[3], w1102, w1103);
  FullAdder U58 (w1103, w1056, IN11[3], w1104, w1105);
  FullAdder U59 (w1105, w1058, IN12[3], w1106, w1107);
  FullAdder U60 (w1107, w1060, IN13[3], w1108, w1109);
  FullAdder U61 (w1109, w1062, IN14[3], w1110, w1111);
  FullAdder U62 (w1111, w1064, IN15[3], w1112, w1113);
  FullAdder U63 (w1113, w1066, IN16[3], w1114, w1115);
  FullAdder U64 (w1115, w1068, IN17[3], w1116, w1117);
  FullAdder U65 (w1117, w1070, IN18[3], w1118, w1119);
  FullAdder U66 (w1119, w1072, IN19[3], w1120, w1121);
  FullAdder U67 (w1121, w1074, IN20[3], w1122, w1123);
  FullAdder U68 (w1123, w1076, IN21[3], w1124, w1125);
  FullAdder U69 (w1125, w1078, IN22[3], w1126, w1127);
  FullAdder U70 (w1127, w1080, IN23[3], w1128, w1129);
  FullAdder U71 (w1129, w1082, IN24[3], w1130, w1131);
  FullAdder U72 (w1131, w1084, IN25[3], w1132, w1133);
  FullAdder U73 (w1133, w1086, IN26[1], w1134, w1135);
  FullAdder U74 (w1135, w1087, IN27[0], w1136, w1137);
  HalfAdder U75 (w1090, IN4[4], Out1[4], w1139);
  FullAdder U76 (w1139, w1092, IN5[4], w1140, w1141);
  FullAdder U77 (w1141, w1094, IN6[4], w1142, w1143);
  FullAdder U78 (w1143, w1096, IN7[4], w1144, w1145);
  FullAdder U79 (w1145, w1098, IN8[4], w1146, w1147);
  FullAdder U80 (w1147, w1100, IN9[4], w1148, w1149);
  FullAdder U81 (w1149, w1102, IN10[4], w1150, w1151);
  FullAdder U82 (w1151, w1104, IN11[4], w1152, w1153);
  FullAdder U83 (w1153, w1106, IN12[4], w1154, w1155);
  FullAdder U84 (w1155, w1108, IN13[4], w1156, w1157);
  FullAdder U85 (w1157, w1110, IN14[4], w1158, w1159);
  FullAdder U86 (w1159, w1112, IN15[4], w1160, w1161);
  FullAdder U87 (w1161, w1114, IN16[4], w1162, w1163);
  FullAdder U88 (w1163, w1116, IN17[4], w1164, w1165);
  FullAdder U89 (w1165, w1118, IN18[4], w1166, w1167);
  FullAdder U90 (w1167, w1120, IN19[4], w1168, w1169);
  FullAdder U91 (w1169, w1122, IN20[4], w1170, w1171);
  FullAdder U92 (w1171, w1124, IN21[4], w1172, w1173);
  FullAdder U93 (w1173, w1126, IN22[4], w1174, w1175);
  FullAdder U94 (w1175, w1128, IN23[4], w1176, w1177);
  FullAdder U95 (w1177, w1130, IN24[4], w1178, w1179);
  FullAdder U96 (w1179, w1132, IN25[4], w1180, w1181);
  FullAdder U97 (w1181, w1134, IN26[2], w1182, w1183);
  FullAdder U98 (w1183, w1136, IN27[1], w1184, w1185);
  FullAdder U99 (w1185, w1137, IN28[0], w1186, w1187);
  HalfAdder U100 (w1140, IN5[5], Out1[5], w1189);
  FullAdder U101 (w1189, w1142, IN6[5], w1190, w1191);
  FullAdder U102 (w1191, w1144, IN7[5], w1192, w1193);
  FullAdder U103 (w1193, w1146, IN8[5], w1194, w1195);
  FullAdder U104 (w1195, w1148, IN9[5], w1196, w1197);
  FullAdder U105 (w1197, w1150, IN10[5], w1198, w1199);
  FullAdder U106 (w1199, w1152, IN11[5], w1200, w1201);
  FullAdder U107 (w1201, w1154, IN12[5], w1202, w1203);
  FullAdder U108 (w1203, w1156, IN13[5], w1204, w1205);
  FullAdder U109 (w1205, w1158, IN14[5], w1206, w1207);
  FullAdder U110 (w1207, w1160, IN15[5], w1208, w1209);
  FullAdder U111 (w1209, w1162, IN16[5], w1210, w1211);
  FullAdder U112 (w1211, w1164, IN17[5], w1212, w1213);
  FullAdder U113 (w1213, w1166, IN18[5], w1214, w1215);
  FullAdder U114 (w1215, w1168, IN19[5], w1216, w1217);
  FullAdder U115 (w1217, w1170, IN20[5], w1218, w1219);
  FullAdder U116 (w1219, w1172, IN21[5], w1220, w1221);
  FullAdder U117 (w1221, w1174, IN22[5], w1222, w1223);
  FullAdder U118 (w1223, w1176, IN23[5], w1224, w1225);
  FullAdder U119 (w1225, w1178, IN24[5], w1226, w1227);
  FullAdder U120 (w1227, w1180, IN25[5], w1228, w1229);
  FullAdder U121 (w1229, w1182, IN26[3], w1230, w1231);
  FullAdder U122 (w1231, w1184, IN27[2], w1232, w1233);
  FullAdder U123 (w1233, w1186, IN28[1], w1234, w1235);
  FullAdder U124 (w1235, w1187, IN29[0], w1236, w1237);
  HalfAdder U125 (w1190, IN6[6], Out1[6], w1239);
  FullAdder U126 (w1239, w1192, IN7[6], w1240, w1241);
  FullAdder U127 (w1241, w1194, IN8[6], w1242, w1243);
  FullAdder U128 (w1243, w1196, IN9[6], w1244, w1245);
  FullAdder U129 (w1245, w1198, IN10[6], w1246, w1247);
  FullAdder U130 (w1247, w1200, IN11[6], w1248, w1249);
  FullAdder U131 (w1249, w1202, IN12[6], w1250, w1251);
  FullAdder U132 (w1251, w1204, IN13[6], w1252, w1253);
  FullAdder U133 (w1253, w1206, IN14[6], w1254, w1255);
  FullAdder U134 (w1255, w1208, IN15[6], w1256, w1257);
  FullAdder U135 (w1257, w1210, IN16[6], w1258, w1259);
  FullAdder U136 (w1259, w1212, IN17[6], w1260, w1261);
  FullAdder U137 (w1261, w1214, IN18[6], w1262, w1263);
  FullAdder U138 (w1263, w1216, IN19[6], w1264, w1265);
  FullAdder U139 (w1265, w1218, IN20[6], w1266, w1267);
  FullAdder U140 (w1267, w1220, IN21[6], w1268, w1269);
  FullAdder U141 (w1269, w1222, IN22[6], w1270, w1271);
  FullAdder U142 (w1271, w1224, IN23[6], w1272, w1273);
  FullAdder U143 (w1273, w1226, IN24[6], w1274, w1275);
  FullAdder U144 (w1275, w1228, IN25[6], w1276, w1277);
  FullAdder U145 (w1277, w1230, IN26[4], w1278, w1279);
  FullAdder U146 (w1279, w1232, IN27[3], w1280, w1281);
  FullAdder U147 (w1281, w1234, IN28[2], w1282, w1283);
  FullAdder U148 (w1283, w1236, IN29[1], w1284, w1285);
  FullAdder U149 (w1285, w1237, IN30[0], w1286, w1287);
  HalfAdder U150 (w1240, IN7[7], Out1[7], w1289);
  FullAdder U151 (w1289, w1242, IN8[7], w1290, w1291);
  FullAdder U152 (w1291, w1244, IN9[7], w1292, w1293);
  FullAdder U153 (w1293, w1246, IN10[7], w1294, w1295);
  FullAdder U154 (w1295, w1248, IN11[7], w1296, w1297);
  FullAdder U155 (w1297, w1250, IN12[7], w1298, w1299);
  FullAdder U156 (w1299, w1252, IN13[7], w1300, w1301);
  FullAdder U157 (w1301, w1254, IN14[7], w1302, w1303);
  FullAdder U158 (w1303, w1256, IN15[7], w1304, w1305);
  FullAdder U159 (w1305, w1258, IN16[7], w1306, w1307);
  FullAdder U160 (w1307, w1260, IN17[7], w1308, w1309);
  FullAdder U161 (w1309, w1262, IN18[7], w1310, w1311);
  FullAdder U162 (w1311, w1264, IN19[7], w1312, w1313);
  FullAdder U163 (w1313, w1266, IN20[7], w1314, w1315);
  FullAdder U164 (w1315, w1268, IN21[7], w1316, w1317);
  FullAdder U165 (w1317, w1270, IN22[7], w1318, w1319);
  FullAdder U166 (w1319, w1272, IN23[7], w1320, w1321);
  FullAdder U167 (w1321, w1274, IN24[7], w1322, w1323);
  FullAdder U168 (w1323, w1276, IN25[7], w1324, w1325);
  FullAdder U169 (w1325, w1278, IN26[5], w1326, w1327);
  FullAdder U170 (w1327, w1280, IN27[4], w1328, w1329);
  FullAdder U171 (w1329, w1282, IN28[3], w1330, w1331);
  FullAdder U172 (w1331, w1284, IN29[2], w1332, w1333);
  FullAdder U173 (w1333, w1286, IN30[1], w1334, w1335);
  FullAdder U174 (w1335, w1287, IN31[0], w1336, w1337);
  HalfAdder U175 (w1290, IN8[8], Out1[8], w1339);
  FullAdder U176 (w1339, w1292, IN9[8], w1340, w1341);
  FullAdder U177 (w1341, w1294, IN10[8], w1342, w1343);
  FullAdder U178 (w1343, w1296, IN11[8], w1344, w1345);
  FullAdder U179 (w1345, w1298, IN12[8], w1346, w1347);
  FullAdder U180 (w1347, w1300, IN13[8], w1348, w1349);
  FullAdder U181 (w1349, w1302, IN14[8], w1350, w1351);
  FullAdder U182 (w1351, w1304, IN15[8], w1352, w1353);
  FullAdder U183 (w1353, w1306, IN16[8], w1354, w1355);
  FullAdder U184 (w1355, w1308, IN17[8], w1356, w1357);
  FullAdder U185 (w1357, w1310, IN18[8], w1358, w1359);
  FullAdder U186 (w1359, w1312, IN19[8], w1360, w1361);
  FullAdder U187 (w1361, w1314, IN20[8], w1362, w1363);
  FullAdder U188 (w1363, w1316, IN21[8], w1364, w1365);
  FullAdder U189 (w1365, w1318, IN22[8], w1366, w1367);
  FullAdder U190 (w1367, w1320, IN23[8], w1368, w1369);
  FullAdder U191 (w1369, w1322, IN24[8], w1370, w1371);
  FullAdder U192 (w1371, w1324, IN25[8], w1372, w1373);
  FullAdder U193 (w1373, w1326, IN26[6], w1374, w1375);
  FullAdder U194 (w1375, w1328, IN27[5], w1376, w1377);
  FullAdder U195 (w1377, w1330, IN28[4], w1378, w1379);
  FullAdder U196 (w1379, w1332, IN29[3], w1380, w1381);
  FullAdder U197 (w1381, w1334, IN30[2], w1382, w1383);
  FullAdder U198 (w1383, w1336, IN31[1], w1384, w1385);
  FullAdder U199 (w1385, w1337, IN32[0], w1386, w1387);
  HalfAdder U200 (w1340, IN9[9], Out1[9], w1389);
  FullAdder U201 (w1389, w1342, IN10[9], w1390, w1391);
  FullAdder U202 (w1391, w1344, IN11[9], w1392, w1393);
  FullAdder U203 (w1393, w1346, IN12[9], w1394, w1395);
  FullAdder U204 (w1395, w1348, IN13[9], w1396, w1397);
  FullAdder U205 (w1397, w1350, IN14[9], w1398, w1399);
  FullAdder U206 (w1399, w1352, IN15[9], w1400, w1401);
  FullAdder U207 (w1401, w1354, IN16[9], w1402, w1403);
  FullAdder U208 (w1403, w1356, IN17[9], w1404, w1405);
  FullAdder U209 (w1405, w1358, IN18[9], w1406, w1407);
  FullAdder U210 (w1407, w1360, IN19[9], w1408, w1409);
  FullAdder U211 (w1409, w1362, IN20[9], w1410, w1411);
  FullAdder U212 (w1411, w1364, IN21[9], w1412, w1413);
  FullAdder U213 (w1413, w1366, IN22[9], w1414, w1415);
  FullAdder U214 (w1415, w1368, IN23[9], w1416, w1417);
  FullAdder U215 (w1417, w1370, IN24[9], w1418, w1419);
  FullAdder U216 (w1419, w1372, IN25[9], w1420, w1421);
  FullAdder U217 (w1421, w1374, IN26[7], w1422, w1423);
  FullAdder U218 (w1423, w1376, IN27[6], w1424, w1425);
  FullAdder U219 (w1425, w1378, IN28[5], w1426, w1427);
  FullAdder U220 (w1427, w1380, IN29[4], w1428, w1429);
  FullAdder U221 (w1429, w1382, IN30[3], w1430, w1431);
  FullAdder U222 (w1431, w1384, IN31[2], w1432, w1433);
  FullAdder U223 (w1433, w1386, IN32[1], w1434, w1435);
  FullAdder U224 (w1435, w1387, IN33[0], w1436, w1437);
  HalfAdder U225 (w1390, IN10[10], Out1[10], w1439);
  FullAdder U226 (w1439, w1392, IN11[10], w1440, w1441);
  FullAdder U227 (w1441, w1394, IN12[10], w1442, w1443);
  FullAdder U228 (w1443, w1396, IN13[10], w1444, w1445);
  FullAdder U229 (w1445, w1398, IN14[10], w1446, w1447);
  FullAdder U230 (w1447, w1400, IN15[10], w1448, w1449);
  FullAdder U231 (w1449, w1402, IN16[10], w1450, w1451);
  FullAdder U232 (w1451, w1404, IN17[10], w1452, w1453);
  FullAdder U233 (w1453, w1406, IN18[10], w1454, w1455);
  FullAdder U234 (w1455, w1408, IN19[10], w1456, w1457);
  FullAdder U235 (w1457, w1410, IN20[10], w1458, w1459);
  FullAdder U236 (w1459, w1412, IN21[10], w1460, w1461);
  FullAdder U237 (w1461, w1414, IN22[10], w1462, w1463);
  FullAdder U238 (w1463, w1416, IN23[10], w1464, w1465);
  FullAdder U239 (w1465, w1418, IN24[10], w1466, w1467);
  FullAdder U240 (w1467, w1420, IN25[10], w1468, w1469);
  FullAdder U241 (w1469, w1422, IN26[8], w1470, w1471);
  FullAdder U242 (w1471, w1424, IN27[7], w1472, w1473);
  FullAdder U243 (w1473, w1426, IN28[6], w1474, w1475);
  FullAdder U244 (w1475, w1428, IN29[5], w1476, w1477);
  FullAdder U245 (w1477, w1430, IN30[4], w1478, w1479);
  FullAdder U246 (w1479, w1432, IN31[3], w1480, w1481);
  FullAdder U247 (w1481, w1434, IN32[2], w1482, w1483);
  FullAdder U248 (w1483, w1436, IN33[1], w1484, w1485);
  FullAdder U249 (w1485, w1437, IN34[0], w1486, w1487);
  HalfAdder U250 (w1440, IN11[11], Out1[11], w1489);
  FullAdder U251 (w1489, w1442, IN12[11], w1490, w1491);
  FullAdder U252 (w1491, w1444, IN13[11], w1492, w1493);
  FullAdder U253 (w1493, w1446, IN14[11], w1494, w1495);
  FullAdder U254 (w1495, w1448, IN15[11], w1496, w1497);
  FullAdder U255 (w1497, w1450, IN16[11], w1498, w1499);
  FullAdder U256 (w1499, w1452, IN17[11], w1500, w1501);
  FullAdder U257 (w1501, w1454, IN18[11], w1502, w1503);
  FullAdder U258 (w1503, w1456, IN19[11], w1504, w1505);
  FullAdder U259 (w1505, w1458, IN20[11], w1506, w1507);
  FullAdder U260 (w1507, w1460, IN21[11], w1508, w1509);
  FullAdder U261 (w1509, w1462, IN22[11], w1510, w1511);
  FullAdder U262 (w1511, w1464, IN23[11], w1512, w1513);
  FullAdder U263 (w1513, w1466, IN24[11], w1514, w1515);
  FullAdder U264 (w1515, w1468, IN25[11], w1516, w1517);
  FullAdder U265 (w1517, w1470, IN26[9], w1518, w1519);
  FullAdder U266 (w1519, w1472, IN27[8], w1520, w1521);
  FullAdder U267 (w1521, w1474, IN28[7], w1522, w1523);
  FullAdder U268 (w1523, w1476, IN29[6], w1524, w1525);
  FullAdder U269 (w1525, w1478, IN30[5], w1526, w1527);
  FullAdder U270 (w1527, w1480, IN31[4], w1528, w1529);
  FullAdder U271 (w1529, w1482, IN32[3], w1530, w1531);
  FullAdder U272 (w1531, w1484, IN33[2], w1532, w1533);
  FullAdder U273 (w1533, w1486, IN34[1], w1534, w1535);
  FullAdder U274 (w1535, w1487, IN35[0], w1536, w1537);
  HalfAdder U275 (w1490, IN12[12], Out1[12], w1539);
  FullAdder U276 (w1539, w1492, IN13[12], w1540, w1541);
  FullAdder U277 (w1541, w1494, IN14[12], w1542, w1543);
  FullAdder U278 (w1543, w1496, IN15[12], w1544, w1545);
  FullAdder U279 (w1545, w1498, IN16[12], w1546, w1547);
  FullAdder U280 (w1547, w1500, IN17[12], w1548, w1549);
  FullAdder U281 (w1549, w1502, IN18[12], w1550, w1551);
  FullAdder U282 (w1551, w1504, IN19[12], w1552, w1553);
  FullAdder U283 (w1553, w1506, IN20[12], w1554, w1555);
  FullAdder U284 (w1555, w1508, IN21[12], w1556, w1557);
  FullAdder U285 (w1557, w1510, IN22[12], w1558, w1559);
  FullAdder U286 (w1559, w1512, IN23[12], w1560, w1561);
  FullAdder U287 (w1561, w1514, IN24[12], w1562, w1563);
  FullAdder U288 (w1563, w1516, IN25[12], w1564, w1565);
  FullAdder U289 (w1565, w1518, IN26[10], w1566, w1567);
  FullAdder U290 (w1567, w1520, IN27[9], w1568, w1569);
  FullAdder U291 (w1569, w1522, IN28[8], w1570, w1571);
  FullAdder U292 (w1571, w1524, IN29[7], w1572, w1573);
  FullAdder U293 (w1573, w1526, IN30[6], w1574, w1575);
  FullAdder U294 (w1575, w1528, IN31[5], w1576, w1577);
  FullAdder U295 (w1577, w1530, IN32[4], w1578, w1579);
  FullAdder U296 (w1579, w1532, IN33[3], w1580, w1581);
  FullAdder U297 (w1581, w1534, IN34[2], w1582, w1583);
  FullAdder U298 (w1583, w1536, IN35[1], w1584, w1585);
  FullAdder U299 (w1585, w1537, IN36[0], w1586, w1587);
  HalfAdder U300 (w1540, IN13[13], Out1[13], w1589);
  FullAdder U301 (w1589, w1542, IN14[13], w1590, w1591);
  FullAdder U302 (w1591, w1544, IN15[13], w1592, w1593);
  FullAdder U303 (w1593, w1546, IN16[13], w1594, w1595);
  FullAdder U304 (w1595, w1548, IN17[13], w1596, w1597);
  FullAdder U305 (w1597, w1550, IN18[13], w1598, w1599);
  FullAdder U306 (w1599, w1552, IN19[13], w1600, w1601);
  FullAdder U307 (w1601, w1554, IN20[13], w1602, w1603);
  FullAdder U308 (w1603, w1556, IN21[13], w1604, w1605);
  FullAdder U309 (w1605, w1558, IN22[13], w1606, w1607);
  FullAdder U310 (w1607, w1560, IN23[13], w1608, w1609);
  FullAdder U311 (w1609, w1562, IN24[13], w1610, w1611);
  FullAdder U312 (w1611, w1564, IN25[13], w1612, w1613);
  FullAdder U313 (w1613, w1566, IN26[11], w1614, w1615);
  FullAdder U314 (w1615, w1568, IN27[10], w1616, w1617);
  FullAdder U315 (w1617, w1570, IN28[9], w1618, w1619);
  FullAdder U316 (w1619, w1572, IN29[8], w1620, w1621);
  FullAdder U317 (w1621, w1574, IN30[7], w1622, w1623);
  FullAdder U318 (w1623, w1576, IN31[6], w1624, w1625);
  FullAdder U319 (w1625, w1578, IN32[5], w1626, w1627);
  FullAdder U320 (w1627, w1580, IN33[4], w1628, w1629);
  FullAdder U321 (w1629, w1582, IN34[3], w1630, w1631);
  FullAdder U322 (w1631, w1584, IN35[2], w1632, w1633);
  FullAdder U323 (w1633, w1586, IN36[1], w1634, w1635);
  FullAdder U324 (w1635, w1587, IN37[0], w1636, w1637);
  HalfAdder U325 (w1590, IN14[14], Out1[14], w1639);
  FullAdder U326 (w1639, w1592, IN15[14], w1640, w1641);
  FullAdder U327 (w1641, w1594, IN16[14], w1642, w1643);
  FullAdder U328 (w1643, w1596, IN17[14], w1644, w1645);
  FullAdder U329 (w1645, w1598, IN18[14], w1646, w1647);
  FullAdder U330 (w1647, w1600, IN19[14], w1648, w1649);
  FullAdder U331 (w1649, w1602, IN20[14], w1650, w1651);
  FullAdder U332 (w1651, w1604, IN21[14], w1652, w1653);
  FullAdder U333 (w1653, w1606, IN22[14], w1654, w1655);
  FullAdder U334 (w1655, w1608, IN23[14], w1656, w1657);
  FullAdder U335 (w1657, w1610, IN24[14], w1658, w1659);
  FullAdder U336 (w1659, w1612, IN25[14], w1660, w1661);
  FullAdder U337 (w1661, w1614, IN26[12], w1662, w1663);
  FullAdder U338 (w1663, w1616, IN27[11], w1664, w1665);
  FullAdder U339 (w1665, w1618, IN28[10], w1666, w1667);
  FullAdder U340 (w1667, w1620, IN29[9], w1668, w1669);
  FullAdder U341 (w1669, w1622, IN30[8], w1670, w1671);
  FullAdder U342 (w1671, w1624, IN31[7], w1672, w1673);
  FullAdder U343 (w1673, w1626, IN32[6], w1674, w1675);
  FullAdder U344 (w1675, w1628, IN33[5], w1676, w1677);
  FullAdder U345 (w1677, w1630, IN34[4], w1678, w1679);
  FullAdder U346 (w1679, w1632, IN35[3], w1680, w1681);
  FullAdder U347 (w1681, w1634, IN36[2], w1682, w1683);
  FullAdder U348 (w1683, w1636, IN37[1], w1684, w1685);
  FullAdder U349 (w1685, w1637, IN38[0], w1686, w1687);
  HalfAdder U350 (w1640, IN15[15], Out1[15], w1689);
  FullAdder U351 (w1689, w1642, IN16[15], w1690, w1691);
  FullAdder U352 (w1691, w1644, IN17[15], w1692, w1693);
  FullAdder U353 (w1693, w1646, IN18[15], w1694, w1695);
  FullAdder U354 (w1695, w1648, IN19[15], w1696, w1697);
  FullAdder U355 (w1697, w1650, IN20[15], w1698, w1699);
  FullAdder U356 (w1699, w1652, IN21[15], w1700, w1701);
  FullAdder U357 (w1701, w1654, IN22[15], w1702, w1703);
  FullAdder U358 (w1703, w1656, IN23[15], w1704, w1705);
  FullAdder U359 (w1705, w1658, IN24[15], w1706, w1707);
  FullAdder U360 (w1707, w1660, IN25[15], w1708, w1709);
  FullAdder U361 (w1709, w1662, IN26[13], w1710, w1711);
  FullAdder U362 (w1711, w1664, IN27[12], w1712, w1713);
  FullAdder U363 (w1713, w1666, IN28[11], w1714, w1715);
  FullAdder U364 (w1715, w1668, IN29[10], w1716, w1717);
  FullAdder U365 (w1717, w1670, IN30[9], w1718, w1719);
  FullAdder U366 (w1719, w1672, IN31[8], w1720, w1721);
  FullAdder U367 (w1721, w1674, IN32[7], w1722, w1723);
  FullAdder U368 (w1723, w1676, IN33[6], w1724, w1725);
  FullAdder U369 (w1725, w1678, IN34[5], w1726, w1727);
  FullAdder U370 (w1727, w1680, IN35[4], w1728, w1729);
  FullAdder U371 (w1729, w1682, IN36[3], w1730, w1731);
  FullAdder U372 (w1731, w1684, IN37[2], w1732, w1733);
  FullAdder U373 (w1733, w1686, IN38[1], w1734, w1735);
  FullAdder U374 (w1735, w1687, IN39[0], w1736, w1737);
  HalfAdder U375 (w1690, IN16[16], Out1[16], w1739);
  FullAdder U376 (w1739, w1692, IN17[16], w1740, w1741);
  FullAdder U377 (w1741, w1694, IN18[16], w1742, w1743);
  FullAdder U378 (w1743, w1696, IN19[16], w1744, w1745);
  FullAdder U379 (w1745, w1698, IN20[16], w1746, w1747);
  FullAdder U380 (w1747, w1700, IN21[16], w1748, w1749);
  FullAdder U381 (w1749, w1702, IN22[16], w1750, w1751);
  FullAdder U382 (w1751, w1704, IN23[16], w1752, w1753);
  FullAdder U383 (w1753, w1706, IN24[16], w1754, w1755);
  FullAdder U384 (w1755, w1708, IN25[16], w1756, w1757);
  FullAdder U385 (w1757, w1710, IN26[14], w1758, w1759);
  FullAdder U386 (w1759, w1712, IN27[13], w1760, w1761);
  FullAdder U387 (w1761, w1714, IN28[12], w1762, w1763);
  FullAdder U388 (w1763, w1716, IN29[11], w1764, w1765);
  FullAdder U389 (w1765, w1718, IN30[10], w1766, w1767);
  FullAdder U390 (w1767, w1720, IN31[9], w1768, w1769);
  FullAdder U391 (w1769, w1722, IN32[8], w1770, w1771);
  FullAdder U392 (w1771, w1724, IN33[7], w1772, w1773);
  FullAdder U393 (w1773, w1726, IN34[6], w1774, w1775);
  FullAdder U394 (w1775, w1728, IN35[5], w1776, w1777);
  FullAdder U395 (w1777, w1730, IN36[4], w1778, w1779);
  FullAdder U396 (w1779, w1732, IN37[3], w1780, w1781);
  FullAdder U397 (w1781, w1734, IN38[2], w1782, w1783);
  FullAdder U398 (w1783, w1736, IN39[1], w1784, w1785);
  FullAdder U399 (w1785, w1737, IN40[0], w1786, w1787);
  HalfAdder U400 (w1740, IN17[17], Out1[17], w1789);
  FullAdder U401 (w1789, w1742, IN18[17], w1790, w1791);
  FullAdder U402 (w1791, w1744, IN19[17], w1792, w1793);
  FullAdder U403 (w1793, w1746, IN20[17], w1794, w1795);
  FullAdder U404 (w1795, w1748, IN21[17], w1796, w1797);
  FullAdder U405 (w1797, w1750, IN22[17], w1798, w1799);
  FullAdder U406 (w1799, w1752, IN23[17], w1800, w1801);
  FullAdder U407 (w1801, w1754, IN24[17], w1802, w1803);
  FullAdder U408 (w1803, w1756, IN25[17], w1804, w1805);
  FullAdder U409 (w1805, w1758, IN26[15], w1806, w1807);
  FullAdder U410 (w1807, w1760, IN27[14], w1808, w1809);
  FullAdder U411 (w1809, w1762, IN28[13], w1810, w1811);
  FullAdder U412 (w1811, w1764, IN29[12], w1812, w1813);
  FullAdder U413 (w1813, w1766, IN30[11], w1814, w1815);
  FullAdder U414 (w1815, w1768, IN31[10], w1816, w1817);
  FullAdder U415 (w1817, w1770, IN32[9], w1818, w1819);
  FullAdder U416 (w1819, w1772, IN33[8], w1820, w1821);
  FullAdder U417 (w1821, w1774, IN34[7], w1822, w1823);
  FullAdder U418 (w1823, w1776, IN35[6], w1824, w1825);
  FullAdder U419 (w1825, w1778, IN36[5], w1826, w1827);
  FullAdder U420 (w1827, w1780, IN37[4], w1828, w1829);
  FullAdder U421 (w1829, w1782, IN38[3], w1830, w1831);
  FullAdder U422 (w1831, w1784, IN39[2], w1832, w1833);
  FullAdder U423 (w1833, w1786, IN40[1], w1834, w1835);
  FullAdder U424 (w1835, w1787, IN41[0], w1836, w1837);
  HalfAdder U425 (w1790, IN18[18], Out1[18], w1839);
  FullAdder U426 (w1839, w1792, IN19[18], w1840, w1841);
  FullAdder U427 (w1841, w1794, IN20[18], w1842, w1843);
  FullAdder U428 (w1843, w1796, IN21[18], w1844, w1845);
  FullAdder U429 (w1845, w1798, IN22[18], w1846, w1847);
  FullAdder U430 (w1847, w1800, IN23[18], w1848, w1849);
  FullAdder U431 (w1849, w1802, IN24[18], w1850, w1851);
  FullAdder U432 (w1851, w1804, IN25[18], w1852, w1853);
  FullAdder U433 (w1853, w1806, IN26[16], w1854, w1855);
  FullAdder U434 (w1855, w1808, IN27[15], w1856, w1857);
  FullAdder U435 (w1857, w1810, IN28[14], w1858, w1859);
  FullAdder U436 (w1859, w1812, IN29[13], w1860, w1861);
  FullAdder U437 (w1861, w1814, IN30[12], w1862, w1863);
  FullAdder U438 (w1863, w1816, IN31[11], w1864, w1865);
  FullAdder U439 (w1865, w1818, IN32[10], w1866, w1867);
  FullAdder U440 (w1867, w1820, IN33[9], w1868, w1869);
  FullAdder U441 (w1869, w1822, IN34[8], w1870, w1871);
  FullAdder U442 (w1871, w1824, IN35[7], w1872, w1873);
  FullAdder U443 (w1873, w1826, IN36[6], w1874, w1875);
  FullAdder U444 (w1875, w1828, IN37[5], w1876, w1877);
  FullAdder U445 (w1877, w1830, IN38[4], w1878, w1879);
  FullAdder U446 (w1879, w1832, IN39[3], w1880, w1881);
  FullAdder U447 (w1881, w1834, IN40[2], w1882, w1883);
  FullAdder U448 (w1883, w1836, IN41[1], w1884, w1885);
  FullAdder U449 (w1885, w1837, IN42[0], w1886, w1887);
  HalfAdder U450 (w1840, IN19[19], Out1[19], w1889);
  FullAdder U451 (w1889, w1842, IN20[19], w1890, w1891);
  FullAdder U452 (w1891, w1844, IN21[19], w1892, w1893);
  FullAdder U453 (w1893, w1846, IN22[19], w1894, w1895);
  FullAdder U454 (w1895, w1848, IN23[19], w1896, w1897);
  FullAdder U455 (w1897, w1850, IN24[19], w1898, w1899);
  FullAdder U456 (w1899, w1852, IN25[19], w1900, w1901);
  FullAdder U457 (w1901, w1854, IN26[17], w1902, w1903);
  FullAdder U458 (w1903, w1856, IN27[16], w1904, w1905);
  FullAdder U459 (w1905, w1858, IN28[15], w1906, w1907);
  FullAdder U460 (w1907, w1860, IN29[14], w1908, w1909);
  FullAdder U461 (w1909, w1862, IN30[13], w1910, w1911);
  FullAdder U462 (w1911, w1864, IN31[12], w1912, w1913);
  FullAdder U463 (w1913, w1866, IN32[11], w1914, w1915);
  FullAdder U464 (w1915, w1868, IN33[10], w1916, w1917);
  FullAdder U465 (w1917, w1870, IN34[9], w1918, w1919);
  FullAdder U466 (w1919, w1872, IN35[8], w1920, w1921);
  FullAdder U467 (w1921, w1874, IN36[7], w1922, w1923);
  FullAdder U468 (w1923, w1876, IN37[6], w1924, w1925);
  FullAdder U469 (w1925, w1878, IN38[5], w1926, w1927);
  FullAdder U470 (w1927, w1880, IN39[4], w1928, w1929);
  FullAdder U471 (w1929, w1882, IN40[3], w1930, w1931);
  FullAdder U472 (w1931, w1884, IN41[2], w1932, w1933);
  FullAdder U473 (w1933, w1886, IN42[1], w1934, w1935);
  FullAdder U474 (w1935, w1887, IN43[0], w1936, w1937);
  HalfAdder U475 (w1890, IN20[20], Out1[20], w1939);
  FullAdder U476 (w1939, w1892, IN21[20], w1940, w1941);
  FullAdder U477 (w1941, w1894, IN22[20], w1942, w1943);
  FullAdder U478 (w1943, w1896, IN23[20], w1944, w1945);
  FullAdder U479 (w1945, w1898, IN24[20], w1946, w1947);
  FullAdder U480 (w1947, w1900, IN25[20], w1948, w1949);
  FullAdder U481 (w1949, w1902, IN26[18], w1950, w1951);
  FullAdder U482 (w1951, w1904, IN27[17], w1952, w1953);
  FullAdder U483 (w1953, w1906, IN28[16], w1954, w1955);
  FullAdder U484 (w1955, w1908, IN29[15], w1956, w1957);
  FullAdder U485 (w1957, w1910, IN30[14], w1958, w1959);
  FullAdder U486 (w1959, w1912, IN31[13], w1960, w1961);
  FullAdder U487 (w1961, w1914, IN32[12], w1962, w1963);
  FullAdder U488 (w1963, w1916, IN33[11], w1964, w1965);
  FullAdder U489 (w1965, w1918, IN34[10], w1966, w1967);
  FullAdder U490 (w1967, w1920, IN35[9], w1968, w1969);
  FullAdder U491 (w1969, w1922, IN36[8], w1970, w1971);
  FullAdder U492 (w1971, w1924, IN37[7], w1972, w1973);
  FullAdder U493 (w1973, w1926, IN38[6], w1974, w1975);
  FullAdder U494 (w1975, w1928, IN39[5], w1976, w1977);
  FullAdder U495 (w1977, w1930, IN40[4], w1978, w1979);
  FullAdder U496 (w1979, w1932, IN41[3], w1980, w1981);
  FullAdder U497 (w1981, w1934, IN42[2], w1982, w1983);
  FullAdder U498 (w1983, w1936, IN43[1], w1984, w1985);
  FullAdder U499 (w1985, w1937, IN44[0], w1986, w1987);
  HalfAdder U500 (w1940, IN21[21], Out1[21], w1989);
  FullAdder U501 (w1989, w1942, IN22[21], w1990, w1991);
  FullAdder U502 (w1991, w1944, IN23[21], w1992, w1993);
  FullAdder U503 (w1993, w1946, IN24[21], w1994, w1995);
  FullAdder U504 (w1995, w1948, IN25[21], w1996, w1997);
  FullAdder U505 (w1997, w1950, IN26[19], w1998, w1999);
  FullAdder U506 (w1999, w1952, IN27[18], w2000, w2001);
  FullAdder U507 (w2001, w1954, IN28[17], w2002, w2003);
  FullAdder U508 (w2003, w1956, IN29[16], w2004, w2005);
  FullAdder U509 (w2005, w1958, IN30[15], w2006, w2007);
  FullAdder U510 (w2007, w1960, IN31[14], w2008, w2009);
  FullAdder U511 (w2009, w1962, IN32[13], w2010, w2011);
  FullAdder U512 (w2011, w1964, IN33[12], w2012, w2013);
  FullAdder U513 (w2013, w1966, IN34[11], w2014, w2015);
  FullAdder U514 (w2015, w1968, IN35[10], w2016, w2017);
  FullAdder U515 (w2017, w1970, IN36[9], w2018, w2019);
  FullAdder U516 (w2019, w1972, IN37[8], w2020, w2021);
  FullAdder U517 (w2021, w1974, IN38[7], w2022, w2023);
  FullAdder U518 (w2023, w1976, IN39[6], w2024, w2025);
  FullAdder U519 (w2025, w1978, IN40[5], w2026, w2027);
  FullAdder U520 (w2027, w1980, IN41[4], w2028, w2029);
  FullAdder U521 (w2029, w1982, IN42[3], w2030, w2031);
  FullAdder U522 (w2031, w1984, IN43[2], w2032, w2033);
  FullAdder U523 (w2033, w1986, IN44[1], w2034, w2035);
  FullAdder U524 (w2035, w1987, IN45[0], w2036, w2037);
  HalfAdder U525 (w1990, IN22[22], Out1[22], w2039);
  FullAdder U526 (w2039, w1992, IN23[22], w2040, w2041);
  FullAdder U527 (w2041, w1994, IN24[22], w2042, w2043);
  FullAdder U528 (w2043, w1996, IN25[22], w2044, w2045);
  FullAdder U529 (w2045, w1998, IN26[20], w2046, w2047);
  FullAdder U530 (w2047, w2000, IN27[19], w2048, w2049);
  FullAdder U531 (w2049, w2002, IN28[18], w2050, w2051);
  FullAdder U532 (w2051, w2004, IN29[17], w2052, w2053);
  FullAdder U533 (w2053, w2006, IN30[16], w2054, w2055);
  FullAdder U534 (w2055, w2008, IN31[15], w2056, w2057);
  FullAdder U535 (w2057, w2010, IN32[14], w2058, w2059);
  FullAdder U536 (w2059, w2012, IN33[13], w2060, w2061);
  FullAdder U537 (w2061, w2014, IN34[12], w2062, w2063);
  FullAdder U538 (w2063, w2016, IN35[11], w2064, w2065);
  FullAdder U539 (w2065, w2018, IN36[10], w2066, w2067);
  FullAdder U540 (w2067, w2020, IN37[9], w2068, w2069);
  FullAdder U541 (w2069, w2022, IN38[8], w2070, w2071);
  FullAdder U542 (w2071, w2024, IN39[7], w2072, w2073);
  FullAdder U543 (w2073, w2026, IN40[6], w2074, w2075);
  FullAdder U544 (w2075, w2028, IN41[5], w2076, w2077);
  FullAdder U545 (w2077, w2030, IN42[4], w2078, w2079);
  FullAdder U546 (w2079, w2032, IN43[3], w2080, w2081);
  FullAdder U547 (w2081, w2034, IN44[2], w2082, w2083);
  FullAdder U548 (w2083, w2036, IN45[1], w2084, w2085);
  FullAdder U549 (w2085, w2037, IN46[0], w2086, w2087);
  HalfAdder U550 (w2040, IN23[23], Out1[23], w2089);
  FullAdder U551 (w2089, w2042, IN24[23], w2090, w2091);
  FullAdder U552 (w2091, w2044, IN25[23], w2092, w2093);
  FullAdder U553 (w2093, w2046, IN26[21], w2094, w2095);
  FullAdder U554 (w2095, w2048, IN27[20], w2096, w2097);
  FullAdder U555 (w2097, w2050, IN28[19], w2098, w2099);
  FullAdder U556 (w2099, w2052, IN29[18], w2100, w2101);
  FullAdder U557 (w2101, w2054, IN30[17], w2102, w2103);
  FullAdder U558 (w2103, w2056, IN31[16], w2104, w2105);
  FullAdder U559 (w2105, w2058, IN32[15], w2106, w2107);
  FullAdder U560 (w2107, w2060, IN33[14], w2108, w2109);
  FullAdder U561 (w2109, w2062, IN34[13], w2110, w2111);
  FullAdder U562 (w2111, w2064, IN35[12], w2112, w2113);
  FullAdder U563 (w2113, w2066, IN36[11], w2114, w2115);
  FullAdder U564 (w2115, w2068, IN37[10], w2116, w2117);
  FullAdder U565 (w2117, w2070, IN38[9], w2118, w2119);
  FullAdder U566 (w2119, w2072, IN39[8], w2120, w2121);
  FullAdder U567 (w2121, w2074, IN40[7], w2122, w2123);
  FullAdder U568 (w2123, w2076, IN41[6], w2124, w2125);
  FullAdder U569 (w2125, w2078, IN42[5], w2126, w2127);
  FullAdder U570 (w2127, w2080, IN43[4], w2128, w2129);
  FullAdder U571 (w2129, w2082, IN44[3], w2130, w2131);
  FullAdder U572 (w2131, w2084, IN45[2], w2132, w2133);
  FullAdder U573 (w2133, w2086, IN46[1], w2134, w2135);
  FullAdder U574 (w2135, w2087, IN47[0], w2136, w2137);
  HalfAdder U575 (w2090, IN24[24], Out1[24], w2139);
  FullAdder U576 (w2139, w2092, IN25[24], w2140, w2141);
  FullAdder U577 (w2141, w2094, IN26[22], w2142, w2143);
  FullAdder U578 (w2143, w2096, IN27[21], w2144, w2145);
  FullAdder U579 (w2145, w2098, IN28[20], w2146, w2147);
  FullAdder U580 (w2147, w2100, IN29[19], w2148, w2149);
  FullAdder U581 (w2149, w2102, IN30[18], w2150, w2151);
  FullAdder U582 (w2151, w2104, IN31[17], w2152, w2153);
  FullAdder U583 (w2153, w2106, IN32[16], w2154, w2155);
  FullAdder U584 (w2155, w2108, IN33[15], w2156, w2157);
  FullAdder U585 (w2157, w2110, IN34[14], w2158, w2159);
  FullAdder U586 (w2159, w2112, IN35[13], w2160, w2161);
  FullAdder U587 (w2161, w2114, IN36[12], w2162, w2163);
  FullAdder U588 (w2163, w2116, IN37[11], w2164, w2165);
  FullAdder U589 (w2165, w2118, IN38[10], w2166, w2167);
  FullAdder U590 (w2167, w2120, IN39[9], w2168, w2169);
  FullAdder U591 (w2169, w2122, IN40[8], w2170, w2171);
  FullAdder U592 (w2171, w2124, IN41[7], w2172, w2173);
  FullAdder U593 (w2173, w2126, IN42[6], w2174, w2175);
  FullAdder U594 (w2175, w2128, IN43[5], w2176, w2177);
  FullAdder U595 (w2177, w2130, IN44[4], w2178, w2179);
  FullAdder U596 (w2179, w2132, IN45[3], w2180, w2181);
  FullAdder U597 (w2181, w2134, IN46[2], w2182, w2183);
  FullAdder U598 (w2183, w2136, IN47[1], w2184, w2185);
  FullAdder U599 (w2185, w2137, IN48[0], w2186, w2187);
  HalfAdder U600 (w2140, IN25[25], Out1[25], w2189);
  FullAdder U601 (w2189, w2142, IN26[23], w2190, w2191);
  FullAdder U602 (w2191, w2144, IN27[22], w2192, w2193);
  FullAdder U603 (w2193, w2146, IN28[21], w2194, w2195);
  FullAdder U604 (w2195, w2148, IN29[20], w2196, w2197);
  FullAdder U605 (w2197, w2150, IN30[19], w2198, w2199);
  FullAdder U606 (w2199, w2152, IN31[18], w2200, w2201);
  FullAdder U607 (w2201, w2154, IN32[17], w2202, w2203);
  FullAdder U608 (w2203, w2156, IN33[16], w2204, w2205);
  FullAdder U609 (w2205, w2158, IN34[15], w2206, w2207);
  FullAdder U610 (w2207, w2160, IN35[14], w2208, w2209);
  FullAdder U611 (w2209, w2162, IN36[13], w2210, w2211);
  FullAdder U612 (w2211, w2164, IN37[12], w2212, w2213);
  FullAdder U613 (w2213, w2166, IN38[11], w2214, w2215);
  FullAdder U614 (w2215, w2168, IN39[10], w2216, w2217);
  FullAdder U615 (w2217, w2170, IN40[9], w2218, w2219);
  FullAdder U616 (w2219, w2172, IN41[8], w2220, w2221);
  FullAdder U617 (w2221, w2174, IN42[7], w2222, w2223);
  FullAdder U618 (w2223, w2176, IN43[6], w2224, w2225);
  FullAdder U619 (w2225, w2178, IN44[5], w2226, w2227);
  FullAdder U620 (w2227, w2180, IN45[4], w2228, w2229);
  FullAdder U621 (w2229, w2182, IN46[3], w2230, w2231);
  FullAdder U622 (w2231, w2184, IN47[2], w2232, w2233);
  FullAdder U623 (w2233, w2186, IN48[1], w2234, w2235);
  FullAdder U624 (w2235, w2187, IN49[0], w2236, w2237);
  HalfAdder U625 (w2190, IN26[24], Out1[26], w2239);
  FullAdder U626 (w2239, w2192, IN27[23], w2240, w2241);
  FullAdder U627 (w2241, w2194, IN28[22], w2242, w2243);
  FullAdder U628 (w2243, w2196, IN29[21], w2244, w2245);
  FullAdder U629 (w2245, w2198, IN30[20], w2246, w2247);
  FullAdder U630 (w2247, w2200, IN31[19], w2248, w2249);
  FullAdder U631 (w2249, w2202, IN32[18], w2250, w2251);
  FullAdder U632 (w2251, w2204, IN33[17], w2252, w2253);
  FullAdder U633 (w2253, w2206, IN34[16], w2254, w2255);
  FullAdder U634 (w2255, w2208, IN35[15], w2256, w2257);
  FullAdder U635 (w2257, w2210, IN36[14], w2258, w2259);
  FullAdder U636 (w2259, w2212, IN37[13], w2260, w2261);
  FullAdder U637 (w2261, w2214, IN38[12], w2262, w2263);
  FullAdder U638 (w2263, w2216, IN39[11], w2264, w2265);
  FullAdder U639 (w2265, w2218, IN40[10], w2266, w2267);
  FullAdder U640 (w2267, w2220, IN41[9], w2268, w2269);
  FullAdder U641 (w2269, w2222, IN42[8], w2270, w2271);
  FullAdder U642 (w2271, w2224, IN43[7], w2272, w2273);
  FullAdder U643 (w2273, w2226, IN44[6], w2274, w2275);
  FullAdder U644 (w2275, w2228, IN45[5], w2276, w2277);
  FullAdder U645 (w2277, w2230, IN46[4], w2278, w2279);
  FullAdder U646 (w2279, w2232, IN47[3], w2280, w2281);
  FullAdder U647 (w2281, w2234, IN48[2], w2282, w2283);
  FullAdder U648 (w2283, w2236, IN49[1], w2284, w2285);
  FullAdder U649 (w2285, w2237, IN50[0], w2286, w2287);
  HalfAdder U650 (w2240, IN27[24], Out1[27], w2289);
  FullAdder U651 (w2289, w2242, IN28[23], w2290, w2291);
  FullAdder U652 (w2291, w2244, IN29[22], w2292, w2293);
  FullAdder U653 (w2293, w2246, IN30[21], w2294, w2295);
  FullAdder U654 (w2295, w2248, IN31[20], w2296, w2297);
  FullAdder U655 (w2297, w2250, IN32[19], w2298, w2299);
  FullAdder U656 (w2299, w2252, IN33[18], w2300, w2301);
  FullAdder U657 (w2301, w2254, IN34[17], w2302, w2303);
  FullAdder U658 (w2303, w2256, IN35[16], w2304, w2305);
  FullAdder U659 (w2305, w2258, IN36[15], w2306, w2307);
  FullAdder U660 (w2307, w2260, IN37[14], w2308, w2309);
  FullAdder U661 (w2309, w2262, IN38[13], w2310, w2311);
  FullAdder U662 (w2311, w2264, IN39[12], w2312, w2313);
  FullAdder U663 (w2313, w2266, IN40[11], w2314, w2315);
  FullAdder U664 (w2315, w2268, IN41[10], w2316, w2317);
  FullAdder U665 (w2317, w2270, IN42[9], w2318, w2319);
  FullAdder U666 (w2319, w2272, IN43[8], w2320, w2321);
  FullAdder U667 (w2321, w2274, IN44[7], w2322, w2323);
  FullAdder U668 (w2323, w2276, IN45[6], w2324, w2325);
  FullAdder U669 (w2325, w2278, IN46[5], w2326, w2327);
  FullAdder U670 (w2327, w2280, IN47[4], w2328, w2329);
  FullAdder U671 (w2329, w2282, IN48[3], w2330, w2331);
  FullAdder U672 (w2331, w2284, IN49[2], w2332, w2333);
  FullAdder U673 (w2333, w2286, IN50[1], w2334, w2335);
  FullAdder U674 (w2335, w2287, IN51[0], w2336, w2337);
  HalfAdder U675 (w2290, IN28[24], Out1[28], w2339);
  FullAdder U676 (w2339, w2292, IN29[23], w2340, w2341);
  FullAdder U677 (w2341, w2294, IN30[22], w2342, w2343);
  FullAdder U678 (w2343, w2296, IN31[21], w2344, w2345);
  FullAdder U679 (w2345, w2298, IN32[20], w2346, w2347);
  FullAdder U680 (w2347, w2300, IN33[19], w2348, w2349);
  FullAdder U681 (w2349, w2302, IN34[18], w2350, w2351);
  FullAdder U682 (w2351, w2304, IN35[17], w2352, w2353);
  FullAdder U683 (w2353, w2306, IN36[16], w2354, w2355);
  FullAdder U684 (w2355, w2308, IN37[15], w2356, w2357);
  FullAdder U685 (w2357, w2310, IN38[14], w2358, w2359);
  FullAdder U686 (w2359, w2312, IN39[13], w2360, w2361);
  FullAdder U687 (w2361, w2314, IN40[12], w2362, w2363);
  FullAdder U688 (w2363, w2316, IN41[11], w2364, w2365);
  FullAdder U689 (w2365, w2318, IN42[10], w2366, w2367);
  FullAdder U690 (w2367, w2320, IN43[9], w2368, w2369);
  FullAdder U691 (w2369, w2322, IN44[8], w2370, w2371);
  FullAdder U692 (w2371, w2324, IN45[7], w2372, w2373);
  FullAdder U693 (w2373, w2326, IN46[6], w2374, w2375);
  FullAdder U694 (w2375, w2328, IN47[5], w2376, w2377);
  FullAdder U695 (w2377, w2330, IN48[4], w2378, w2379);
  FullAdder U696 (w2379, w2332, IN49[3], w2380, w2381);
  FullAdder U697 (w2381, w2334, IN50[2], w2382, w2383);
  FullAdder U698 (w2383, w2336, IN51[1], w2384, w2385);
  FullAdder U699 (w2385, w2337, IN52[0], w2386, w2387);
  HalfAdder U700 (w2340, IN29[24], Out1[29], w2389);
  FullAdder U701 (w2389, w2342, IN30[23], w2390, w2391);
  FullAdder U702 (w2391, w2344, IN31[22], w2392, w2393);
  FullAdder U703 (w2393, w2346, IN32[21], w2394, w2395);
  FullAdder U704 (w2395, w2348, IN33[20], w2396, w2397);
  FullAdder U705 (w2397, w2350, IN34[19], w2398, w2399);
  FullAdder U706 (w2399, w2352, IN35[18], w2400, w2401);
  FullAdder U707 (w2401, w2354, IN36[17], w2402, w2403);
  FullAdder U708 (w2403, w2356, IN37[16], w2404, w2405);
  FullAdder U709 (w2405, w2358, IN38[15], w2406, w2407);
  FullAdder U710 (w2407, w2360, IN39[14], w2408, w2409);
  FullAdder U711 (w2409, w2362, IN40[13], w2410, w2411);
  FullAdder U712 (w2411, w2364, IN41[12], w2412, w2413);
  FullAdder U713 (w2413, w2366, IN42[11], w2414, w2415);
  FullAdder U714 (w2415, w2368, IN43[10], w2416, w2417);
  FullAdder U715 (w2417, w2370, IN44[9], w2418, w2419);
  FullAdder U716 (w2419, w2372, IN45[8], w2420, w2421);
  FullAdder U717 (w2421, w2374, IN46[7], w2422, w2423);
  FullAdder U718 (w2423, w2376, IN47[6], w2424, w2425);
  FullAdder U719 (w2425, w2378, IN48[5], w2426, w2427);
  FullAdder U720 (w2427, w2380, IN49[4], w2428, w2429);
  FullAdder U721 (w2429, w2382, IN50[3], w2430, w2431);
  FullAdder U722 (w2431, w2384, IN51[2], w2432, w2433);
  FullAdder U723 (w2433, w2386, IN52[1], w2434, w2435);
  FullAdder U724 (w2435, w2387, IN53[0], w2436, w2437);
  HalfAdder U725 (w2390, IN30[24], Out1[30], w2439);
  FullAdder U726 (w2439, w2392, IN31[23], w2440, w2441);
  FullAdder U727 (w2441, w2394, IN32[22], w2442, w2443);
  FullAdder U728 (w2443, w2396, IN33[21], w2444, w2445);
  FullAdder U729 (w2445, w2398, IN34[20], w2446, w2447);
  FullAdder U730 (w2447, w2400, IN35[19], w2448, w2449);
  FullAdder U731 (w2449, w2402, IN36[18], w2450, w2451);
  FullAdder U732 (w2451, w2404, IN37[17], w2452, w2453);
  FullAdder U733 (w2453, w2406, IN38[16], w2454, w2455);
  FullAdder U734 (w2455, w2408, IN39[15], w2456, w2457);
  FullAdder U735 (w2457, w2410, IN40[14], w2458, w2459);
  FullAdder U736 (w2459, w2412, IN41[13], w2460, w2461);
  FullAdder U737 (w2461, w2414, IN42[12], w2462, w2463);
  FullAdder U738 (w2463, w2416, IN43[11], w2464, w2465);
  FullAdder U739 (w2465, w2418, IN44[10], w2466, w2467);
  FullAdder U740 (w2467, w2420, IN45[9], w2468, w2469);
  FullAdder U741 (w2469, w2422, IN46[8], w2470, w2471);
  FullAdder U742 (w2471, w2424, IN47[7], w2472, w2473);
  FullAdder U743 (w2473, w2426, IN48[6], w2474, w2475);
  FullAdder U744 (w2475, w2428, IN49[5], w2476, w2477);
  FullAdder U745 (w2477, w2430, IN50[4], w2478, w2479);
  FullAdder U746 (w2479, w2432, IN51[3], w2480, w2481);
  FullAdder U747 (w2481, w2434, IN52[2], w2482, w2483);
  FullAdder U748 (w2483, w2436, IN53[1], w2484, w2485);
  FullAdder U749 (w2485, w2437, IN54[0], w2486, w2487);
  HalfAdder U750 (w2440, IN31[24], Out1[31], w2489);
  FullAdder U751 (w2489, w2442, IN32[23], w2490, w2491);
  FullAdder U752 (w2491, w2444, IN33[22], w2492, w2493);
  FullAdder U753 (w2493, w2446, IN34[21], w2494, w2495);
  FullAdder U754 (w2495, w2448, IN35[20], w2496, w2497);
  FullAdder U755 (w2497, w2450, IN36[19], w2498, w2499);
  FullAdder U756 (w2499, w2452, IN37[18], w2500, w2501);
  FullAdder U757 (w2501, w2454, IN38[17], w2502, w2503);
  FullAdder U758 (w2503, w2456, IN39[16], w2504, w2505);
  FullAdder U759 (w2505, w2458, IN40[15], w2506, w2507);
  FullAdder U760 (w2507, w2460, IN41[14], w2508, w2509);
  FullAdder U761 (w2509, w2462, IN42[13], w2510, w2511);
  FullAdder U762 (w2511, w2464, IN43[12], w2512, w2513);
  FullAdder U763 (w2513, w2466, IN44[11], w2514, w2515);
  FullAdder U764 (w2515, w2468, IN45[10], w2516, w2517);
  FullAdder U765 (w2517, w2470, IN46[9], w2518, w2519);
  FullAdder U766 (w2519, w2472, IN47[8], w2520, w2521);
  FullAdder U767 (w2521, w2474, IN48[7], w2522, w2523);
  FullAdder U768 (w2523, w2476, IN49[6], w2524, w2525);
  FullAdder U769 (w2525, w2478, IN50[5], w2526, w2527);
  FullAdder U770 (w2527, w2480, IN51[4], w2528, w2529);
  FullAdder U771 (w2529, w2482, IN52[3], w2530, w2531);
  FullAdder U772 (w2531, w2484, IN53[2], w2532, w2533);
  FullAdder U773 (w2533, w2486, IN54[1], w2534, w2535);
  FullAdder U774 (w2535, w2487, IN55[0], w2536, w2537);
  HalfAdder U775 (w2490, IN32[24], Out1[32], w2539);
  FullAdder U776 (w2539, w2492, IN33[23], w2540, w2541);
  FullAdder U777 (w2541, w2494, IN34[22], w2542, w2543);
  FullAdder U778 (w2543, w2496, IN35[21], w2544, w2545);
  FullAdder U779 (w2545, w2498, IN36[20], w2546, w2547);
  FullAdder U780 (w2547, w2500, IN37[19], w2548, w2549);
  FullAdder U781 (w2549, w2502, IN38[18], w2550, w2551);
  FullAdder U782 (w2551, w2504, IN39[17], w2552, w2553);
  FullAdder U783 (w2553, w2506, IN40[16], w2554, w2555);
  FullAdder U784 (w2555, w2508, IN41[15], w2556, w2557);
  FullAdder U785 (w2557, w2510, IN42[14], w2558, w2559);
  FullAdder U786 (w2559, w2512, IN43[13], w2560, w2561);
  FullAdder U787 (w2561, w2514, IN44[12], w2562, w2563);
  FullAdder U788 (w2563, w2516, IN45[11], w2564, w2565);
  FullAdder U789 (w2565, w2518, IN46[10], w2566, w2567);
  FullAdder U790 (w2567, w2520, IN47[9], w2568, w2569);
  FullAdder U791 (w2569, w2522, IN48[8], w2570, w2571);
  FullAdder U792 (w2571, w2524, IN49[7], w2572, w2573);
  FullAdder U793 (w2573, w2526, IN50[6], w2574, w2575);
  FullAdder U794 (w2575, w2528, IN51[5], w2576, w2577);
  FullAdder U795 (w2577, w2530, IN52[4], w2578, w2579);
  FullAdder U796 (w2579, w2532, IN53[3], w2580, w2581);
  FullAdder U797 (w2581, w2534, IN54[2], w2582, w2583);
  FullAdder U798 (w2583, w2536, IN55[1], w2584, w2585);
  FullAdder U799 (w2585, w2537, IN56[0], w2586, w2587);
  HalfAdder U800 (w2540, IN33[24], Out1[33], w2589);
  FullAdder U801 (w2589, w2542, IN34[23], w2590, w2591);
  FullAdder U802 (w2591, w2544, IN35[22], w2592, w2593);
  FullAdder U803 (w2593, w2546, IN36[21], w2594, w2595);
  FullAdder U804 (w2595, w2548, IN37[20], w2596, w2597);
  FullAdder U805 (w2597, w2550, IN38[19], w2598, w2599);
  FullAdder U806 (w2599, w2552, IN39[18], w2600, w2601);
  FullAdder U807 (w2601, w2554, IN40[17], w2602, w2603);
  FullAdder U808 (w2603, w2556, IN41[16], w2604, w2605);
  FullAdder U809 (w2605, w2558, IN42[15], w2606, w2607);
  FullAdder U810 (w2607, w2560, IN43[14], w2608, w2609);
  FullAdder U811 (w2609, w2562, IN44[13], w2610, w2611);
  FullAdder U812 (w2611, w2564, IN45[12], w2612, w2613);
  FullAdder U813 (w2613, w2566, IN46[11], w2614, w2615);
  FullAdder U814 (w2615, w2568, IN47[10], w2616, w2617);
  FullAdder U815 (w2617, w2570, IN48[9], w2618, w2619);
  FullAdder U816 (w2619, w2572, IN49[8], w2620, w2621);
  FullAdder U817 (w2621, w2574, IN50[7], w2622, w2623);
  FullAdder U818 (w2623, w2576, IN51[6], w2624, w2625);
  FullAdder U819 (w2625, w2578, IN52[5], w2626, w2627);
  FullAdder U820 (w2627, w2580, IN53[4], w2628, w2629);
  FullAdder U821 (w2629, w2582, IN54[3], w2630, w2631);
  FullAdder U822 (w2631, w2584, IN55[2], w2632, w2633);
  FullAdder U823 (w2633, w2586, IN56[1], w2634, w2635);
  FullAdder U824 (w2635, w2587, IN57[0], w2636, w2637);
  HalfAdder U825 (w2590, IN34[24], Out1[34], w2639);
  FullAdder U826 (w2639, w2592, IN35[23], w2640, w2641);
  FullAdder U827 (w2641, w2594, IN36[22], w2642, w2643);
  FullAdder U828 (w2643, w2596, IN37[21], w2644, w2645);
  FullAdder U829 (w2645, w2598, IN38[20], w2646, w2647);
  FullAdder U830 (w2647, w2600, IN39[19], w2648, w2649);
  FullAdder U831 (w2649, w2602, IN40[18], w2650, w2651);
  FullAdder U832 (w2651, w2604, IN41[17], w2652, w2653);
  FullAdder U833 (w2653, w2606, IN42[16], w2654, w2655);
  FullAdder U834 (w2655, w2608, IN43[15], w2656, w2657);
  FullAdder U835 (w2657, w2610, IN44[14], w2658, w2659);
  FullAdder U836 (w2659, w2612, IN45[13], w2660, w2661);
  FullAdder U837 (w2661, w2614, IN46[12], w2662, w2663);
  FullAdder U838 (w2663, w2616, IN47[11], w2664, w2665);
  FullAdder U839 (w2665, w2618, IN48[10], w2666, w2667);
  FullAdder U840 (w2667, w2620, IN49[9], w2668, w2669);
  FullAdder U841 (w2669, w2622, IN50[8], w2670, w2671);
  FullAdder U842 (w2671, w2624, IN51[7], w2672, w2673);
  FullAdder U843 (w2673, w2626, IN52[6], w2674, w2675);
  FullAdder U844 (w2675, w2628, IN53[5], w2676, w2677);
  FullAdder U845 (w2677, w2630, IN54[4], w2678, w2679);
  FullAdder U846 (w2679, w2632, IN55[3], w2680, w2681);
  FullAdder U847 (w2681, w2634, IN56[2], w2682, w2683);
  FullAdder U848 (w2683, w2636, IN57[1], w2684, w2685);
  FullAdder U849 (w2685, w2637, IN58[0], w2686, w2687);
  HalfAdder U850 (w2640, IN35[24], Out1[35], w2689);
  FullAdder U851 (w2689, w2642, IN36[23], w2690, w2691);
  FullAdder U852 (w2691, w2644, IN37[22], w2692, w2693);
  FullAdder U853 (w2693, w2646, IN38[21], w2694, w2695);
  FullAdder U854 (w2695, w2648, IN39[20], w2696, w2697);
  FullAdder U855 (w2697, w2650, IN40[19], w2698, w2699);
  FullAdder U856 (w2699, w2652, IN41[18], w2700, w2701);
  FullAdder U857 (w2701, w2654, IN42[17], w2702, w2703);
  FullAdder U858 (w2703, w2656, IN43[16], w2704, w2705);
  FullAdder U859 (w2705, w2658, IN44[15], w2706, w2707);
  FullAdder U860 (w2707, w2660, IN45[14], w2708, w2709);
  FullAdder U861 (w2709, w2662, IN46[13], w2710, w2711);
  FullAdder U862 (w2711, w2664, IN47[12], w2712, w2713);
  FullAdder U863 (w2713, w2666, IN48[11], w2714, w2715);
  FullAdder U864 (w2715, w2668, IN49[10], w2716, w2717);
  FullAdder U865 (w2717, w2670, IN50[9], w2718, w2719);
  FullAdder U866 (w2719, w2672, IN51[8], w2720, w2721);
  FullAdder U867 (w2721, w2674, IN52[7], w2722, w2723);
  FullAdder U868 (w2723, w2676, IN53[6], w2724, w2725);
  FullAdder U869 (w2725, w2678, IN54[5], w2726, w2727);
  FullAdder U870 (w2727, w2680, IN55[4], w2728, w2729);
  FullAdder U871 (w2729, w2682, IN56[3], w2730, w2731);
  FullAdder U872 (w2731, w2684, IN57[2], w2732, w2733);
  FullAdder U873 (w2733, w2686, IN58[1], w2734, w2735);
  FullAdder U874 (w2735, w2687, IN59[0], w2736, w2737);
  HalfAdder U875 (w2690, IN36[24], Out1[36], w2739);
  FullAdder U876 (w2739, w2692, IN37[23], w2740, w2741);
  FullAdder U877 (w2741, w2694, IN38[22], w2742, w2743);
  FullAdder U878 (w2743, w2696, IN39[21], w2744, w2745);
  FullAdder U879 (w2745, w2698, IN40[20], w2746, w2747);
  FullAdder U880 (w2747, w2700, IN41[19], w2748, w2749);
  FullAdder U881 (w2749, w2702, IN42[18], w2750, w2751);
  FullAdder U882 (w2751, w2704, IN43[17], w2752, w2753);
  FullAdder U883 (w2753, w2706, IN44[16], w2754, w2755);
  FullAdder U884 (w2755, w2708, IN45[15], w2756, w2757);
  FullAdder U885 (w2757, w2710, IN46[14], w2758, w2759);
  FullAdder U886 (w2759, w2712, IN47[13], w2760, w2761);
  FullAdder U887 (w2761, w2714, IN48[12], w2762, w2763);
  FullAdder U888 (w2763, w2716, IN49[11], w2764, w2765);
  FullAdder U889 (w2765, w2718, IN50[10], w2766, w2767);
  FullAdder U890 (w2767, w2720, IN51[9], w2768, w2769);
  FullAdder U891 (w2769, w2722, IN52[8], w2770, w2771);
  FullAdder U892 (w2771, w2724, IN53[7], w2772, w2773);
  FullAdder U893 (w2773, w2726, IN54[6], w2774, w2775);
  FullAdder U894 (w2775, w2728, IN55[5], w2776, w2777);
  FullAdder U895 (w2777, w2730, IN56[4], w2778, w2779);
  FullAdder U896 (w2779, w2732, IN57[3], w2780, w2781);
  FullAdder U897 (w2781, w2734, IN58[2], w2782, w2783);
  FullAdder U898 (w2783, w2736, IN59[1], w2784, w2785);
  FullAdder U899 (w2785, w2737, IN60[0], w2786, w2787);
  HalfAdder U900 (w2740, IN37[24], Out1[37], w2789);
  FullAdder U901 (w2789, w2742, IN38[23], Out1[38], w2791);
  FullAdder U902 (w2791, w2744, IN39[22], Out1[39], w2793);
  FullAdder U903 (w2793, w2746, IN40[21], Out1[40], w2795);
  FullAdder U904 (w2795, w2748, IN41[20], Out1[41], w2797);
  FullAdder U905 (w2797, w2750, IN42[19], Out1[42], w2799);
  FullAdder U906 (w2799, w2752, IN43[18], Out1[43], w2801);
  FullAdder U907 (w2801, w2754, IN44[17], Out1[44], w2803);
  FullAdder U908 (w2803, w2756, IN45[16], Out1[45], w2805);
  FullAdder U909 (w2805, w2758, IN46[15], Out1[46], w2807);
  FullAdder U910 (w2807, w2760, IN47[14], Out1[47], w2809);
  FullAdder U911 (w2809, w2762, IN48[13], Out1[48], w2811);
  FullAdder U912 (w2811, w2764, IN49[12], Out1[49], w2813);
  FullAdder U913 (w2813, w2766, IN50[11], Out1[50], w2815);
  FullAdder U914 (w2815, w2768, IN51[10], Out1[51], w2817);
  FullAdder U915 (w2817, w2770, IN52[9], Out1[52], w2819);
  FullAdder U916 (w2819, w2772, IN53[8], Out1[53], w2821);
  FullAdder U917 (w2821, w2774, IN54[7], Out1[54], w2823);
  FullAdder U918 (w2823, w2776, IN55[6], Out1[55], w2825);
  FullAdder U919 (w2825, w2778, IN56[5], Out1[56], w2827);
  FullAdder U920 (w2827, w2780, IN57[4], Out1[57], w2829);
  FullAdder U921 (w2829, w2782, IN58[3], Out1[58], w2831);
  FullAdder U922 (w2831, w2784, IN59[2], Out1[59], w2833);
  FullAdder U923 (w2833, w2786, IN60[1], Out1[60], w2835);
  FullAdder U924 (w2835, w2787, IN61[0], Out1[61], Out1[62]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN26[25];
  assign Out2[1] = IN27[25];
  assign Out2[2] = IN28[25];
  assign Out2[3] = IN29[25];
  assign Out2[4] = IN30[25];
  assign Out2[5] = IN31[25];
  assign Out2[6] = IN32[25];
  assign Out2[7] = IN33[25];
  assign Out2[8] = IN34[25];
  assign Out2[9] = IN35[25];
  assign Out2[10] = IN36[25];
  assign Out2[11] = IN37[25];
  assign Out2[12] = IN38[24];
  assign Out2[13] = IN39[23];
  assign Out2[14] = IN40[22];
  assign Out2[15] = IN41[21];
  assign Out2[16] = IN42[20];
  assign Out2[17] = IN43[19];
  assign Out2[18] = IN44[18];
  assign Out2[19] = IN45[17];
  assign Out2[20] = IN46[16];
  assign Out2[21] = IN47[15];
  assign Out2[22] = IN48[14];
  assign Out2[23] = IN49[13];
  assign Out2[24] = IN50[12];
  assign Out2[25] = IN51[11];
  assign Out2[26] = IN52[10];
  assign Out2[27] = IN53[9];
  assign Out2[28] = IN54[8];
  assign Out2[29] = IN55[7];
  assign Out2[30] = IN56[6];
  assign Out2[31] = IN57[5];
  assign Out2[32] = IN58[4];
  assign Out2[33] = IN59[3];
  assign Out2[34] = IN60[2];
  assign Out2[35] = IN61[1];
  assign Out2[36] = IN62[0];

endmodule
module RC_37_37(IN1, IN2, Out);
  input [36:0] IN1;
  input [36:0] IN2;
  output [37:0] Out;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w75);
  FullAdder U1 (IN1[1], IN2[1], w75, Out[1], w77);
  FullAdder U2 (IN1[2], IN2[2], w77, Out[2], w79);
  FullAdder U3 (IN1[3], IN2[3], w79, Out[3], w81);
  FullAdder U4 (IN1[4], IN2[4], w81, Out[4], w83);
  FullAdder U5 (IN1[5], IN2[5], w83, Out[5], w85);
  FullAdder U6 (IN1[6], IN2[6], w85, Out[6], w87);
  FullAdder U7 (IN1[7], IN2[7], w87, Out[7], w89);
  FullAdder U8 (IN1[8], IN2[8], w89, Out[8], w91);
  FullAdder U9 (IN1[9], IN2[9], w91, Out[9], w93);
  FullAdder U10 (IN1[10], IN2[10], w93, Out[10], w95);
  FullAdder U11 (IN1[11], IN2[11], w95, Out[11], w97);
  FullAdder U12 (IN1[12], IN2[12], w97, Out[12], w99);
  FullAdder U13 (IN1[13], IN2[13], w99, Out[13], w101);
  FullAdder U14 (IN1[14], IN2[14], w101, Out[14], w103);
  FullAdder U15 (IN1[15], IN2[15], w103, Out[15], w105);
  FullAdder U16 (IN1[16], IN2[16], w105, Out[16], w107);
  FullAdder U17 (IN1[17], IN2[17], w107, Out[17], w109);
  FullAdder U18 (IN1[18], IN2[18], w109, Out[18], w111);
  FullAdder U19 (IN1[19], IN2[19], w111, Out[19], w113);
  FullAdder U20 (IN1[20], IN2[20], w113, Out[20], w115);
  FullAdder U21 (IN1[21], IN2[21], w115, Out[21], w117);
  FullAdder U22 (IN1[22], IN2[22], w117, Out[22], w119);
  FullAdder U23 (IN1[23], IN2[23], w119, Out[23], w121);
  FullAdder U24 (IN1[24], IN2[24], w121, Out[24], w123);
  FullAdder U25 (IN1[25], IN2[25], w123, Out[25], w125);
  FullAdder U26 (IN1[26], IN2[26], w125, Out[26], w127);
  FullAdder U27 (IN1[27], IN2[27], w127, Out[27], w129);
  FullAdder U28 (IN1[28], IN2[28], w129, Out[28], w131);
  FullAdder U29 (IN1[29], IN2[29], w131, Out[29], w133);
  FullAdder U30 (IN1[30], IN2[30], w133, Out[30], w135);
  FullAdder U31 (IN1[31], IN2[31], w135, Out[31], w137);
  FullAdder U32 (IN1[32], IN2[32], w137, Out[32], w139);
  FullAdder U33 (IN1[33], IN2[33], w139, Out[33], w141);
  FullAdder U34 (IN1[34], IN2[34], w141, Out[34], w143);
  FullAdder U35 (IN1[35], IN2[35], w143, Out[35], w145);
  FullAdder U36 (IN1[36], IN2[36], w145, Out[36], Out[37]);

endmodule
module NR_26_38(IN1, IN2, Out);
  input [25:0] IN1;
  input [37:0] IN2;
  output [63:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [25:0] P26;
  wire [25:0] P27;
  wire [25:0] P28;
  wire [25:0] P29;
  wire [25:0] P30;
  wire [25:0] P31;
  wire [25:0] P32;
  wire [25:0] P33;
  wire [25:0] P34;
  wire [25:0] P35;
  wire [25:0] P36;
  wire [25:0] P37;
  wire [24:0] P38;
  wire [23:0] P39;
  wire [22:0] P40;
  wire [21:0] P41;
  wire [20:0] P42;
  wire [19:0] P43;
  wire [18:0] P44;
  wire [17:0] P45;
  wire [16:0] P46;
  wire [15:0] P47;
  wire [14:0] P48;
  wire [13:0] P49;
  wire [12:0] P50;
  wire [11:0] P51;
  wire [10:0] P52;
  wire [9:0] P53;
  wire [8:0] P54;
  wire [7:0] P55;
  wire [6:0] P56;
  wire [5:0] P57;
  wire [4:0] P58;
  wire [3:0] P59;
  wire [2:0] P60;
  wire [1:0] P61;
  wire [0:0] P62;
  wire [62:0] R1;
  wire [36:0] R2;
  wire [63:0] aOut;
  U_SP_26_38 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, R1, R2);
  RC_37_37 S2 (R1[62:26], R2, aOut[63:26]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign Out = aOut[63:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
