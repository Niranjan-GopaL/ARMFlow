
module NR_1_61(
    input [0:0]IN1,
    input [60:0]IN2,
    output [60:0]Out
);
    assign Out = IN2;
endmodule
