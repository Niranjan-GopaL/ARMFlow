
module customAdder34_0(
    input [33 : 0] A,
    input [33 : 0] B,
    output [34 : 0] Sum
);

    assign Sum = A+B;

endmodule
