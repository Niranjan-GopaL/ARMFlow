
module NR_1_64(
    input [0:0]IN1,
    input [63:0]IN2,
    output [63:0]Out
);
    assign Out = IN2;
endmodule
