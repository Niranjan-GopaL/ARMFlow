
module NR_1_44(
    input [0:0]IN1,
    input [43:0]IN2,
    output [43:0]Out
);
    assign Out = IN2;
endmodule
