
module multiplier32bit_38(
    input [31:0] A, 
    input [31:0] B, 
    output [63:0] P
);
    
    wire [24:0] A_H, B_H;
    wire [6:0] A_L, B_L;
    
    assign A_H = A[31:7];
    assign B_H = B[31:7];
    assign A_L = A[6:0];
    assign B_L = B[6:0];
    
    
    wire [49:0] P1;
    wire [31:0] P2, P3;
    wire [13:0] P4;
    
    NR_25_25 M1(A_H, B_H, P1);
    NR_25_7 M2(A_H, B_L, P2);
    NR_7_25 M3(A_L, B_H, P3);
    rr_7x7_4 M4(A_L, B_L, P4);
    
    wire[6:0] P4_L;
    wire[6:0] P4_H;

    wire[56:0] operand1;
    wire[32:0] operand2;
    wire[57:0] out;
    
    assign P4_L = P4[6:0];
    assign P4_H = P4[13:7];
    assign operand1 = {P1,P4_H};

    customAdder32_0 adder1(
        P2,
        P3,
        operand2
    );

    customAdder57_24 adder2(
        operand1,
        operand2,
        out
    );
    assign P = {out[56:0],P4_L};
endmodule
        
module rr_7x7_4(
    input [6:0] A, 
    input [6:0] B, 
    output [13:0] P
);
    
    wire [1:0] A_H, B_H;
    wire [4:0] A_L, B_L;
    
    assign A_H = A[6:5];
    assign B_H = B[6:5];
    assign A_L = A[4:0];
    assign B_L = B[4:0];
    
    wire [3:0] P1;
    wire [6:0] P2, P3;
    wire [9:0] P4;
    
    NR_2_2 M1(A_H, B_H, P1);
    NR_2_5 M2(A_H, B_L, P2);
    NR_5_2 M3(A_L, B_H, P3);
    NR_5_5 M4(A_L, B_L, P4);
    
    wire[4:0] P4_L;
    wire[4:0] P4_H;

    wire[8:0] operand1;
    wire[7:0] operand2;
    wire[9:0] out;
    
    assign P4_L = P4[4:0];
    assign P4_H = P4[9:5];
    assign operand1 = {P1,P4_H};

    customAdder7_0 adder1(
        P2,
        P3,
        operand2
    );

    customAdder9_1 adder2(
        operand1,
        operand2,
        out
    );
    assign P = {out[8:0],P4_L};
endmodule
        