
module NR_63_1(
    input [62:0]IN1,
    input [0:0]IN2,
    output [62:0]Out
);
    assign Out = IN2;
endmodule
