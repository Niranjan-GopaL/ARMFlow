//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 51
  second input length: 35
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_51_35(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84);
  input [50:0] IN1;
  input [34:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [29:0] P29;
  output [30:0] P30;
  output [31:0] P31;
  output [32:0] P32;
  output [33:0] P33;
  output [34:0] P34;
  output [34:0] P35;
  output [34:0] P36;
  output [34:0] P37;
  output [34:0] P38;
  output [34:0] P39;
  output [34:0] P40;
  output [34:0] P41;
  output [34:0] P42;
  output [34:0] P43;
  output [34:0] P44;
  output [34:0] P45;
  output [34:0] P46;
  output [34:0] P47;
  output [34:0] P48;
  output [34:0] P49;
  output [34:0] P50;
  output [33:0] P51;
  output [32:0] P52;
  output [31:0] P53;
  output [30:0] P54;
  output [29:0] P55;
  output [28:0] P56;
  output [27:0] P57;
  output [26:0] P58;
  output [25:0] P59;
  output [24:0] P60;
  output [23:0] P61;
  output [22:0] P62;
  output [21:0] P63;
  output [20:0] P64;
  output [19:0] P65;
  output [18:0] P66;
  output [17:0] P67;
  output [16:0] P68;
  output [15:0] P69;
  output [14:0] P70;
  output [13:0] P71;
  output [12:0] P72;
  output [11:0] P73;
  output [10:0] P74;
  output [9:0] P75;
  output [8:0] P76;
  output [7:0] P77;
  output [6:0] P78;
  output [5:0] P79;
  output [4:0] P80;
  output [3:0] P81;
  output [2:0] P82;
  output [1:0] P83;
  output [0:0] P84;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[0] = IN1[1]&IN2[34];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[1] = IN1[2]&IN2[33];
  assign P36[0] = IN1[2]&IN2[34];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[2] = IN1[3]&IN2[32];
  assign P36[1] = IN1[3]&IN2[33];
  assign P37[0] = IN1[3]&IN2[34];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[3] = IN1[4]&IN2[31];
  assign P36[2] = IN1[4]&IN2[32];
  assign P37[1] = IN1[4]&IN2[33];
  assign P38[0] = IN1[4]&IN2[34];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[4] = IN1[5]&IN2[30];
  assign P36[3] = IN1[5]&IN2[31];
  assign P37[2] = IN1[5]&IN2[32];
  assign P38[1] = IN1[5]&IN2[33];
  assign P39[0] = IN1[5]&IN2[34];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[5] = IN1[6]&IN2[29];
  assign P36[4] = IN1[6]&IN2[30];
  assign P37[3] = IN1[6]&IN2[31];
  assign P38[2] = IN1[6]&IN2[32];
  assign P39[1] = IN1[6]&IN2[33];
  assign P40[0] = IN1[6]&IN2[34];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[6] = IN1[7]&IN2[28];
  assign P36[5] = IN1[7]&IN2[29];
  assign P37[4] = IN1[7]&IN2[30];
  assign P38[3] = IN1[7]&IN2[31];
  assign P39[2] = IN1[7]&IN2[32];
  assign P40[1] = IN1[7]&IN2[33];
  assign P41[0] = IN1[7]&IN2[34];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[7] = IN1[8]&IN2[27];
  assign P36[6] = IN1[8]&IN2[28];
  assign P37[5] = IN1[8]&IN2[29];
  assign P38[4] = IN1[8]&IN2[30];
  assign P39[3] = IN1[8]&IN2[31];
  assign P40[2] = IN1[8]&IN2[32];
  assign P41[1] = IN1[8]&IN2[33];
  assign P42[0] = IN1[8]&IN2[34];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[8] = IN1[9]&IN2[26];
  assign P36[7] = IN1[9]&IN2[27];
  assign P37[6] = IN1[9]&IN2[28];
  assign P38[5] = IN1[9]&IN2[29];
  assign P39[4] = IN1[9]&IN2[30];
  assign P40[3] = IN1[9]&IN2[31];
  assign P41[2] = IN1[9]&IN2[32];
  assign P42[1] = IN1[9]&IN2[33];
  assign P43[0] = IN1[9]&IN2[34];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[9] = IN1[10]&IN2[25];
  assign P36[8] = IN1[10]&IN2[26];
  assign P37[7] = IN1[10]&IN2[27];
  assign P38[6] = IN1[10]&IN2[28];
  assign P39[5] = IN1[10]&IN2[29];
  assign P40[4] = IN1[10]&IN2[30];
  assign P41[3] = IN1[10]&IN2[31];
  assign P42[2] = IN1[10]&IN2[32];
  assign P43[1] = IN1[10]&IN2[33];
  assign P44[0] = IN1[10]&IN2[34];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[10] = IN1[11]&IN2[24];
  assign P36[9] = IN1[11]&IN2[25];
  assign P37[8] = IN1[11]&IN2[26];
  assign P38[7] = IN1[11]&IN2[27];
  assign P39[6] = IN1[11]&IN2[28];
  assign P40[5] = IN1[11]&IN2[29];
  assign P41[4] = IN1[11]&IN2[30];
  assign P42[3] = IN1[11]&IN2[31];
  assign P43[2] = IN1[11]&IN2[32];
  assign P44[1] = IN1[11]&IN2[33];
  assign P45[0] = IN1[11]&IN2[34];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[11] = IN1[12]&IN2[23];
  assign P36[10] = IN1[12]&IN2[24];
  assign P37[9] = IN1[12]&IN2[25];
  assign P38[8] = IN1[12]&IN2[26];
  assign P39[7] = IN1[12]&IN2[27];
  assign P40[6] = IN1[12]&IN2[28];
  assign P41[5] = IN1[12]&IN2[29];
  assign P42[4] = IN1[12]&IN2[30];
  assign P43[3] = IN1[12]&IN2[31];
  assign P44[2] = IN1[12]&IN2[32];
  assign P45[1] = IN1[12]&IN2[33];
  assign P46[0] = IN1[12]&IN2[34];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[12] = IN1[13]&IN2[22];
  assign P36[11] = IN1[13]&IN2[23];
  assign P37[10] = IN1[13]&IN2[24];
  assign P38[9] = IN1[13]&IN2[25];
  assign P39[8] = IN1[13]&IN2[26];
  assign P40[7] = IN1[13]&IN2[27];
  assign P41[6] = IN1[13]&IN2[28];
  assign P42[5] = IN1[13]&IN2[29];
  assign P43[4] = IN1[13]&IN2[30];
  assign P44[3] = IN1[13]&IN2[31];
  assign P45[2] = IN1[13]&IN2[32];
  assign P46[1] = IN1[13]&IN2[33];
  assign P47[0] = IN1[13]&IN2[34];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[13] = IN1[14]&IN2[21];
  assign P36[12] = IN1[14]&IN2[22];
  assign P37[11] = IN1[14]&IN2[23];
  assign P38[10] = IN1[14]&IN2[24];
  assign P39[9] = IN1[14]&IN2[25];
  assign P40[8] = IN1[14]&IN2[26];
  assign P41[7] = IN1[14]&IN2[27];
  assign P42[6] = IN1[14]&IN2[28];
  assign P43[5] = IN1[14]&IN2[29];
  assign P44[4] = IN1[14]&IN2[30];
  assign P45[3] = IN1[14]&IN2[31];
  assign P46[2] = IN1[14]&IN2[32];
  assign P47[1] = IN1[14]&IN2[33];
  assign P48[0] = IN1[14]&IN2[34];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[14] = IN1[15]&IN2[20];
  assign P36[13] = IN1[15]&IN2[21];
  assign P37[12] = IN1[15]&IN2[22];
  assign P38[11] = IN1[15]&IN2[23];
  assign P39[10] = IN1[15]&IN2[24];
  assign P40[9] = IN1[15]&IN2[25];
  assign P41[8] = IN1[15]&IN2[26];
  assign P42[7] = IN1[15]&IN2[27];
  assign P43[6] = IN1[15]&IN2[28];
  assign P44[5] = IN1[15]&IN2[29];
  assign P45[4] = IN1[15]&IN2[30];
  assign P46[3] = IN1[15]&IN2[31];
  assign P47[2] = IN1[15]&IN2[32];
  assign P48[1] = IN1[15]&IN2[33];
  assign P49[0] = IN1[15]&IN2[34];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[15] = IN1[16]&IN2[19];
  assign P36[14] = IN1[16]&IN2[20];
  assign P37[13] = IN1[16]&IN2[21];
  assign P38[12] = IN1[16]&IN2[22];
  assign P39[11] = IN1[16]&IN2[23];
  assign P40[10] = IN1[16]&IN2[24];
  assign P41[9] = IN1[16]&IN2[25];
  assign P42[8] = IN1[16]&IN2[26];
  assign P43[7] = IN1[16]&IN2[27];
  assign P44[6] = IN1[16]&IN2[28];
  assign P45[5] = IN1[16]&IN2[29];
  assign P46[4] = IN1[16]&IN2[30];
  assign P47[3] = IN1[16]&IN2[31];
  assign P48[2] = IN1[16]&IN2[32];
  assign P49[1] = IN1[16]&IN2[33];
  assign P50[0] = IN1[16]&IN2[34];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[16] = IN1[17]&IN2[18];
  assign P36[15] = IN1[17]&IN2[19];
  assign P37[14] = IN1[17]&IN2[20];
  assign P38[13] = IN1[17]&IN2[21];
  assign P39[12] = IN1[17]&IN2[22];
  assign P40[11] = IN1[17]&IN2[23];
  assign P41[10] = IN1[17]&IN2[24];
  assign P42[9] = IN1[17]&IN2[25];
  assign P43[8] = IN1[17]&IN2[26];
  assign P44[7] = IN1[17]&IN2[27];
  assign P45[6] = IN1[17]&IN2[28];
  assign P46[5] = IN1[17]&IN2[29];
  assign P47[4] = IN1[17]&IN2[30];
  assign P48[3] = IN1[17]&IN2[31];
  assign P49[2] = IN1[17]&IN2[32];
  assign P50[1] = IN1[17]&IN2[33];
  assign P51[0] = IN1[17]&IN2[34];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[17] = IN1[18]&IN2[17];
  assign P36[16] = IN1[18]&IN2[18];
  assign P37[15] = IN1[18]&IN2[19];
  assign P38[14] = IN1[18]&IN2[20];
  assign P39[13] = IN1[18]&IN2[21];
  assign P40[12] = IN1[18]&IN2[22];
  assign P41[11] = IN1[18]&IN2[23];
  assign P42[10] = IN1[18]&IN2[24];
  assign P43[9] = IN1[18]&IN2[25];
  assign P44[8] = IN1[18]&IN2[26];
  assign P45[7] = IN1[18]&IN2[27];
  assign P46[6] = IN1[18]&IN2[28];
  assign P47[5] = IN1[18]&IN2[29];
  assign P48[4] = IN1[18]&IN2[30];
  assign P49[3] = IN1[18]&IN2[31];
  assign P50[2] = IN1[18]&IN2[32];
  assign P51[1] = IN1[18]&IN2[33];
  assign P52[0] = IN1[18]&IN2[34];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[18] = IN1[19]&IN2[16];
  assign P36[17] = IN1[19]&IN2[17];
  assign P37[16] = IN1[19]&IN2[18];
  assign P38[15] = IN1[19]&IN2[19];
  assign P39[14] = IN1[19]&IN2[20];
  assign P40[13] = IN1[19]&IN2[21];
  assign P41[12] = IN1[19]&IN2[22];
  assign P42[11] = IN1[19]&IN2[23];
  assign P43[10] = IN1[19]&IN2[24];
  assign P44[9] = IN1[19]&IN2[25];
  assign P45[8] = IN1[19]&IN2[26];
  assign P46[7] = IN1[19]&IN2[27];
  assign P47[6] = IN1[19]&IN2[28];
  assign P48[5] = IN1[19]&IN2[29];
  assign P49[4] = IN1[19]&IN2[30];
  assign P50[3] = IN1[19]&IN2[31];
  assign P51[2] = IN1[19]&IN2[32];
  assign P52[1] = IN1[19]&IN2[33];
  assign P53[0] = IN1[19]&IN2[34];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[19] = IN1[20]&IN2[15];
  assign P36[18] = IN1[20]&IN2[16];
  assign P37[17] = IN1[20]&IN2[17];
  assign P38[16] = IN1[20]&IN2[18];
  assign P39[15] = IN1[20]&IN2[19];
  assign P40[14] = IN1[20]&IN2[20];
  assign P41[13] = IN1[20]&IN2[21];
  assign P42[12] = IN1[20]&IN2[22];
  assign P43[11] = IN1[20]&IN2[23];
  assign P44[10] = IN1[20]&IN2[24];
  assign P45[9] = IN1[20]&IN2[25];
  assign P46[8] = IN1[20]&IN2[26];
  assign P47[7] = IN1[20]&IN2[27];
  assign P48[6] = IN1[20]&IN2[28];
  assign P49[5] = IN1[20]&IN2[29];
  assign P50[4] = IN1[20]&IN2[30];
  assign P51[3] = IN1[20]&IN2[31];
  assign P52[2] = IN1[20]&IN2[32];
  assign P53[1] = IN1[20]&IN2[33];
  assign P54[0] = IN1[20]&IN2[34];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[20] = IN1[21]&IN2[14];
  assign P36[19] = IN1[21]&IN2[15];
  assign P37[18] = IN1[21]&IN2[16];
  assign P38[17] = IN1[21]&IN2[17];
  assign P39[16] = IN1[21]&IN2[18];
  assign P40[15] = IN1[21]&IN2[19];
  assign P41[14] = IN1[21]&IN2[20];
  assign P42[13] = IN1[21]&IN2[21];
  assign P43[12] = IN1[21]&IN2[22];
  assign P44[11] = IN1[21]&IN2[23];
  assign P45[10] = IN1[21]&IN2[24];
  assign P46[9] = IN1[21]&IN2[25];
  assign P47[8] = IN1[21]&IN2[26];
  assign P48[7] = IN1[21]&IN2[27];
  assign P49[6] = IN1[21]&IN2[28];
  assign P50[5] = IN1[21]&IN2[29];
  assign P51[4] = IN1[21]&IN2[30];
  assign P52[3] = IN1[21]&IN2[31];
  assign P53[2] = IN1[21]&IN2[32];
  assign P54[1] = IN1[21]&IN2[33];
  assign P55[0] = IN1[21]&IN2[34];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[21] = IN1[22]&IN2[13];
  assign P36[20] = IN1[22]&IN2[14];
  assign P37[19] = IN1[22]&IN2[15];
  assign P38[18] = IN1[22]&IN2[16];
  assign P39[17] = IN1[22]&IN2[17];
  assign P40[16] = IN1[22]&IN2[18];
  assign P41[15] = IN1[22]&IN2[19];
  assign P42[14] = IN1[22]&IN2[20];
  assign P43[13] = IN1[22]&IN2[21];
  assign P44[12] = IN1[22]&IN2[22];
  assign P45[11] = IN1[22]&IN2[23];
  assign P46[10] = IN1[22]&IN2[24];
  assign P47[9] = IN1[22]&IN2[25];
  assign P48[8] = IN1[22]&IN2[26];
  assign P49[7] = IN1[22]&IN2[27];
  assign P50[6] = IN1[22]&IN2[28];
  assign P51[5] = IN1[22]&IN2[29];
  assign P52[4] = IN1[22]&IN2[30];
  assign P53[3] = IN1[22]&IN2[31];
  assign P54[2] = IN1[22]&IN2[32];
  assign P55[1] = IN1[22]&IN2[33];
  assign P56[0] = IN1[22]&IN2[34];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[22] = IN1[23]&IN2[12];
  assign P36[21] = IN1[23]&IN2[13];
  assign P37[20] = IN1[23]&IN2[14];
  assign P38[19] = IN1[23]&IN2[15];
  assign P39[18] = IN1[23]&IN2[16];
  assign P40[17] = IN1[23]&IN2[17];
  assign P41[16] = IN1[23]&IN2[18];
  assign P42[15] = IN1[23]&IN2[19];
  assign P43[14] = IN1[23]&IN2[20];
  assign P44[13] = IN1[23]&IN2[21];
  assign P45[12] = IN1[23]&IN2[22];
  assign P46[11] = IN1[23]&IN2[23];
  assign P47[10] = IN1[23]&IN2[24];
  assign P48[9] = IN1[23]&IN2[25];
  assign P49[8] = IN1[23]&IN2[26];
  assign P50[7] = IN1[23]&IN2[27];
  assign P51[6] = IN1[23]&IN2[28];
  assign P52[5] = IN1[23]&IN2[29];
  assign P53[4] = IN1[23]&IN2[30];
  assign P54[3] = IN1[23]&IN2[31];
  assign P55[2] = IN1[23]&IN2[32];
  assign P56[1] = IN1[23]&IN2[33];
  assign P57[0] = IN1[23]&IN2[34];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[23] = IN1[24]&IN2[11];
  assign P36[22] = IN1[24]&IN2[12];
  assign P37[21] = IN1[24]&IN2[13];
  assign P38[20] = IN1[24]&IN2[14];
  assign P39[19] = IN1[24]&IN2[15];
  assign P40[18] = IN1[24]&IN2[16];
  assign P41[17] = IN1[24]&IN2[17];
  assign P42[16] = IN1[24]&IN2[18];
  assign P43[15] = IN1[24]&IN2[19];
  assign P44[14] = IN1[24]&IN2[20];
  assign P45[13] = IN1[24]&IN2[21];
  assign P46[12] = IN1[24]&IN2[22];
  assign P47[11] = IN1[24]&IN2[23];
  assign P48[10] = IN1[24]&IN2[24];
  assign P49[9] = IN1[24]&IN2[25];
  assign P50[8] = IN1[24]&IN2[26];
  assign P51[7] = IN1[24]&IN2[27];
  assign P52[6] = IN1[24]&IN2[28];
  assign P53[5] = IN1[24]&IN2[29];
  assign P54[4] = IN1[24]&IN2[30];
  assign P55[3] = IN1[24]&IN2[31];
  assign P56[2] = IN1[24]&IN2[32];
  assign P57[1] = IN1[24]&IN2[33];
  assign P58[0] = IN1[24]&IN2[34];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[24] = IN1[25]&IN2[10];
  assign P36[23] = IN1[25]&IN2[11];
  assign P37[22] = IN1[25]&IN2[12];
  assign P38[21] = IN1[25]&IN2[13];
  assign P39[20] = IN1[25]&IN2[14];
  assign P40[19] = IN1[25]&IN2[15];
  assign P41[18] = IN1[25]&IN2[16];
  assign P42[17] = IN1[25]&IN2[17];
  assign P43[16] = IN1[25]&IN2[18];
  assign P44[15] = IN1[25]&IN2[19];
  assign P45[14] = IN1[25]&IN2[20];
  assign P46[13] = IN1[25]&IN2[21];
  assign P47[12] = IN1[25]&IN2[22];
  assign P48[11] = IN1[25]&IN2[23];
  assign P49[10] = IN1[25]&IN2[24];
  assign P50[9] = IN1[25]&IN2[25];
  assign P51[8] = IN1[25]&IN2[26];
  assign P52[7] = IN1[25]&IN2[27];
  assign P53[6] = IN1[25]&IN2[28];
  assign P54[5] = IN1[25]&IN2[29];
  assign P55[4] = IN1[25]&IN2[30];
  assign P56[3] = IN1[25]&IN2[31];
  assign P57[2] = IN1[25]&IN2[32];
  assign P58[1] = IN1[25]&IN2[33];
  assign P59[0] = IN1[25]&IN2[34];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[26] = IN1[26]&IN2[3];
  assign P30[26] = IN1[26]&IN2[4];
  assign P31[26] = IN1[26]&IN2[5];
  assign P32[26] = IN1[26]&IN2[6];
  assign P33[26] = IN1[26]&IN2[7];
  assign P34[26] = IN1[26]&IN2[8];
  assign P35[25] = IN1[26]&IN2[9];
  assign P36[24] = IN1[26]&IN2[10];
  assign P37[23] = IN1[26]&IN2[11];
  assign P38[22] = IN1[26]&IN2[12];
  assign P39[21] = IN1[26]&IN2[13];
  assign P40[20] = IN1[26]&IN2[14];
  assign P41[19] = IN1[26]&IN2[15];
  assign P42[18] = IN1[26]&IN2[16];
  assign P43[17] = IN1[26]&IN2[17];
  assign P44[16] = IN1[26]&IN2[18];
  assign P45[15] = IN1[26]&IN2[19];
  assign P46[14] = IN1[26]&IN2[20];
  assign P47[13] = IN1[26]&IN2[21];
  assign P48[12] = IN1[26]&IN2[22];
  assign P49[11] = IN1[26]&IN2[23];
  assign P50[10] = IN1[26]&IN2[24];
  assign P51[9] = IN1[26]&IN2[25];
  assign P52[8] = IN1[26]&IN2[26];
  assign P53[7] = IN1[26]&IN2[27];
  assign P54[6] = IN1[26]&IN2[28];
  assign P55[5] = IN1[26]&IN2[29];
  assign P56[4] = IN1[26]&IN2[30];
  assign P57[3] = IN1[26]&IN2[31];
  assign P58[2] = IN1[26]&IN2[32];
  assign P59[1] = IN1[26]&IN2[33];
  assign P60[0] = IN1[26]&IN2[34];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[27] = IN1[27]&IN2[2];
  assign P30[27] = IN1[27]&IN2[3];
  assign P31[27] = IN1[27]&IN2[4];
  assign P32[27] = IN1[27]&IN2[5];
  assign P33[27] = IN1[27]&IN2[6];
  assign P34[27] = IN1[27]&IN2[7];
  assign P35[26] = IN1[27]&IN2[8];
  assign P36[25] = IN1[27]&IN2[9];
  assign P37[24] = IN1[27]&IN2[10];
  assign P38[23] = IN1[27]&IN2[11];
  assign P39[22] = IN1[27]&IN2[12];
  assign P40[21] = IN1[27]&IN2[13];
  assign P41[20] = IN1[27]&IN2[14];
  assign P42[19] = IN1[27]&IN2[15];
  assign P43[18] = IN1[27]&IN2[16];
  assign P44[17] = IN1[27]&IN2[17];
  assign P45[16] = IN1[27]&IN2[18];
  assign P46[15] = IN1[27]&IN2[19];
  assign P47[14] = IN1[27]&IN2[20];
  assign P48[13] = IN1[27]&IN2[21];
  assign P49[12] = IN1[27]&IN2[22];
  assign P50[11] = IN1[27]&IN2[23];
  assign P51[10] = IN1[27]&IN2[24];
  assign P52[9] = IN1[27]&IN2[25];
  assign P53[8] = IN1[27]&IN2[26];
  assign P54[7] = IN1[27]&IN2[27];
  assign P55[6] = IN1[27]&IN2[28];
  assign P56[5] = IN1[27]&IN2[29];
  assign P57[4] = IN1[27]&IN2[30];
  assign P58[3] = IN1[27]&IN2[31];
  assign P59[2] = IN1[27]&IN2[32];
  assign P60[1] = IN1[27]&IN2[33];
  assign P61[0] = IN1[27]&IN2[34];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[28] = IN1[28]&IN2[1];
  assign P30[28] = IN1[28]&IN2[2];
  assign P31[28] = IN1[28]&IN2[3];
  assign P32[28] = IN1[28]&IN2[4];
  assign P33[28] = IN1[28]&IN2[5];
  assign P34[28] = IN1[28]&IN2[6];
  assign P35[27] = IN1[28]&IN2[7];
  assign P36[26] = IN1[28]&IN2[8];
  assign P37[25] = IN1[28]&IN2[9];
  assign P38[24] = IN1[28]&IN2[10];
  assign P39[23] = IN1[28]&IN2[11];
  assign P40[22] = IN1[28]&IN2[12];
  assign P41[21] = IN1[28]&IN2[13];
  assign P42[20] = IN1[28]&IN2[14];
  assign P43[19] = IN1[28]&IN2[15];
  assign P44[18] = IN1[28]&IN2[16];
  assign P45[17] = IN1[28]&IN2[17];
  assign P46[16] = IN1[28]&IN2[18];
  assign P47[15] = IN1[28]&IN2[19];
  assign P48[14] = IN1[28]&IN2[20];
  assign P49[13] = IN1[28]&IN2[21];
  assign P50[12] = IN1[28]&IN2[22];
  assign P51[11] = IN1[28]&IN2[23];
  assign P52[10] = IN1[28]&IN2[24];
  assign P53[9] = IN1[28]&IN2[25];
  assign P54[8] = IN1[28]&IN2[26];
  assign P55[7] = IN1[28]&IN2[27];
  assign P56[6] = IN1[28]&IN2[28];
  assign P57[5] = IN1[28]&IN2[29];
  assign P58[4] = IN1[28]&IN2[30];
  assign P59[3] = IN1[28]&IN2[31];
  assign P60[2] = IN1[28]&IN2[32];
  assign P61[1] = IN1[28]&IN2[33];
  assign P62[0] = IN1[28]&IN2[34];
  assign P29[29] = IN1[29]&IN2[0];
  assign P30[29] = IN1[29]&IN2[1];
  assign P31[29] = IN1[29]&IN2[2];
  assign P32[29] = IN1[29]&IN2[3];
  assign P33[29] = IN1[29]&IN2[4];
  assign P34[29] = IN1[29]&IN2[5];
  assign P35[28] = IN1[29]&IN2[6];
  assign P36[27] = IN1[29]&IN2[7];
  assign P37[26] = IN1[29]&IN2[8];
  assign P38[25] = IN1[29]&IN2[9];
  assign P39[24] = IN1[29]&IN2[10];
  assign P40[23] = IN1[29]&IN2[11];
  assign P41[22] = IN1[29]&IN2[12];
  assign P42[21] = IN1[29]&IN2[13];
  assign P43[20] = IN1[29]&IN2[14];
  assign P44[19] = IN1[29]&IN2[15];
  assign P45[18] = IN1[29]&IN2[16];
  assign P46[17] = IN1[29]&IN2[17];
  assign P47[16] = IN1[29]&IN2[18];
  assign P48[15] = IN1[29]&IN2[19];
  assign P49[14] = IN1[29]&IN2[20];
  assign P50[13] = IN1[29]&IN2[21];
  assign P51[12] = IN1[29]&IN2[22];
  assign P52[11] = IN1[29]&IN2[23];
  assign P53[10] = IN1[29]&IN2[24];
  assign P54[9] = IN1[29]&IN2[25];
  assign P55[8] = IN1[29]&IN2[26];
  assign P56[7] = IN1[29]&IN2[27];
  assign P57[6] = IN1[29]&IN2[28];
  assign P58[5] = IN1[29]&IN2[29];
  assign P59[4] = IN1[29]&IN2[30];
  assign P60[3] = IN1[29]&IN2[31];
  assign P61[2] = IN1[29]&IN2[32];
  assign P62[1] = IN1[29]&IN2[33];
  assign P63[0] = IN1[29]&IN2[34];
  assign P30[30] = IN1[30]&IN2[0];
  assign P31[30] = IN1[30]&IN2[1];
  assign P32[30] = IN1[30]&IN2[2];
  assign P33[30] = IN1[30]&IN2[3];
  assign P34[30] = IN1[30]&IN2[4];
  assign P35[29] = IN1[30]&IN2[5];
  assign P36[28] = IN1[30]&IN2[6];
  assign P37[27] = IN1[30]&IN2[7];
  assign P38[26] = IN1[30]&IN2[8];
  assign P39[25] = IN1[30]&IN2[9];
  assign P40[24] = IN1[30]&IN2[10];
  assign P41[23] = IN1[30]&IN2[11];
  assign P42[22] = IN1[30]&IN2[12];
  assign P43[21] = IN1[30]&IN2[13];
  assign P44[20] = IN1[30]&IN2[14];
  assign P45[19] = IN1[30]&IN2[15];
  assign P46[18] = IN1[30]&IN2[16];
  assign P47[17] = IN1[30]&IN2[17];
  assign P48[16] = IN1[30]&IN2[18];
  assign P49[15] = IN1[30]&IN2[19];
  assign P50[14] = IN1[30]&IN2[20];
  assign P51[13] = IN1[30]&IN2[21];
  assign P52[12] = IN1[30]&IN2[22];
  assign P53[11] = IN1[30]&IN2[23];
  assign P54[10] = IN1[30]&IN2[24];
  assign P55[9] = IN1[30]&IN2[25];
  assign P56[8] = IN1[30]&IN2[26];
  assign P57[7] = IN1[30]&IN2[27];
  assign P58[6] = IN1[30]&IN2[28];
  assign P59[5] = IN1[30]&IN2[29];
  assign P60[4] = IN1[30]&IN2[30];
  assign P61[3] = IN1[30]&IN2[31];
  assign P62[2] = IN1[30]&IN2[32];
  assign P63[1] = IN1[30]&IN2[33];
  assign P64[0] = IN1[30]&IN2[34];
  assign P31[31] = IN1[31]&IN2[0];
  assign P32[31] = IN1[31]&IN2[1];
  assign P33[31] = IN1[31]&IN2[2];
  assign P34[31] = IN1[31]&IN2[3];
  assign P35[30] = IN1[31]&IN2[4];
  assign P36[29] = IN1[31]&IN2[5];
  assign P37[28] = IN1[31]&IN2[6];
  assign P38[27] = IN1[31]&IN2[7];
  assign P39[26] = IN1[31]&IN2[8];
  assign P40[25] = IN1[31]&IN2[9];
  assign P41[24] = IN1[31]&IN2[10];
  assign P42[23] = IN1[31]&IN2[11];
  assign P43[22] = IN1[31]&IN2[12];
  assign P44[21] = IN1[31]&IN2[13];
  assign P45[20] = IN1[31]&IN2[14];
  assign P46[19] = IN1[31]&IN2[15];
  assign P47[18] = IN1[31]&IN2[16];
  assign P48[17] = IN1[31]&IN2[17];
  assign P49[16] = IN1[31]&IN2[18];
  assign P50[15] = IN1[31]&IN2[19];
  assign P51[14] = IN1[31]&IN2[20];
  assign P52[13] = IN1[31]&IN2[21];
  assign P53[12] = IN1[31]&IN2[22];
  assign P54[11] = IN1[31]&IN2[23];
  assign P55[10] = IN1[31]&IN2[24];
  assign P56[9] = IN1[31]&IN2[25];
  assign P57[8] = IN1[31]&IN2[26];
  assign P58[7] = IN1[31]&IN2[27];
  assign P59[6] = IN1[31]&IN2[28];
  assign P60[5] = IN1[31]&IN2[29];
  assign P61[4] = IN1[31]&IN2[30];
  assign P62[3] = IN1[31]&IN2[31];
  assign P63[2] = IN1[31]&IN2[32];
  assign P64[1] = IN1[31]&IN2[33];
  assign P65[0] = IN1[31]&IN2[34];
  assign P32[32] = IN1[32]&IN2[0];
  assign P33[32] = IN1[32]&IN2[1];
  assign P34[32] = IN1[32]&IN2[2];
  assign P35[31] = IN1[32]&IN2[3];
  assign P36[30] = IN1[32]&IN2[4];
  assign P37[29] = IN1[32]&IN2[5];
  assign P38[28] = IN1[32]&IN2[6];
  assign P39[27] = IN1[32]&IN2[7];
  assign P40[26] = IN1[32]&IN2[8];
  assign P41[25] = IN1[32]&IN2[9];
  assign P42[24] = IN1[32]&IN2[10];
  assign P43[23] = IN1[32]&IN2[11];
  assign P44[22] = IN1[32]&IN2[12];
  assign P45[21] = IN1[32]&IN2[13];
  assign P46[20] = IN1[32]&IN2[14];
  assign P47[19] = IN1[32]&IN2[15];
  assign P48[18] = IN1[32]&IN2[16];
  assign P49[17] = IN1[32]&IN2[17];
  assign P50[16] = IN1[32]&IN2[18];
  assign P51[15] = IN1[32]&IN2[19];
  assign P52[14] = IN1[32]&IN2[20];
  assign P53[13] = IN1[32]&IN2[21];
  assign P54[12] = IN1[32]&IN2[22];
  assign P55[11] = IN1[32]&IN2[23];
  assign P56[10] = IN1[32]&IN2[24];
  assign P57[9] = IN1[32]&IN2[25];
  assign P58[8] = IN1[32]&IN2[26];
  assign P59[7] = IN1[32]&IN2[27];
  assign P60[6] = IN1[32]&IN2[28];
  assign P61[5] = IN1[32]&IN2[29];
  assign P62[4] = IN1[32]&IN2[30];
  assign P63[3] = IN1[32]&IN2[31];
  assign P64[2] = IN1[32]&IN2[32];
  assign P65[1] = IN1[32]&IN2[33];
  assign P66[0] = IN1[32]&IN2[34];
  assign P33[33] = IN1[33]&IN2[0];
  assign P34[33] = IN1[33]&IN2[1];
  assign P35[32] = IN1[33]&IN2[2];
  assign P36[31] = IN1[33]&IN2[3];
  assign P37[30] = IN1[33]&IN2[4];
  assign P38[29] = IN1[33]&IN2[5];
  assign P39[28] = IN1[33]&IN2[6];
  assign P40[27] = IN1[33]&IN2[7];
  assign P41[26] = IN1[33]&IN2[8];
  assign P42[25] = IN1[33]&IN2[9];
  assign P43[24] = IN1[33]&IN2[10];
  assign P44[23] = IN1[33]&IN2[11];
  assign P45[22] = IN1[33]&IN2[12];
  assign P46[21] = IN1[33]&IN2[13];
  assign P47[20] = IN1[33]&IN2[14];
  assign P48[19] = IN1[33]&IN2[15];
  assign P49[18] = IN1[33]&IN2[16];
  assign P50[17] = IN1[33]&IN2[17];
  assign P51[16] = IN1[33]&IN2[18];
  assign P52[15] = IN1[33]&IN2[19];
  assign P53[14] = IN1[33]&IN2[20];
  assign P54[13] = IN1[33]&IN2[21];
  assign P55[12] = IN1[33]&IN2[22];
  assign P56[11] = IN1[33]&IN2[23];
  assign P57[10] = IN1[33]&IN2[24];
  assign P58[9] = IN1[33]&IN2[25];
  assign P59[8] = IN1[33]&IN2[26];
  assign P60[7] = IN1[33]&IN2[27];
  assign P61[6] = IN1[33]&IN2[28];
  assign P62[5] = IN1[33]&IN2[29];
  assign P63[4] = IN1[33]&IN2[30];
  assign P64[3] = IN1[33]&IN2[31];
  assign P65[2] = IN1[33]&IN2[32];
  assign P66[1] = IN1[33]&IN2[33];
  assign P67[0] = IN1[33]&IN2[34];
  assign P34[34] = IN1[34]&IN2[0];
  assign P35[33] = IN1[34]&IN2[1];
  assign P36[32] = IN1[34]&IN2[2];
  assign P37[31] = IN1[34]&IN2[3];
  assign P38[30] = IN1[34]&IN2[4];
  assign P39[29] = IN1[34]&IN2[5];
  assign P40[28] = IN1[34]&IN2[6];
  assign P41[27] = IN1[34]&IN2[7];
  assign P42[26] = IN1[34]&IN2[8];
  assign P43[25] = IN1[34]&IN2[9];
  assign P44[24] = IN1[34]&IN2[10];
  assign P45[23] = IN1[34]&IN2[11];
  assign P46[22] = IN1[34]&IN2[12];
  assign P47[21] = IN1[34]&IN2[13];
  assign P48[20] = IN1[34]&IN2[14];
  assign P49[19] = IN1[34]&IN2[15];
  assign P50[18] = IN1[34]&IN2[16];
  assign P51[17] = IN1[34]&IN2[17];
  assign P52[16] = IN1[34]&IN2[18];
  assign P53[15] = IN1[34]&IN2[19];
  assign P54[14] = IN1[34]&IN2[20];
  assign P55[13] = IN1[34]&IN2[21];
  assign P56[12] = IN1[34]&IN2[22];
  assign P57[11] = IN1[34]&IN2[23];
  assign P58[10] = IN1[34]&IN2[24];
  assign P59[9] = IN1[34]&IN2[25];
  assign P60[8] = IN1[34]&IN2[26];
  assign P61[7] = IN1[34]&IN2[27];
  assign P62[6] = IN1[34]&IN2[28];
  assign P63[5] = IN1[34]&IN2[29];
  assign P64[4] = IN1[34]&IN2[30];
  assign P65[3] = IN1[34]&IN2[31];
  assign P66[2] = IN1[34]&IN2[32];
  assign P67[1] = IN1[34]&IN2[33];
  assign P68[0] = IN1[34]&IN2[34];
  assign P35[34] = IN1[35]&IN2[0];
  assign P36[33] = IN1[35]&IN2[1];
  assign P37[32] = IN1[35]&IN2[2];
  assign P38[31] = IN1[35]&IN2[3];
  assign P39[30] = IN1[35]&IN2[4];
  assign P40[29] = IN1[35]&IN2[5];
  assign P41[28] = IN1[35]&IN2[6];
  assign P42[27] = IN1[35]&IN2[7];
  assign P43[26] = IN1[35]&IN2[8];
  assign P44[25] = IN1[35]&IN2[9];
  assign P45[24] = IN1[35]&IN2[10];
  assign P46[23] = IN1[35]&IN2[11];
  assign P47[22] = IN1[35]&IN2[12];
  assign P48[21] = IN1[35]&IN2[13];
  assign P49[20] = IN1[35]&IN2[14];
  assign P50[19] = IN1[35]&IN2[15];
  assign P51[18] = IN1[35]&IN2[16];
  assign P52[17] = IN1[35]&IN2[17];
  assign P53[16] = IN1[35]&IN2[18];
  assign P54[15] = IN1[35]&IN2[19];
  assign P55[14] = IN1[35]&IN2[20];
  assign P56[13] = IN1[35]&IN2[21];
  assign P57[12] = IN1[35]&IN2[22];
  assign P58[11] = IN1[35]&IN2[23];
  assign P59[10] = IN1[35]&IN2[24];
  assign P60[9] = IN1[35]&IN2[25];
  assign P61[8] = IN1[35]&IN2[26];
  assign P62[7] = IN1[35]&IN2[27];
  assign P63[6] = IN1[35]&IN2[28];
  assign P64[5] = IN1[35]&IN2[29];
  assign P65[4] = IN1[35]&IN2[30];
  assign P66[3] = IN1[35]&IN2[31];
  assign P67[2] = IN1[35]&IN2[32];
  assign P68[1] = IN1[35]&IN2[33];
  assign P69[0] = IN1[35]&IN2[34];
  assign P36[34] = IN1[36]&IN2[0];
  assign P37[33] = IN1[36]&IN2[1];
  assign P38[32] = IN1[36]&IN2[2];
  assign P39[31] = IN1[36]&IN2[3];
  assign P40[30] = IN1[36]&IN2[4];
  assign P41[29] = IN1[36]&IN2[5];
  assign P42[28] = IN1[36]&IN2[6];
  assign P43[27] = IN1[36]&IN2[7];
  assign P44[26] = IN1[36]&IN2[8];
  assign P45[25] = IN1[36]&IN2[9];
  assign P46[24] = IN1[36]&IN2[10];
  assign P47[23] = IN1[36]&IN2[11];
  assign P48[22] = IN1[36]&IN2[12];
  assign P49[21] = IN1[36]&IN2[13];
  assign P50[20] = IN1[36]&IN2[14];
  assign P51[19] = IN1[36]&IN2[15];
  assign P52[18] = IN1[36]&IN2[16];
  assign P53[17] = IN1[36]&IN2[17];
  assign P54[16] = IN1[36]&IN2[18];
  assign P55[15] = IN1[36]&IN2[19];
  assign P56[14] = IN1[36]&IN2[20];
  assign P57[13] = IN1[36]&IN2[21];
  assign P58[12] = IN1[36]&IN2[22];
  assign P59[11] = IN1[36]&IN2[23];
  assign P60[10] = IN1[36]&IN2[24];
  assign P61[9] = IN1[36]&IN2[25];
  assign P62[8] = IN1[36]&IN2[26];
  assign P63[7] = IN1[36]&IN2[27];
  assign P64[6] = IN1[36]&IN2[28];
  assign P65[5] = IN1[36]&IN2[29];
  assign P66[4] = IN1[36]&IN2[30];
  assign P67[3] = IN1[36]&IN2[31];
  assign P68[2] = IN1[36]&IN2[32];
  assign P69[1] = IN1[36]&IN2[33];
  assign P70[0] = IN1[36]&IN2[34];
  assign P37[34] = IN1[37]&IN2[0];
  assign P38[33] = IN1[37]&IN2[1];
  assign P39[32] = IN1[37]&IN2[2];
  assign P40[31] = IN1[37]&IN2[3];
  assign P41[30] = IN1[37]&IN2[4];
  assign P42[29] = IN1[37]&IN2[5];
  assign P43[28] = IN1[37]&IN2[6];
  assign P44[27] = IN1[37]&IN2[7];
  assign P45[26] = IN1[37]&IN2[8];
  assign P46[25] = IN1[37]&IN2[9];
  assign P47[24] = IN1[37]&IN2[10];
  assign P48[23] = IN1[37]&IN2[11];
  assign P49[22] = IN1[37]&IN2[12];
  assign P50[21] = IN1[37]&IN2[13];
  assign P51[20] = IN1[37]&IN2[14];
  assign P52[19] = IN1[37]&IN2[15];
  assign P53[18] = IN1[37]&IN2[16];
  assign P54[17] = IN1[37]&IN2[17];
  assign P55[16] = IN1[37]&IN2[18];
  assign P56[15] = IN1[37]&IN2[19];
  assign P57[14] = IN1[37]&IN2[20];
  assign P58[13] = IN1[37]&IN2[21];
  assign P59[12] = IN1[37]&IN2[22];
  assign P60[11] = IN1[37]&IN2[23];
  assign P61[10] = IN1[37]&IN2[24];
  assign P62[9] = IN1[37]&IN2[25];
  assign P63[8] = IN1[37]&IN2[26];
  assign P64[7] = IN1[37]&IN2[27];
  assign P65[6] = IN1[37]&IN2[28];
  assign P66[5] = IN1[37]&IN2[29];
  assign P67[4] = IN1[37]&IN2[30];
  assign P68[3] = IN1[37]&IN2[31];
  assign P69[2] = IN1[37]&IN2[32];
  assign P70[1] = IN1[37]&IN2[33];
  assign P71[0] = IN1[37]&IN2[34];
  assign P38[34] = IN1[38]&IN2[0];
  assign P39[33] = IN1[38]&IN2[1];
  assign P40[32] = IN1[38]&IN2[2];
  assign P41[31] = IN1[38]&IN2[3];
  assign P42[30] = IN1[38]&IN2[4];
  assign P43[29] = IN1[38]&IN2[5];
  assign P44[28] = IN1[38]&IN2[6];
  assign P45[27] = IN1[38]&IN2[7];
  assign P46[26] = IN1[38]&IN2[8];
  assign P47[25] = IN1[38]&IN2[9];
  assign P48[24] = IN1[38]&IN2[10];
  assign P49[23] = IN1[38]&IN2[11];
  assign P50[22] = IN1[38]&IN2[12];
  assign P51[21] = IN1[38]&IN2[13];
  assign P52[20] = IN1[38]&IN2[14];
  assign P53[19] = IN1[38]&IN2[15];
  assign P54[18] = IN1[38]&IN2[16];
  assign P55[17] = IN1[38]&IN2[17];
  assign P56[16] = IN1[38]&IN2[18];
  assign P57[15] = IN1[38]&IN2[19];
  assign P58[14] = IN1[38]&IN2[20];
  assign P59[13] = IN1[38]&IN2[21];
  assign P60[12] = IN1[38]&IN2[22];
  assign P61[11] = IN1[38]&IN2[23];
  assign P62[10] = IN1[38]&IN2[24];
  assign P63[9] = IN1[38]&IN2[25];
  assign P64[8] = IN1[38]&IN2[26];
  assign P65[7] = IN1[38]&IN2[27];
  assign P66[6] = IN1[38]&IN2[28];
  assign P67[5] = IN1[38]&IN2[29];
  assign P68[4] = IN1[38]&IN2[30];
  assign P69[3] = IN1[38]&IN2[31];
  assign P70[2] = IN1[38]&IN2[32];
  assign P71[1] = IN1[38]&IN2[33];
  assign P72[0] = IN1[38]&IN2[34];
  assign P39[34] = IN1[39]&IN2[0];
  assign P40[33] = IN1[39]&IN2[1];
  assign P41[32] = IN1[39]&IN2[2];
  assign P42[31] = IN1[39]&IN2[3];
  assign P43[30] = IN1[39]&IN2[4];
  assign P44[29] = IN1[39]&IN2[5];
  assign P45[28] = IN1[39]&IN2[6];
  assign P46[27] = IN1[39]&IN2[7];
  assign P47[26] = IN1[39]&IN2[8];
  assign P48[25] = IN1[39]&IN2[9];
  assign P49[24] = IN1[39]&IN2[10];
  assign P50[23] = IN1[39]&IN2[11];
  assign P51[22] = IN1[39]&IN2[12];
  assign P52[21] = IN1[39]&IN2[13];
  assign P53[20] = IN1[39]&IN2[14];
  assign P54[19] = IN1[39]&IN2[15];
  assign P55[18] = IN1[39]&IN2[16];
  assign P56[17] = IN1[39]&IN2[17];
  assign P57[16] = IN1[39]&IN2[18];
  assign P58[15] = IN1[39]&IN2[19];
  assign P59[14] = IN1[39]&IN2[20];
  assign P60[13] = IN1[39]&IN2[21];
  assign P61[12] = IN1[39]&IN2[22];
  assign P62[11] = IN1[39]&IN2[23];
  assign P63[10] = IN1[39]&IN2[24];
  assign P64[9] = IN1[39]&IN2[25];
  assign P65[8] = IN1[39]&IN2[26];
  assign P66[7] = IN1[39]&IN2[27];
  assign P67[6] = IN1[39]&IN2[28];
  assign P68[5] = IN1[39]&IN2[29];
  assign P69[4] = IN1[39]&IN2[30];
  assign P70[3] = IN1[39]&IN2[31];
  assign P71[2] = IN1[39]&IN2[32];
  assign P72[1] = IN1[39]&IN2[33];
  assign P73[0] = IN1[39]&IN2[34];
  assign P40[34] = IN1[40]&IN2[0];
  assign P41[33] = IN1[40]&IN2[1];
  assign P42[32] = IN1[40]&IN2[2];
  assign P43[31] = IN1[40]&IN2[3];
  assign P44[30] = IN1[40]&IN2[4];
  assign P45[29] = IN1[40]&IN2[5];
  assign P46[28] = IN1[40]&IN2[6];
  assign P47[27] = IN1[40]&IN2[7];
  assign P48[26] = IN1[40]&IN2[8];
  assign P49[25] = IN1[40]&IN2[9];
  assign P50[24] = IN1[40]&IN2[10];
  assign P51[23] = IN1[40]&IN2[11];
  assign P52[22] = IN1[40]&IN2[12];
  assign P53[21] = IN1[40]&IN2[13];
  assign P54[20] = IN1[40]&IN2[14];
  assign P55[19] = IN1[40]&IN2[15];
  assign P56[18] = IN1[40]&IN2[16];
  assign P57[17] = IN1[40]&IN2[17];
  assign P58[16] = IN1[40]&IN2[18];
  assign P59[15] = IN1[40]&IN2[19];
  assign P60[14] = IN1[40]&IN2[20];
  assign P61[13] = IN1[40]&IN2[21];
  assign P62[12] = IN1[40]&IN2[22];
  assign P63[11] = IN1[40]&IN2[23];
  assign P64[10] = IN1[40]&IN2[24];
  assign P65[9] = IN1[40]&IN2[25];
  assign P66[8] = IN1[40]&IN2[26];
  assign P67[7] = IN1[40]&IN2[27];
  assign P68[6] = IN1[40]&IN2[28];
  assign P69[5] = IN1[40]&IN2[29];
  assign P70[4] = IN1[40]&IN2[30];
  assign P71[3] = IN1[40]&IN2[31];
  assign P72[2] = IN1[40]&IN2[32];
  assign P73[1] = IN1[40]&IN2[33];
  assign P74[0] = IN1[40]&IN2[34];
  assign P41[34] = IN1[41]&IN2[0];
  assign P42[33] = IN1[41]&IN2[1];
  assign P43[32] = IN1[41]&IN2[2];
  assign P44[31] = IN1[41]&IN2[3];
  assign P45[30] = IN1[41]&IN2[4];
  assign P46[29] = IN1[41]&IN2[5];
  assign P47[28] = IN1[41]&IN2[6];
  assign P48[27] = IN1[41]&IN2[7];
  assign P49[26] = IN1[41]&IN2[8];
  assign P50[25] = IN1[41]&IN2[9];
  assign P51[24] = IN1[41]&IN2[10];
  assign P52[23] = IN1[41]&IN2[11];
  assign P53[22] = IN1[41]&IN2[12];
  assign P54[21] = IN1[41]&IN2[13];
  assign P55[20] = IN1[41]&IN2[14];
  assign P56[19] = IN1[41]&IN2[15];
  assign P57[18] = IN1[41]&IN2[16];
  assign P58[17] = IN1[41]&IN2[17];
  assign P59[16] = IN1[41]&IN2[18];
  assign P60[15] = IN1[41]&IN2[19];
  assign P61[14] = IN1[41]&IN2[20];
  assign P62[13] = IN1[41]&IN2[21];
  assign P63[12] = IN1[41]&IN2[22];
  assign P64[11] = IN1[41]&IN2[23];
  assign P65[10] = IN1[41]&IN2[24];
  assign P66[9] = IN1[41]&IN2[25];
  assign P67[8] = IN1[41]&IN2[26];
  assign P68[7] = IN1[41]&IN2[27];
  assign P69[6] = IN1[41]&IN2[28];
  assign P70[5] = IN1[41]&IN2[29];
  assign P71[4] = IN1[41]&IN2[30];
  assign P72[3] = IN1[41]&IN2[31];
  assign P73[2] = IN1[41]&IN2[32];
  assign P74[1] = IN1[41]&IN2[33];
  assign P75[0] = IN1[41]&IN2[34];
  assign P42[34] = IN1[42]&IN2[0];
  assign P43[33] = IN1[42]&IN2[1];
  assign P44[32] = IN1[42]&IN2[2];
  assign P45[31] = IN1[42]&IN2[3];
  assign P46[30] = IN1[42]&IN2[4];
  assign P47[29] = IN1[42]&IN2[5];
  assign P48[28] = IN1[42]&IN2[6];
  assign P49[27] = IN1[42]&IN2[7];
  assign P50[26] = IN1[42]&IN2[8];
  assign P51[25] = IN1[42]&IN2[9];
  assign P52[24] = IN1[42]&IN2[10];
  assign P53[23] = IN1[42]&IN2[11];
  assign P54[22] = IN1[42]&IN2[12];
  assign P55[21] = IN1[42]&IN2[13];
  assign P56[20] = IN1[42]&IN2[14];
  assign P57[19] = IN1[42]&IN2[15];
  assign P58[18] = IN1[42]&IN2[16];
  assign P59[17] = IN1[42]&IN2[17];
  assign P60[16] = IN1[42]&IN2[18];
  assign P61[15] = IN1[42]&IN2[19];
  assign P62[14] = IN1[42]&IN2[20];
  assign P63[13] = IN1[42]&IN2[21];
  assign P64[12] = IN1[42]&IN2[22];
  assign P65[11] = IN1[42]&IN2[23];
  assign P66[10] = IN1[42]&IN2[24];
  assign P67[9] = IN1[42]&IN2[25];
  assign P68[8] = IN1[42]&IN2[26];
  assign P69[7] = IN1[42]&IN2[27];
  assign P70[6] = IN1[42]&IN2[28];
  assign P71[5] = IN1[42]&IN2[29];
  assign P72[4] = IN1[42]&IN2[30];
  assign P73[3] = IN1[42]&IN2[31];
  assign P74[2] = IN1[42]&IN2[32];
  assign P75[1] = IN1[42]&IN2[33];
  assign P76[0] = IN1[42]&IN2[34];
  assign P43[34] = IN1[43]&IN2[0];
  assign P44[33] = IN1[43]&IN2[1];
  assign P45[32] = IN1[43]&IN2[2];
  assign P46[31] = IN1[43]&IN2[3];
  assign P47[30] = IN1[43]&IN2[4];
  assign P48[29] = IN1[43]&IN2[5];
  assign P49[28] = IN1[43]&IN2[6];
  assign P50[27] = IN1[43]&IN2[7];
  assign P51[26] = IN1[43]&IN2[8];
  assign P52[25] = IN1[43]&IN2[9];
  assign P53[24] = IN1[43]&IN2[10];
  assign P54[23] = IN1[43]&IN2[11];
  assign P55[22] = IN1[43]&IN2[12];
  assign P56[21] = IN1[43]&IN2[13];
  assign P57[20] = IN1[43]&IN2[14];
  assign P58[19] = IN1[43]&IN2[15];
  assign P59[18] = IN1[43]&IN2[16];
  assign P60[17] = IN1[43]&IN2[17];
  assign P61[16] = IN1[43]&IN2[18];
  assign P62[15] = IN1[43]&IN2[19];
  assign P63[14] = IN1[43]&IN2[20];
  assign P64[13] = IN1[43]&IN2[21];
  assign P65[12] = IN1[43]&IN2[22];
  assign P66[11] = IN1[43]&IN2[23];
  assign P67[10] = IN1[43]&IN2[24];
  assign P68[9] = IN1[43]&IN2[25];
  assign P69[8] = IN1[43]&IN2[26];
  assign P70[7] = IN1[43]&IN2[27];
  assign P71[6] = IN1[43]&IN2[28];
  assign P72[5] = IN1[43]&IN2[29];
  assign P73[4] = IN1[43]&IN2[30];
  assign P74[3] = IN1[43]&IN2[31];
  assign P75[2] = IN1[43]&IN2[32];
  assign P76[1] = IN1[43]&IN2[33];
  assign P77[0] = IN1[43]&IN2[34];
  assign P44[34] = IN1[44]&IN2[0];
  assign P45[33] = IN1[44]&IN2[1];
  assign P46[32] = IN1[44]&IN2[2];
  assign P47[31] = IN1[44]&IN2[3];
  assign P48[30] = IN1[44]&IN2[4];
  assign P49[29] = IN1[44]&IN2[5];
  assign P50[28] = IN1[44]&IN2[6];
  assign P51[27] = IN1[44]&IN2[7];
  assign P52[26] = IN1[44]&IN2[8];
  assign P53[25] = IN1[44]&IN2[9];
  assign P54[24] = IN1[44]&IN2[10];
  assign P55[23] = IN1[44]&IN2[11];
  assign P56[22] = IN1[44]&IN2[12];
  assign P57[21] = IN1[44]&IN2[13];
  assign P58[20] = IN1[44]&IN2[14];
  assign P59[19] = IN1[44]&IN2[15];
  assign P60[18] = IN1[44]&IN2[16];
  assign P61[17] = IN1[44]&IN2[17];
  assign P62[16] = IN1[44]&IN2[18];
  assign P63[15] = IN1[44]&IN2[19];
  assign P64[14] = IN1[44]&IN2[20];
  assign P65[13] = IN1[44]&IN2[21];
  assign P66[12] = IN1[44]&IN2[22];
  assign P67[11] = IN1[44]&IN2[23];
  assign P68[10] = IN1[44]&IN2[24];
  assign P69[9] = IN1[44]&IN2[25];
  assign P70[8] = IN1[44]&IN2[26];
  assign P71[7] = IN1[44]&IN2[27];
  assign P72[6] = IN1[44]&IN2[28];
  assign P73[5] = IN1[44]&IN2[29];
  assign P74[4] = IN1[44]&IN2[30];
  assign P75[3] = IN1[44]&IN2[31];
  assign P76[2] = IN1[44]&IN2[32];
  assign P77[1] = IN1[44]&IN2[33];
  assign P78[0] = IN1[44]&IN2[34];
  assign P45[34] = IN1[45]&IN2[0];
  assign P46[33] = IN1[45]&IN2[1];
  assign P47[32] = IN1[45]&IN2[2];
  assign P48[31] = IN1[45]&IN2[3];
  assign P49[30] = IN1[45]&IN2[4];
  assign P50[29] = IN1[45]&IN2[5];
  assign P51[28] = IN1[45]&IN2[6];
  assign P52[27] = IN1[45]&IN2[7];
  assign P53[26] = IN1[45]&IN2[8];
  assign P54[25] = IN1[45]&IN2[9];
  assign P55[24] = IN1[45]&IN2[10];
  assign P56[23] = IN1[45]&IN2[11];
  assign P57[22] = IN1[45]&IN2[12];
  assign P58[21] = IN1[45]&IN2[13];
  assign P59[20] = IN1[45]&IN2[14];
  assign P60[19] = IN1[45]&IN2[15];
  assign P61[18] = IN1[45]&IN2[16];
  assign P62[17] = IN1[45]&IN2[17];
  assign P63[16] = IN1[45]&IN2[18];
  assign P64[15] = IN1[45]&IN2[19];
  assign P65[14] = IN1[45]&IN2[20];
  assign P66[13] = IN1[45]&IN2[21];
  assign P67[12] = IN1[45]&IN2[22];
  assign P68[11] = IN1[45]&IN2[23];
  assign P69[10] = IN1[45]&IN2[24];
  assign P70[9] = IN1[45]&IN2[25];
  assign P71[8] = IN1[45]&IN2[26];
  assign P72[7] = IN1[45]&IN2[27];
  assign P73[6] = IN1[45]&IN2[28];
  assign P74[5] = IN1[45]&IN2[29];
  assign P75[4] = IN1[45]&IN2[30];
  assign P76[3] = IN1[45]&IN2[31];
  assign P77[2] = IN1[45]&IN2[32];
  assign P78[1] = IN1[45]&IN2[33];
  assign P79[0] = IN1[45]&IN2[34];
  assign P46[34] = IN1[46]&IN2[0];
  assign P47[33] = IN1[46]&IN2[1];
  assign P48[32] = IN1[46]&IN2[2];
  assign P49[31] = IN1[46]&IN2[3];
  assign P50[30] = IN1[46]&IN2[4];
  assign P51[29] = IN1[46]&IN2[5];
  assign P52[28] = IN1[46]&IN2[6];
  assign P53[27] = IN1[46]&IN2[7];
  assign P54[26] = IN1[46]&IN2[8];
  assign P55[25] = IN1[46]&IN2[9];
  assign P56[24] = IN1[46]&IN2[10];
  assign P57[23] = IN1[46]&IN2[11];
  assign P58[22] = IN1[46]&IN2[12];
  assign P59[21] = IN1[46]&IN2[13];
  assign P60[20] = IN1[46]&IN2[14];
  assign P61[19] = IN1[46]&IN2[15];
  assign P62[18] = IN1[46]&IN2[16];
  assign P63[17] = IN1[46]&IN2[17];
  assign P64[16] = IN1[46]&IN2[18];
  assign P65[15] = IN1[46]&IN2[19];
  assign P66[14] = IN1[46]&IN2[20];
  assign P67[13] = IN1[46]&IN2[21];
  assign P68[12] = IN1[46]&IN2[22];
  assign P69[11] = IN1[46]&IN2[23];
  assign P70[10] = IN1[46]&IN2[24];
  assign P71[9] = IN1[46]&IN2[25];
  assign P72[8] = IN1[46]&IN2[26];
  assign P73[7] = IN1[46]&IN2[27];
  assign P74[6] = IN1[46]&IN2[28];
  assign P75[5] = IN1[46]&IN2[29];
  assign P76[4] = IN1[46]&IN2[30];
  assign P77[3] = IN1[46]&IN2[31];
  assign P78[2] = IN1[46]&IN2[32];
  assign P79[1] = IN1[46]&IN2[33];
  assign P80[0] = IN1[46]&IN2[34];
  assign P47[34] = IN1[47]&IN2[0];
  assign P48[33] = IN1[47]&IN2[1];
  assign P49[32] = IN1[47]&IN2[2];
  assign P50[31] = IN1[47]&IN2[3];
  assign P51[30] = IN1[47]&IN2[4];
  assign P52[29] = IN1[47]&IN2[5];
  assign P53[28] = IN1[47]&IN2[6];
  assign P54[27] = IN1[47]&IN2[7];
  assign P55[26] = IN1[47]&IN2[8];
  assign P56[25] = IN1[47]&IN2[9];
  assign P57[24] = IN1[47]&IN2[10];
  assign P58[23] = IN1[47]&IN2[11];
  assign P59[22] = IN1[47]&IN2[12];
  assign P60[21] = IN1[47]&IN2[13];
  assign P61[20] = IN1[47]&IN2[14];
  assign P62[19] = IN1[47]&IN2[15];
  assign P63[18] = IN1[47]&IN2[16];
  assign P64[17] = IN1[47]&IN2[17];
  assign P65[16] = IN1[47]&IN2[18];
  assign P66[15] = IN1[47]&IN2[19];
  assign P67[14] = IN1[47]&IN2[20];
  assign P68[13] = IN1[47]&IN2[21];
  assign P69[12] = IN1[47]&IN2[22];
  assign P70[11] = IN1[47]&IN2[23];
  assign P71[10] = IN1[47]&IN2[24];
  assign P72[9] = IN1[47]&IN2[25];
  assign P73[8] = IN1[47]&IN2[26];
  assign P74[7] = IN1[47]&IN2[27];
  assign P75[6] = IN1[47]&IN2[28];
  assign P76[5] = IN1[47]&IN2[29];
  assign P77[4] = IN1[47]&IN2[30];
  assign P78[3] = IN1[47]&IN2[31];
  assign P79[2] = IN1[47]&IN2[32];
  assign P80[1] = IN1[47]&IN2[33];
  assign P81[0] = IN1[47]&IN2[34];
  assign P48[34] = IN1[48]&IN2[0];
  assign P49[33] = IN1[48]&IN2[1];
  assign P50[32] = IN1[48]&IN2[2];
  assign P51[31] = IN1[48]&IN2[3];
  assign P52[30] = IN1[48]&IN2[4];
  assign P53[29] = IN1[48]&IN2[5];
  assign P54[28] = IN1[48]&IN2[6];
  assign P55[27] = IN1[48]&IN2[7];
  assign P56[26] = IN1[48]&IN2[8];
  assign P57[25] = IN1[48]&IN2[9];
  assign P58[24] = IN1[48]&IN2[10];
  assign P59[23] = IN1[48]&IN2[11];
  assign P60[22] = IN1[48]&IN2[12];
  assign P61[21] = IN1[48]&IN2[13];
  assign P62[20] = IN1[48]&IN2[14];
  assign P63[19] = IN1[48]&IN2[15];
  assign P64[18] = IN1[48]&IN2[16];
  assign P65[17] = IN1[48]&IN2[17];
  assign P66[16] = IN1[48]&IN2[18];
  assign P67[15] = IN1[48]&IN2[19];
  assign P68[14] = IN1[48]&IN2[20];
  assign P69[13] = IN1[48]&IN2[21];
  assign P70[12] = IN1[48]&IN2[22];
  assign P71[11] = IN1[48]&IN2[23];
  assign P72[10] = IN1[48]&IN2[24];
  assign P73[9] = IN1[48]&IN2[25];
  assign P74[8] = IN1[48]&IN2[26];
  assign P75[7] = IN1[48]&IN2[27];
  assign P76[6] = IN1[48]&IN2[28];
  assign P77[5] = IN1[48]&IN2[29];
  assign P78[4] = IN1[48]&IN2[30];
  assign P79[3] = IN1[48]&IN2[31];
  assign P80[2] = IN1[48]&IN2[32];
  assign P81[1] = IN1[48]&IN2[33];
  assign P82[0] = IN1[48]&IN2[34];
  assign P49[34] = IN1[49]&IN2[0];
  assign P50[33] = IN1[49]&IN2[1];
  assign P51[32] = IN1[49]&IN2[2];
  assign P52[31] = IN1[49]&IN2[3];
  assign P53[30] = IN1[49]&IN2[4];
  assign P54[29] = IN1[49]&IN2[5];
  assign P55[28] = IN1[49]&IN2[6];
  assign P56[27] = IN1[49]&IN2[7];
  assign P57[26] = IN1[49]&IN2[8];
  assign P58[25] = IN1[49]&IN2[9];
  assign P59[24] = IN1[49]&IN2[10];
  assign P60[23] = IN1[49]&IN2[11];
  assign P61[22] = IN1[49]&IN2[12];
  assign P62[21] = IN1[49]&IN2[13];
  assign P63[20] = IN1[49]&IN2[14];
  assign P64[19] = IN1[49]&IN2[15];
  assign P65[18] = IN1[49]&IN2[16];
  assign P66[17] = IN1[49]&IN2[17];
  assign P67[16] = IN1[49]&IN2[18];
  assign P68[15] = IN1[49]&IN2[19];
  assign P69[14] = IN1[49]&IN2[20];
  assign P70[13] = IN1[49]&IN2[21];
  assign P71[12] = IN1[49]&IN2[22];
  assign P72[11] = IN1[49]&IN2[23];
  assign P73[10] = IN1[49]&IN2[24];
  assign P74[9] = IN1[49]&IN2[25];
  assign P75[8] = IN1[49]&IN2[26];
  assign P76[7] = IN1[49]&IN2[27];
  assign P77[6] = IN1[49]&IN2[28];
  assign P78[5] = IN1[49]&IN2[29];
  assign P79[4] = IN1[49]&IN2[30];
  assign P80[3] = IN1[49]&IN2[31];
  assign P81[2] = IN1[49]&IN2[32];
  assign P82[1] = IN1[49]&IN2[33];
  assign P83[0] = IN1[49]&IN2[34];
  assign P50[34] = IN1[50]&IN2[0];
  assign P51[33] = IN1[50]&IN2[1];
  assign P52[32] = IN1[50]&IN2[2];
  assign P53[31] = IN1[50]&IN2[3];
  assign P54[30] = IN1[50]&IN2[4];
  assign P55[29] = IN1[50]&IN2[5];
  assign P56[28] = IN1[50]&IN2[6];
  assign P57[27] = IN1[50]&IN2[7];
  assign P58[26] = IN1[50]&IN2[8];
  assign P59[25] = IN1[50]&IN2[9];
  assign P60[24] = IN1[50]&IN2[10];
  assign P61[23] = IN1[50]&IN2[11];
  assign P62[22] = IN1[50]&IN2[12];
  assign P63[21] = IN1[50]&IN2[13];
  assign P64[20] = IN1[50]&IN2[14];
  assign P65[19] = IN1[50]&IN2[15];
  assign P66[18] = IN1[50]&IN2[16];
  assign P67[17] = IN1[50]&IN2[17];
  assign P68[16] = IN1[50]&IN2[18];
  assign P69[15] = IN1[50]&IN2[19];
  assign P70[14] = IN1[50]&IN2[20];
  assign P71[13] = IN1[50]&IN2[21];
  assign P72[12] = IN1[50]&IN2[22];
  assign P73[11] = IN1[50]&IN2[23];
  assign P74[10] = IN1[50]&IN2[24];
  assign P75[9] = IN1[50]&IN2[25];
  assign P76[8] = IN1[50]&IN2[26];
  assign P77[7] = IN1[50]&IN2[27];
  assign P78[6] = IN1[50]&IN2[28];
  assign P79[5] = IN1[50]&IN2[29];
  assign P80[4] = IN1[50]&IN2[30];
  assign P81[3] = IN1[50]&IN2[31];
  assign P82[2] = IN1[50]&IN2[32];
  assign P83[1] = IN1[50]&IN2[33];
  assign P84[0] = IN1[50]&IN2[34];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, IN79, IN80, IN81, IN82, IN83, IN84, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [29:0] IN29;
  input [30:0] IN30;
  input [31:0] IN31;
  input [32:0] IN32;
  input [33:0] IN33;
  input [34:0] IN34;
  input [34:0] IN35;
  input [34:0] IN36;
  input [34:0] IN37;
  input [34:0] IN38;
  input [34:0] IN39;
  input [34:0] IN40;
  input [34:0] IN41;
  input [34:0] IN42;
  input [34:0] IN43;
  input [34:0] IN44;
  input [34:0] IN45;
  input [34:0] IN46;
  input [34:0] IN47;
  input [34:0] IN48;
  input [34:0] IN49;
  input [34:0] IN50;
  input [33:0] IN51;
  input [32:0] IN52;
  input [31:0] IN53;
  input [30:0] IN54;
  input [29:0] IN55;
  input [28:0] IN56;
  input [27:0] IN57;
  input [26:0] IN58;
  input [25:0] IN59;
  input [24:0] IN60;
  input [23:0] IN61;
  input [22:0] IN62;
  input [21:0] IN63;
  input [20:0] IN64;
  input [19:0] IN65;
  input [18:0] IN66;
  input [17:0] IN67;
  input [16:0] IN68;
  input [15:0] IN69;
  input [14:0] IN70;
  input [13:0] IN71;
  input [12:0] IN72;
  input [11:0] IN73;
  input [10:0] IN74;
  input [9:0] IN75;
  input [8:0] IN76;
  input [7:0] IN77;
  input [6:0] IN78;
  input [5:0] IN79;
  input [4:0] IN80;
  input [3:0] IN81;
  input [2:0] IN82;
  input [1:0] IN83;
  input [0:0] IN84;
  output [84:0] Out1;
  output [33:0] Out2;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1984;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2050;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2086;
  wire w2087;
  wire w2088;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2140;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2586;
  wire w2587;
  wire w2588;
  wire w2589;
  wire w2590;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2614;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2631;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2638;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2680;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2686;
  wire w2687;
  wire w2688;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2694;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2708;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2738;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2747;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2770;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2774;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2786;
  wire w2787;
  wire w2788;
  wire w2789;
  wire w2790;
  wire w2791;
  wire w2792;
  wire w2793;
  wire w2794;
  wire w2795;
  wire w2796;
  wire w2797;
  wire w2798;
  wire w2799;
  wire w2800;
  wire w2801;
  wire w2802;
  wire w2803;
  wire w2804;
  wire w2805;
  wire w2806;
  wire w2807;
  wire w2808;
  wire w2809;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2854;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2860;
  wire w2861;
  wire w2862;
  wire w2863;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2896;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2913;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2934;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2950;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2979;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2990;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3014;
  wire w3015;
  wire w3016;
  wire w3017;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3040;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3084;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3094;
  wire w3095;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3121;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3130;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3225;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3254;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3262;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3272;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3327;
  wire w3328;
  wire w3329;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3334;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3362;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3366;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3414;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3433;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3443;
  wire w3444;
  wire w3445;
  wire w3446;
  wire w3447;
  wire w3448;
  wire w3449;
  wire w3450;
  wire w3451;
  wire w3452;
  wire w3453;
  wire w3454;
  wire w3455;
  wire w3456;
  wire w3457;
  wire w3458;
  wire w3459;
  wire w3460;
  wire w3461;
  wire w3462;
  wire w3463;
  wire w3464;
  wire w3465;
  wire w3466;
  wire w3467;
  wire w3468;
  wire w3469;
  wire w3470;
  wire w3471;
  wire w3472;
  wire w3473;
  wire w3474;
  wire w3475;
  wire w3476;
  wire w3477;
  wire w3478;
  wire w3479;
  wire w3480;
  wire w3481;
  wire w3482;
  wire w3483;
  wire w3484;
  wire w3486;
  wire w3487;
  wire w3488;
  wire w3489;
  wire w3490;
  wire w3491;
  wire w3492;
  wire w3493;
  wire w3494;
  wire w3495;
  wire w3496;
  wire w3497;
  wire w3498;
  wire w3499;
  wire w3500;
  wire w3501;
  wire w3502;
  wire w3503;
  wire w3504;
  wire w3505;
  wire w3506;
  wire w3507;
  wire w3508;
  wire w3509;
  wire w3510;
  wire w3511;
  wire w3512;
  wire w3513;
  wire w3514;
  wire w3515;
  wire w3516;
  wire w3517;
  wire w3518;
  wire w3519;
  wire w3520;
  wire w3521;
  wire w3522;
  wire w3523;
  wire w3524;
  wire w3525;
  wire w3526;
  wire w3527;
  wire w3528;
  wire w3529;
  wire w3530;
  wire w3531;
  wire w3532;
  wire w3533;
  wire w3534;
  wire w3535;
  wire w3536;
  wire w3537;
  wire w3538;
  wire w3539;
  wire w3540;
  wire w3541;
  wire w3542;
  wire w3543;
  wire w3544;
  wire w3545;
  wire w3546;
  wire w3547;
  wire w3548;
  wire w3549;
  wire w3550;
  wire w3551;
  wire w3552;
  wire w3553;
  wire w3554;
  wire w3555;
  wire w3556;
  wire w3557;
  wire w3558;
  wire w3559;
  wire w3560;
  wire w3561;
  wire w3562;
  wire w3563;
  wire w3564;
  wire w3565;
  wire w3566;
  wire w3567;
  wire w3568;
  wire w3569;
  wire w3570;
  wire w3571;
  wire w3572;
  wire w3573;
  wire w3574;
  wire w3575;
  wire w3576;
  wire w3577;
  wire w3578;
  wire w3579;
  wire w3580;
  wire w3581;
  wire w3582;
  wire w3583;
  wire w3584;
  wire w3586;
  wire w3587;
  wire w3588;
  wire w3589;
  wire w3590;
  wire w3591;
  wire w3592;
  wire w3593;
  wire w3594;
  wire w3595;
  wire w3596;
  wire w3597;
  wire w3598;
  wire w3599;
  wire w3600;
  wire w3601;
  wire w3602;
  wire w3603;
  wire w3604;
  wire w3605;
  wire w3606;
  wire w3607;
  wire w3608;
  wire w3609;
  wire w3610;
  wire w3611;
  wire w3612;
  wire w3613;
  wire w3614;
  wire w3615;
  wire w3616;
  wire w3617;
  wire w3618;
  wire w3619;
  wire w3620;
  wire w3621;
  wire w3622;
  wire w3623;
  wire w3624;
  wire w3625;
  wire w3626;
  wire w3627;
  wire w3628;
  wire w3629;
  wire w3630;
  wire w3631;
  wire w3632;
  wire w3633;
  wire w3634;
  wire w3635;
  wire w3636;
  wire w3637;
  wire w3638;
  wire w3639;
  wire w3640;
  wire w3641;
  wire w3642;
  wire w3643;
  wire w3644;
  wire w3645;
  wire w3646;
  wire w3647;
  wire w3648;
  wire w3649;
  wire w3650;
  wire w3651;
  wire w3652;
  wire w3653;
  wire w3654;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3662;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3734;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3742;
  wire w3743;
  wire w3744;
  wire w3745;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3762;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3768;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3814;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3836;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3849;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3862;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3882;
  wire w3883;
  wire w3884;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3894;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3930;
  wire w3931;
  wire w3932;
  wire w3933;
  wire w3934;
  wire w3935;
  wire w3936;
  wire w3937;
  wire w3938;
  wire w3939;
  wire w3940;
  wire w3941;
  wire w3942;
  wire w3943;
  wire w3944;
  wire w3945;
  wire w3946;
  wire w3947;
  wire w3948;
  wire w3949;
  wire w3950;
  wire w3951;
  wire w3952;
  wire w3953;
  wire w3954;
  wire w3955;
  wire w3956;
  wire w3957;
  wire w3958;
  wire w3959;
  wire w3960;
  wire w3961;
  wire w3962;
  wire w3963;
  wire w3964;
  wire w3965;
  wire w3966;
  wire w3967;
  wire w3968;
  wire w3969;
  wire w3970;
  wire w3971;
  wire w3972;
  wire w3973;
  wire w3974;
  wire w3975;
  wire w3976;
  wire w3977;
  wire w3978;
  wire w3979;
  wire w3980;
  wire w3981;
  wire w3982;
  wire w3983;
  wire w3984;
  wire w3986;
  wire w3987;
  wire w3988;
  wire w3989;
  wire w3990;
  wire w3991;
  wire w3992;
  wire w3993;
  wire w3994;
  wire w3995;
  wire w3996;
  wire w3997;
  wire w3998;
  wire w3999;
  wire w4000;
  wire w4001;
  wire w4002;
  wire w4003;
  wire w4004;
  wire w4005;
  wire w4006;
  wire w4007;
  wire w4008;
  wire w4009;
  wire w4010;
  wire w4011;
  wire w4012;
  wire w4013;
  wire w4014;
  wire w4015;
  wire w4016;
  wire w4017;
  wire w4018;
  wire w4019;
  wire w4020;
  wire w4021;
  wire w4022;
  wire w4023;
  wire w4024;
  wire w4025;
  wire w4026;
  wire w4027;
  wire w4028;
  wire w4029;
  wire w4030;
  wire w4031;
  wire w4032;
  wire w4033;
  wire w4034;
  wire w4035;
  wire w4036;
  wire w4037;
  wire w4038;
  wire w4039;
  wire w4040;
  wire w4041;
  wire w4042;
  wire w4043;
  wire w4044;
  wire w4045;
  wire w4046;
  wire w4047;
  wire w4048;
  wire w4049;
  wire w4050;
  wire w4051;
  wire w4052;
  wire w4053;
  wire w4054;
  wire w4055;
  wire w4056;
  wire w4057;
  wire w4058;
  wire w4059;
  wire w4060;
  wire w4061;
  wire w4062;
  wire w4063;
  wire w4064;
  wire w4065;
  wire w4066;
  wire w4067;
  wire w4068;
  wire w4069;
  wire w4070;
  wire w4071;
  wire w4072;
  wire w4073;
  wire w4074;
  wire w4075;
  wire w4076;
  wire w4077;
  wire w4078;
  wire w4079;
  wire w4080;
  wire w4081;
  wire w4082;
  wire w4083;
  wire w4084;
  wire w4086;
  wire w4087;
  wire w4088;
  wire w4089;
  wire w4090;
  wire w4091;
  wire w4092;
  wire w4093;
  wire w4094;
  wire w4095;
  wire w4096;
  wire w4097;
  wire w4098;
  wire w4099;
  wire w4100;
  wire w4101;
  wire w4102;
  wire w4103;
  wire w4104;
  wire w4105;
  wire w4106;
  wire w4107;
  wire w4108;
  wire w4109;
  wire w4110;
  wire w4111;
  wire w4112;
  wire w4113;
  wire w4114;
  wire w4115;
  wire w4116;
  wire w4117;
  wire w4118;
  wire w4119;
  wire w4120;
  wire w4121;
  wire w4122;
  wire w4123;
  wire w4124;
  wire w4125;
  wire w4126;
  wire w4127;
  wire w4128;
  wire w4129;
  wire w4130;
  wire w4131;
  wire w4132;
  wire w4133;
  wire w4134;
  wire w4135;
  wire w4136;
  wire w4137;
  wire w4138;
  wire w4139;
  wire w4140;
  wire w4141;
  wire w4142;
  wire w4143;
  wire w4144;
  wire w4145;
  wire w4146;
  wire w4147;
  wire w4148;
  wire w4149;
  wire w4150;
  wire w4151;
  wire w4152;
  wire w4153;
  wire w4154;
  wire w4155;
  wire w4156;
  wire w4157;
  wire w4158;
  wire w4159;
  wire w4160;
  wire w4161;
  wire w4162;
  wire w4163;
  wire w4164;
  wire w4165;
  wire w4166;
  wire w4167;
  wire w4168;
  wire w4169;
  wire w4170;
  wire w4171;
  wire w4172;
  wire w4173;
  wire w4174;
  wire w4175;
  wire w4176;
  wire w4177;
  wire w4178;
  wire w4179;
  wire w4180;
  wire w4181;
  wire w4182;
  wire w4183;
  wire w4184;
  wire w4186;
  wire w4187;
  wire w4188;
  wire w4189;
  wire w4190;
  wire w4191;
  wire w4192;
  wire w4193;
  wire w4194;
  wire w4195;
  wire w4196;
  wire w4197;
  wire w4198;
  wire w4199;
  wire w4200;
  wire w4201;
  wire w4202;
  wire w4203;
  wire w4204;
  wire w4205;
  wire w4206;
  wire w4207;
  wire w4208;
  wire w4209;
  wire w4210;
  wire w4211;
  wire w4212;
  wire w4213;
  wire w4214;
  wire w4215;
  wire w4216;
  wire w4217;
  wire w4218;
  wire w4219;
  wire w4220;
  wire w4221;
  wire w4222;
  wire w4223;
  wire w4224;
  wire w4225;
  wire w4226;
  wire w4227;
  wire w4228;
  wire w4229;
  wire w4230;
  wire w4231;
  wire w4232;
  wire w4233;
  wire w4234;
  wire w4235;
  wire w4236;
  wire w4237;
  wire w4238;
  wire w4239;
  wire w4240;
  wire w4241;
  wire w4242;
  wire w4243;
  wire w4244;
  wire w4245;
  wire w4246;
  wire w4247;
  wire w4248;
  wire w4249;
  wire w4250;
  wire w4251;
  wire w4252;
  wire w4253;
  wire w4254;
  wire w4255;
  wire w4256;
  wire w4257;
  wire w4258;
  wire w4259;
  wire w4260;
  wire w4261;
  wire w4262;
  wire w4263;
  wire w4264;
  wire w4265;
  wire w4266;
  wire w4267;
  wire w4268;
  wire w4269;
  wire w4270;
  wire w4271;
  wire w4272;
  wire w4273;
  wire w4274;
  wire w4275;
  wire w4276;
  wire w4277;
  wire w4278;
  wire w4279;
  wire w4280;
  wire w4281;
  wire w4282;
  wire w4283;
  wire w4284;
  wire w4286;
  wire w4287;
  wire w4288;
  wire w4289;
  wire w4290;
  wire w4291;
  wire w4292;
  wire w4293;
  wire w4294;
  wire w4295;
  wire w4296;
  wire w4297;
  wire w4298;
  wire w4299;
  wire w4300;
  wire w4301;
  wire w4302;
  wire w4303;
  wire w4304;
  wire w4305;
  wire w4306;
  wire w4307;
  wire w4308;
  wire w4309;
  wire w4310;
  wire w4311;
  wire w4312;
  wire w4313;
  wire w4314;
  wire w4315;
  wire w4316;
  wire w4317;
  wire w4318;
  wire w4319;
  wire w4320;
  wire w4321;
  wire w4322;
  wire w4323;
  wire w4324;
  wire w4325;
  wire w4326;
  wire w4327;
  wire w4328;
  wire w4329;
  wire w4330;
  wire w4331;
  wire w4332;
  wire w4333;
  wire w4334;
  wire w4335;
  wire w4336;
  wire w4337;
  wire w4338;
  wire w4339;
  wire w4340;
  wire w4341;
  wire w4342;
  wire w4343;
  wire w4344;
  wire w4345;
  wire w4346;
  wire w4347;
  wire w4348;
  wire w4349;
  wire w4350;
  wire w4351;
  wire w4352;
  wire w4353;
  wire w4354;
  wire w4355;
  wire w4356;
  wire w4357;
  wire w4358;
  wire w4359;
  wire w4360;
  wire w4361;
  wire w4362;
  wire w4363;
  wire w4364;
  wire w4365;
  wire w4366;
  wire w4367;
  wire w4368;
  wire w4369;
  wire w4370;
  wire w4371;
  wire w4372;
  wire w4373;
  wire w4374;
  wire w4375;
  wire w4376;
  wire w4377;
  wire w4378;
  wire w4379;
  wire w4380;
  wire w4381;
  wire w4382;
  wire w4383;
  wire w4384;
  wire w4386;
  wire w4387;
  wire w4388;
  wire w4389;
  wire w4390;
  wire w4391;
  wire w4392;
  wire w4393;
  wire w4394;
  wire w4395;
  wire w4396;
  wire w4397;
  wire w4398;
  wire w4399;
  wire w4400;
  wire w4401;
  wire w4402;
  wire w4403;
  wire w4404;
  wire w4405;
  wire w4406;
  wire w4407;
  wire w4408;
  wire w4409;
  wire w4410;
  wire w4411;
  wire w4412;
  wire w4413;
  wire w4414;
  wire w4415;
  wire w4416;
  wire w4417;
  wire w4418;
  wire w4419;
  wire w4420;
  wire w4421;
  wire w4422;
  wire w4423;
  wire w4424;
  wire w4425;
  wire w4426;
  wire w4427;
  wire w4428;
  wire w4429;
  wire w4430;
  wire w4431;
  wire w4432;
  wire w4433;
  wire w4434;
  wire w4435;
  wire w4436;
  wire w4437;
  wire w4438;
  wire w4439;
  wire w4440;
  wire w4441;
  wire w4442;
  wire w4443;
  wire w4444;
  wire w4445;
  wire w4446;
  wire w4447;
  wire w4448;
  wire w4449;
  wire w4450;
  wire w4451;
  wire w4452;
  wire w4453;
  wire w4454;
  wire w4455;
  wire w4456;
  wire w4457;
  wire w4458;
  wire w4459;
  wire w4460;
  wire w4461;
  wire w4462;
  wire w4463;
  wire w4464;
  wire w4465;
  wire w4466;
  wire w4467;
  wire w4468;
  wire w4469;
  wire w4470;
  wire w4471;
  wire w4472;
  wire w4473;
  wire w4474;
  wire w4475;
  wire w4476;
  wire w4477;
  wire w4478;
  wire w4479;
  wire w4480;
  wire w4481;
  wire w4482;
  wire w4483;
  wire w4484;
  wire w4486;
  wire w4487;
  wire w4488;
  wire w4489;
  wire w4490;
  wire w4491;
  wire w4492;
  wire w4493;
  wire w4494;
  wire w4495;
  wire w4496;
  wire w4497;
  wire w4498;
  wire w4499;
  wire w4500;
  wire w4501;
  wire w4502;
  wire w4503;
  wire w4504;
  wire w4505;
  wire w4506;
  wire w4507;
  wire w4508;
  wire w4509;
  wire w4510;
  wire w4511;
  wire w4512;
  wire w4513;
  wire w4514;
  wire w4515;
  wire w4516;
  wire w4517;
  wire w4518;
  wire w4519;
  wire w4520;
  wire w4521;
  wire w4522;
  wire w4523;
  wire w4524;
  wire w4525;
  wire w4526;
  wire w4527;
  wire w4528;
  wire w4529;
  wire w4530;
  wire w4531;
  wire w4532;
  wire w4533;
  wire w4534;
  wire w4535;
  wire w4536;
  wire w4537;
  wire w4538;
  wire w4539;
  wire w4540;
  wire w4541;
  wire w4542;
  wire w4543;
  wire w4544;
  wire w4545;
  wire w4546;
  wire w4547;
  wire w4548;
  wire w4549;
  wire w4550;
  wire w4551;
  wire w4552;
  wire w4553;
  wire w4554;
  wire w4555;
  wire w4556;
  wire w4557;
  wire w4558;
  wire w4559;
  wire w4560;
  wire w4561;
  wire w4562;
  wire w4563;
  wire w4564;
  wire w4565;
  wire w4566;
  wire w4567;
  wire w4568;
  wire w4569;
  wire w4570;
  wire w4571;
  wire w4572;
  wire w4573;
  wire w4574;
  wire w4575;
  wire w4576;
  wire w4577;
  wire w4578;
  wire w4579;
  wire w4580;
  wire w4581;
  wire w4582;
  wire w4583;
  wire w4584;
  wire w4586;
  wire w4587;
  wire w4588;
  wire w4589;
  wire w4590;
  wire w4591;
  wire w4592;
  wire w4593;
  wire w4594;
  wire w4595;
  wire w4596;
  wire w4597;
  wire w4598;
  wire w4599;
  wire w4600;
  wire w4601;
  wire w4602;
  wire w4603;
  wire w4604;
  wire w4605;
  wire w4606;
  wire w4607;
  wire w4608;
  wire w4609;
  wire w4610;
  wire w4611;
  wire w4612;
  wire w4613;
  wire w4614;
  wire w4615;
  wire w4616;
  wire w4617;
  wire w4618;
  wire w4619;
  wire w4620;
  wire w4621;
  wire w4622;
  wire w4623;
  wire w4624;
  wire w4625;
  wire w4626;
  wire w4627;
  wire w4628;
  wire w4629;
  wire w4630;
  wire w4631;
  wire w4632;
  wire w4633;
  wire w4634;
  wire w4635;
  wire w4636;
  wire w4637;
  wire w4638;
  wire w4639;
  wire w4640;
  wire w4641;
  wire w4642;
  wire w4643;
  wire w4644;
  wire w4645;
  wire w4646;
  wire w4647;
  wire w4648;
  wire w4649;
  wire w4650;
  wire w4651;
  wire w4652;
  wire w4653;
  wire w4654;
  wire w4655;
  wire w4656;
  wire w4657;
  wire w4658;
  wire w4659;
  wire w4660;
  wire w4661;
  wire w4662;
  wire w4663;
  wire w4664;
  wire w4665;
  wire w4666;
  wire w4667;
  wire w4668;
  wire w4669;
  wire w4670;
  wire w4671;
  wire w4672;
  wire w4673;
  wire w4674;
  wire w4675;
  wire w4676;
  wire w4677;
  wire w4678;
  wire w4679;
  wire w4680;
  wire w4681;
  wire w4682;
  wire w4683;
  wire w4684;
  wire w4686;
  wire w4687;
  wire w4688;
  wire w4689;
  wire w4690;
  wire w4691;
  wire w4692;
  wire w4693;
  wire w4694;
  wire w4695;
  wire w4696;
  wire w4697;
  wire w4698;
  wire w4699;
  wire w4700;
  wire w4701;
  wire w4702;
  wire w4703;
  wire w4704;
  wire w4705;
  wire w4706;
  wire w4707;
  wire w4708;
  wire w4709;
  wire w4710;
  wire w4711;
  wire w4712;
  wire w4713;
  wire w4714;
  wire w4715;
  wire w4716;
  wire w4717;
  wire w4718;
  wire w4719;
  wire w4720;
  wire w4721;
  wire w4722;
  wire w4723;
  wire w4724;
  wire w4725;
  wire w4726;
  wire w4727;
  wire w4728;
  wire w4729;
  wire w4730;
  wire w4731;
  wire w4732;
  wire w4733;
  wire w4734;
  wire w4735;
  wire w4736;
  wire w4737;
  wire w4738;
  wire w4739;
  wire w4740;
  wire w4741;
  wire w4742;
  wire w4743;
  wire w4744;
  wire w4745;
  wire w4746;
  wire w4747;
  wire w4748;
  wire w4749;
  wire w4750;
  wire w4751;
  wire w4752;
  wire w4753;
  wire w4754;
  wire w4755;
  wire w4756;
  wire w4757;
  wire w4758;
  wire w4759;
  wire w4760;
  wire w4761;
  wire w4762;
  wire w4763;
  wire w4764;
  wire w4765;
  wire w4766;
  wire w4767;
  wire w4768;
  wire w4769;
  wire w4770;
  wire w4771;
  wire w4772;
  wire w4773;
  wire w4774;
  wire w4775;
  wire w4776;
  wire w4777;
  wire w4778;
  wire w4779;
  wire w4780;
  wire w4781;
  wire w4782;
  wire w4783;
  wire w4784;
  wire w4786;
  wire w4787;
  wire w4788;
  wire w4789;
  wire w4790;
  wire w4791;
  wire w4792;
  wire w4793;
  wire w4794;
  wire w4795;
  wire w4796;
  wire w4797;
  wire w4798;
  wire w4799;
  wire w4800;
  wire w4801;
  wire w4802;
  wire w4803;
  wire w4804;
  wire w4805;
  wire w4806;
  wire w4807;
  wire w4808;
  wire w4809;
  wire w4810;
  wire w4811;
  wire w4812;
  wire w4813;
  wire w4814;
  wire w4815;
  wire w4816;
  wire w4817;
  wire w4818;
  wire w4819;
  wire w4820;
  wire w4821;
  wire w4822;
  wire w4823;
  wire w4824;
  wire w4825;
  wire w4826;
  wire w4827;
  wire w4828;
  wire w4829;
  wire w4830;
  wire w4831;
  wire w4832;
  wire w4833;
  wire w4834;
  wire w4835;
  wire w4836;
  wire w4837;
  wire w4838;
  wire w4839;
  wire w4840;
  wire w4841;
  wire w4842;
  wire w4843;
  wire w4844;
  wire w4845;
  wire w4846;
  wire w4847;
  wire w4848;
  wire w4849;
  wire w4850;
  wire w4851;
  wire w4852;
  wire w4853;
  wire w4854;
  wire w4855;
  wire w4856;
  wire w4857;
  wire w4858;
  wire w4859;
  wire w4860;
  wire w4861;
  wire w4862;
  wire w4863;
  wire w4864;
  wire w4865;
  wire w4866;
  wire w4867;
  wire w4868;
  wire w4869;
  wire w4870;
  wire w4871;
  wire w4872;
  wire w4873;
  wire w4874;
  wire w4875;
  wire w4876;
  wire w4877;
  wire w4878;
  wire w4879;
  wire w4880;
  wire w4881;
  wire w4882;
  wire w4883;
  wire w4884;
  wire w4886;
  wire w4887;
  wire w4888;
  wire w4889;
  wire w4890;
  wire w4891;
  wire w4892;
  wire w4893;
  wire w4894;
  wire w4895;
  wire w4896;
  wire w4897;
  wire w4898;
  wire w4899;
  wire w4900;
  wire w4901;
  wire w4902;
  wire w4903;
  wire w4904;
  wire w4905;
  wire w4906;
  wire w4907;
  wire w4908;
  wire w4909;
  wire w4910;
  wire w4911;
  wire w4912;
  wire w4913;
  wire w4914;
  wire w4915;
  wire w4916;
  wire w4917;
  wire w4918;
  wire w4919;
  wire w4920;
  wire w4921;
  wire w4922;
  wire w4923;
  wire w4924;
  wire w4925;
  wire w4926;
  wire w4927;
  wire w4928;
  wire w4929;
  wire w4930;
  wire w4931;
  wire w4932;
  wire w4933;
  wire w4934;
  wire w4935;
  wire w4936;
  wire w4937;
  wire w4938;
  wire w4939;
  wire w4940;
  wire w4941;
  wire w4942;
  wire w4943;
  wire w4944;
  wire w4945;
  wire w4946;
  wire w4947;
  wire w4948;
  wire w4949;
  wire w4950;
  wire w4951;
  wire w4952;
  wire w4953;
  wire w4954;
  wire w4955;
  wire w4956;
  wire w4957;
  wire w4958;
  wire w4959;
  wire w4960;
  wire w4961;
  wire w4962;
  wire w4963;
  wire w4964;
  wire w4965;
  wire w4966;
  wire w4967;
  wire w4968;
  wire w4969;
  wire w4970;
  wire w4971;
  wire w4972;
  wire w4973;
  wire w4974;
  wire w4975;
  wire w4976;
  wire w4977;
  wire w4978;
  wire w4979;
  wire w4980;
  wire w4981;
  wire w4982;
  wire w4983;
  wire w4984;
  wire w4986;
  wire w4987;
  wire w4988;
  wire w4989;
  wire w4990;
  wire w4991;
  wire w4992;
  wire w4993;
  wire w4994;
  wire w4995;
  wire w4996;
  wire w4997;
  wire w4998;
  wire w4999;
  wire w5000;
  wire w5001;
  wire w5002;
  wire w5003;
  wire w5004;
  wire w5005;
  wire w5006;
  wire w5007;
  wire w5008;
  wire w5009;
  wire w5010;
  wire w5011;
  wire w5012;
  wire w5013;
  wire w5014;
  wire w5015;
  wire w5016;
  wire w5017;
  wire w5018;
  wire w5019;
  wire w5020;
  wire w5021;
  wire w5022;
  wire w5023;
  wire w5024;
  wire w5025;
  wire w5026;
  wire w5027;
  wire w5028;
  wire w5029;
  wire w5030;
  wire w5031;
  wire w5032;
  wire w5033;
  wire w5034;
  wire w5035;
  wire w5036;
  wire w5037;
  wire w5038;
  wire w5039;
  wire w5040;
  wire w5041;
  wire w5042;
  wire w5043;
  wire w5044;
  wire w5045;
  wire w5046;
  wire w5047;
  wire w5048;
  wire w5049;
  wire w5050;
  wire w5051;
  wire w5052;
  wire w5053;
  wire w5054;
  wire w5055;
  wire w5056;
  wire w5057;
  wire w5058;
  wire w5059;
  wire w5060;
  wire w5061;
  wire w5062;
  wire w5063;
  wire w5064;
  wire w5065;
  wire w5066;
  wire w5067;
  wire w5068;
  wire w5069;
  wire w5070;
  wire w5071;
  wire w5072;
  wire w5073;
  wire w5074;
  wire w5075;
  wire w5076;
  wire w5077;
  wire w5078;
  wire w5079;
  wire w5080;
  wire w5081;
  wire w5082;
  wire w5083;
  wire w5084;
  wire w5086;
  wire w5088;
  wire w5090;
  wire w5092;
  wire w5094;
  wire w5096;
  wire w5098;
  wire w5100;
  wire w5102;
  wire w5104;
  wire w5106;
  wire w5108;
  wire w5110;
  wire w5112;
  wire w5114;
  wire w5116;
  wire w5118;
  wire w5120;
  wire w5122;
  wire w5124;
  wire w5126;
  wire w5128;
  wire w5130;
  wire w5132;
  wire w5134;
  wire w5136;
  wire w5138;
  wire w5140;
  wire w5142;
  wire w5144;
  wire w5146;
  wire w5148;
  wire w5150;
  wire w5152;
  wire w5154;
  wire w5156;
  wire w5158;
  wire w5160;
  wire w5162;
  wire w5164;
  wire w5166;
  wire w5168;
  wire w5170;
  wire w5172;
  wire w5174;
  wire w5176;
  wire w5178;
  wire w5180;
  wire w5182;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w1786);
  FullAdder U1 (w1786, IN2[0], IN2[1], w1787, w1788);
  FullAdder U2 (w1788, IN3[0], IN3[1], w1789, w1790);
  FullAdder U3 (w1790, IN4[0], IN4[1], w1791, w1792);
  FullAdder U4 (w1792, IN5[0], IN5[1], w1793, w1794);
  FullAdder U5 (w1794, IN6[0], IN6[1], w1795, w1796);
  FullAdder U6 (w1796, IN7[0], IN7[1], w1797, w1798);
  FullAdder U7 (w1798, IN8[0], IN8[1], w1799, w1800);
  FullAdder U8 (w1800, IN9[0], IN9[1], w1801, w1802);
  FullAdder U9 (w1802, IN10[0], IN10[1], w1803, w1804);
  FullAdder U10 (w1804, IN11[0], IN11[1], w1805, w1806);
  FullAdder U11 (w1806, IN12[0], IN12[1], w1807, w1808);
  FullAdder U12 (w1808, IN13[0], IN13[1], w1809, w1810);
  FullAdder U13 (w1810, IN14[0], IN14[1], w1811, w1812);
  FullAdder U14 (w1812, IN15[0], IN15[1], w1813, w1814);
  FullAdder U15 (w1814, IN16[0], IN16[1], w1815, w1816);
  FullAdder U16 (w1816, IN17[0], IN17[1], w1817, w1818);
  FullAdder U17 (w1818, IN18[0], IN18[1], w1819, w1820);
  FullAdder U18 (w1820, IN19[0], IN19[1], w1821, w1822);
  FullAdder U19 (w1822, IN20[0], IN20[1], w1823, w1824);
  FullAdder U20 (w1824, IN21[0], IN21[1], w1825, w1826);
  FullAdder U21 (w1826, IN22[0], IN22[1], w1827, w1828);
  FullAdder U22 (w1828, IN23[0], IN23[1], w1829, w1830);
  FullAdder U23 (w1830, IN24[0], IN24[1], w1831, w1832);
  FullAdder U24 (w1832, IN25[0], IN25[1], w1833, w1834);
  FullAdder U25 (w1834, IN26[0], IN26[1], w1835, w1836);
  FullAdder U26 (w1836, IN27[0], IN27[1], w1837, w1838);
  FullAdder U27 (w1838, IN28[0], IN28[1], w1839, w1840);
  FullAdder U28 (w1840, IN29[0], IN29[1], w1841, w1842);
  FullAdder U29 (w1842, IN30[0], IN30[1], w1843, w1844);
  FullAdder U30 (w1844, IN31[0], IN31[1], w1845, w1846);
  FullAdder U31 (w1846, IN32[0], IN32[1], w1847, w1848);
  FullAdder U32 (w1848, IN33[0], IN33[1], w1849, w1850);
  FullAdder U33 (w1850, IN34[0], IN34[1], w1851, w1852);
  FullAdder U34 (w1852, IN35[0], IN35[1], w1853, w1854);
  FullAdder U35 (w1854, IN36[0], IN36[1], w1855, w1856);
  FullAdder U36 (w1856, IN37[0], IN37[1], w1857, w1858);
  FullAdder U37 (w1858, IN38[0], IN38[1], w1859, w1860);
  FullAdder U38 (w1860, IN39[0], IN39[1], w1861, w1862);
  FullAdder U39 (w1862, IN40[0], IN40[1], w1863, w1864);
  FullAdder U40 (w1864, IN41[0], IN41[1], w1865, w1866);
  FullAdder U41 (w1866, IN42[0], IN42[1], w1867, w1868);
  FullAdder U42 (w1868, IN43[0], IN43[1], w1869, w1870);
  FullAdder U43 (w1870, IN44[0], IN44[1], w1871, w1872);
  FullAdder U44 (w1872, IN45[0], IN45[1], w1873, w1874);
  FullAdder U45 (w1874, IN46[0], IN46[1], w1875, w1876);
  FullAdder U46 (w1876, IN47[0], IN47[1], w1877, w1878);
  FullAdder U47 (w1878, IN48[0], IN48[1], w1879, w1880);
  FullAdder U48 (w1880, IN49[0], IN49[1], w1881, w1882);
  FullAdder U49 (w1882, IN50[0], IN50[1], w1883, w1884);
  HalfAdder U50 (w1787, IN2[2], Out1[2], w1886);
  FullAdder U51 (w1886, w1789, IN3[2], w1887, w1888);
  FullAdder U52 (w1888, w1791, IN4[2], w1889, w1890);
  FullAdder U53 (w1890, w1793, IN5[2], w1891, w1892);
  FullAdder U54 (w1892, w1795, IN6[2], w1893, w1894);
  FullAdder U55 (w1894, w1797, IN7[2], w1895, w1896);
  FullAdder U56 (w1896, w1799, IN8[2], w1897, w1898);
  FullAdder U57 (w1898, w1801, IN9[2], w1899, w1900);
  FullAdder U58 (w1900, w1803, IN10[2], w1901, w1902);
  FullAdder U59 (w1902, w1805, IN11[2], w1903, w1904);
  FullAdder U60 (w1904, w1807, IN12[2], w1905, w1906);
  FullAdder U61 (w1906, w1809, IN13[2], w1907, w1908);
  FullAdder U62 (w1908, w1811, IN14[2], w1909, w1910);
  FullAdder U63 (w1910, w1813, IN15[2], w1911, w1912);
  FullAdder U64 (w1912, w1815, IN16[2], w1913, w1914);
  FullAdder U65 (w1914, w1817, IN17[2], w1915, w1916);
  FullAdder U66 (w1916, w1819, IN18[2], w1917, w1918);
  FullAdder U67 (w1918, w1821, IN19[2], w1919, w1920);
  FullAdder U68 (w1920, w1823, IN20[2], w1921, w1922);
  FullAdder U69 (w1922, w1825, IN21[2], w1923, w1924);
  FullAdder U70 (w1924, w1827, IN22[2], w1925, w1926);
  FullAdder U71 (w1926, w1829, IN23[2], w1927, w1928);
  FullAdder U72 (w1928, w1831, IN24[2], w1929, w1930);
  FullAdder U73 (w1930, w1833, IN25[2], w1931, w1932);
  FullAdder U74 (w1932, w1835, IN26[2], w1933, w1934);
  FullAdder U75 (w1934, w1837, IN27[2], w1935, w1936);
  FullAdder U76 (w1936, w1839, IN28[2], w1937, w1938);
  FullAdder U77 (w1938, w1841, IN29[2], w1939, w1940);
  FullAdder U78 (w1940, w1843, IN30[2], w1941, w1942);
  FullAdder U79 (w1942, w1845, IN31[2], w1943, w1944);
  FullAdder U80 (w1944, w1847, IN32[2], w1945, w1946);
  FullAdder U81 (w1946, w1849, IN33[2], w1947, w1948);
  FullAdder U82 (w1948, w1851, IN34[2], w1949, w1950);
  FullAdder U83 (w1950, w1853, IN35[2], w1951, w1952);
  FullAdder U84 (w1952, w1855, IN36[2], w1953, w1954);
  FullAdder U85 (w1954, w1857, IN37[2], w1955, w1956);
  FullAdder U86 (w1956, w1859, IN38[2], w1957, w1958);
  FullAdder U87 (w1958, w1861, IN39[2], w1959, w1960);
  FullAdder U88 (w1960, w1863, IN40[2], w1961, w1962);
  FullAdder U89 (w1962, w1865, IN41[2], w1963, w1964);
  FullAdder U90 (w1964, w1867, IN42[2], w1965, w1966);
  FullAdder U91 (w1966, w1869, IN43[2], w1967, w1968);
  FullAdder U92 (w1968, w1871, IN44[2], w1969, w1970);
  FullAdder U93 (w1970, w1873, IN45[2], w1971, w1972);
  FullAdder U94 (w1972, w1875, IN46[2], w1973, w1974);
  FullAdder U95 (w1974, w1877, IN47[2], w1975, w1976);
  FullAdder U96 (w1976, w1879, IN48[2], w1977, w1978);
  FullAdder U97 (w1978, w1881, IN49[2], w1979, w1980);
  FullAdder U98 (w1980, w1883, IN50[2], w1981, w1982);
  FullAdder U99 (w1982, w1884, IN51[0], w1983, w1984);
  HalfAdder U100 (w1887, IN3[3], Out1[3], w1986);
  FullAdder U101 (w1986, w1889, IN4[3], w1987, w1988);
  FullAdder U102 (w1988, w1891, IN5[3], w1989, w1990);
  FullAdder U103 (w1990, w1893, IN6[3], w1991, w1992);
  FullAdder U104 (w1992, w1895, IN7[3], w1993, w1994);
  FullAdder U105 (w1994, w1897, IN8[3], w1995, w1996);
  FullAdder U106 (w1996, w1899, IN9[3], w1997, w1998);
  FullAdder U107 (w1998, w1901, IN10[3], w1999, w2000);
  FullAdder U108 (w2000, w1903, IN11[3], w2001, w2002);
  FullAdder U109 (w2002, w1905, IN12[3], w2003, w2004);
  FullAdder U110 (w2004, w1907, IN13[3], w2005, w2006);
  FullAdder U111 (w2006, w1909, IN14[3], w2007, w2008);
  FullAdder U112 (w2008, w1911, IN15[3], w2009, w2010);
  FullAdder U113 (w2010, w1913, IN16[3], w2011, w2012);
  FullAdder U114 (w2012, w1915, IN17[3], w2013, w2014);
  FullAdder U115 (w2014, w1917, IN18[3], w2015, w2016);
  FullAdder U116 (w2016, w1919, IN19[3], w2017, w2018);
  FullAdder U117 (w2018, w1921, IN20[3], w2019, w2020);
  FullAdder U118 (w2020, w1923, IN21[3], w2021, w2022);
  FullAdder U119 (w2022, w1925, IN22[3], w2023, w2024);
  FullAdder U120 (w2024, w1927, IN23[3], w2025, w2026);
  FullAdder U121 (w2026, w1929, IN24[3], w2027, w2028);
  FullAdder U122 (w2028, w1931, IN25[3], w2029, w2030);
  FullAdder U123 (w2030, w1933, IN26[3], w2031, w2032);
  FullAdder U124 (w2032, w1935, IN27[3], w2033, w2034);
  FullAdder U125 (w2034, w1937, IN28[3], w2035, w2036);
  FullAdder U126 (w2036, w1939, IN29[3], w2037, w2038);
  FullAdder U127 (w2038, w1941, IN30[3], w2039, w2040);
  FullAdder U128 (w2040, w1943, IN31[3], w2041, w2042);
  FullAdder U129 (w2042, w1945, IN32[3], w2043, w2044);
  FullAdder U130 (w2044, w1947, IN33[3], w2045, w2046);
  FullAdder U131 (w2046, w1949, IN34[3], w2047, w2048);
  FullAdder U132 (w2048, w1951, IN35[3], w2049, w2050);
  FullAdder U133 (w2050, w1953, IN36[3], w2051, w2052);
  FullAdder U134 (w2052, w1955, IN37[3], w2053, w2054);
  FullAdder U135 (w2054, w1957, IN38[3], w2055, w2056);
  FullAdder U136 (w2056, w1959, IN39[3], w2057, w2058);
  FullAdder U137 (w2058, w1961, IN40[3], w2059, w2060);
  FullAdder U138 (w2060, w1963, IN41[3], w2061, w2062);
  FullAdder U139 (w2062, w1965, IN42[3], w2063, w2064);
  FullAdder U140 (w2064, w1967, IN43[3], w2065, w2066);
  FullAdder U141 (w2066, w1969, IN44[3], w2067, w2068);
  FullAdder U142 (w2068, w1971, IN45[3], w2069, w2070);
  FullAdder U143 (w2070, w1973, IN46[3], w2071, w2072);
  FullAdder U144 (w2072, w1975, IN47[3], w2073, w2074);
  FullAdder U145 (w2074, w1977, IN48[3], w2075, w2076);
  FullAdder U146 (w2076, w1979, IN49[3], w2077, w2078);
  FullAdder U147 (w2078, w1981, IN50[3], w2079, w2080);
  FullAdder U148 (w2080, w1983, IN51[1], w2081, w2082);
  FullAdder U149 (w2082, w1984, IN52[0], w2083, w2084);
  HalfAdder U150 (w1987, IN4[4], Out1[4], w2086);
  FullAdder U151 (w2086, w1989, IN5[4], w2087, w2088);
  FullAdder U152 (w2088, w1991, IN6[4], w2089, w2090);
  FullAdder U153 (w2090, w1993, IN7[4], w2091, w2092);
  FullAdder U154 (w2092, w1995, IN8[4], w2093, w2094);
  FullAdder U155 (w2094, w1997, IN9[4], w2095, w2096);
  FullAdder U156 (w2096, w1999, IN10[4], w2097, w2098);
  FullAdder U157 (w2098, w2001, IN11[4], w2099, w2100);
  FullAdder U158 (w2100, w2003, IN12[4], w2101, w2102);
  FullAdder U159 (w2102, w2005, IN13[4], w2103, w2104);
  FullAdder U160 (w2104, w2007, IN14[4], w2105, w2106);
  FullAdder U161 (w2106, w2009, IN15[4], w2107, w2108);
  FullAdder U162 (w2108, w2011, IN16[4], w2109, w2110);
  FullAdder U163 (w2110, w2013, IN17[4], w2111, w2112);
  FullAdder U164 (w2112, w2015, IN18[4], w2113, w2114);
  FullAdder U165 (w2114, w2017, IN19[4], w2115, w2116);
  FullAdder U166 (w2116, w2019, IN20[4], w2117, w2118);
  FullAdder U167 (w2118, w2021, IN21[4], w2119, w2120);
  FullAdder U168 (w2120, w2023, IN22[4], w2121, w2122);
  FullAdder U169 (w2122, w2025, IN23[4], w2123, w2124);
  FullAdder U170 (w2124, w2027, IN24[4], w2125, w2126);
  FullAdder U171 (w2126, w2029, IN25[4], w2127, w2128);
  FullAdder U172 (w2128, w2031, IN26[4], w2129, w2130);
  FullAdder U173 (w2130, w2033, IN27[4], w2131, w2132);
  FullAdder U174 (w2132, w2035, IN28[4], w2133, w2134);
  FullAdder U175 (w2134, w2037, IN29[4], w2135, w2136);
  FullAdder U176 (w2136, w2039, IN30[4], w2137, w2138);
  FullAdder U177 (w2138, w2041, IN31[4], w2139, w2140);
  FullAdder U178 (w2140, w2043, IN32[4], w2141, w2142);
  FullAdder U179 (w2142, w2045, IN33[4], w2143, w2144);
  FullAdder U180 (w2144, w2047, IN34[4], w2145, w2146);
  FullAdder U181 (w2146, w2049, IN35[4], w2147, w2148);
  FullAdder U182 (w2148, w2051, IN36[4], w2149, w2150);
  FullAdder U183 (w2150, w2053, IN37[4], w2151, w2152);
  FullAdder U184 (w2152, w2055, IN38[4], w2153, w2154);
  FullAdder U185 (w2154, w2057, IN39[4], w2155, w2156);
  FullAdder U186 (w2156, w2059, IN40[4], w2157, w2158);
  FullAdder U187 (w2158, w2061, IN41[4], w2159, w2160);
  FullAdder U188 (w2160, w2063, IN42[4], w2161, w2162);
  FullAdder U189 (w2162, w2065, IN43[4], w2163, w2164);
  FullAdder U190 (w2164, w2067, IN44[4], w2165, w2166);
  FullAdder U191 (w2166, w2069, IN45[4], w2167, w2168);
  FullAdder U192 (w2168, w2071, IN46[4], w2169, w2170);
  FullAdder U193 (w2170, w2073, IN47[4], w2171, w2172);
  FullAdder U194 (w2172, w2075, IN48[4], w2173, w2174);
  FullAdder U195 (w2174, w2077, IN49[4], w2175, w2176);
  FullAdder U196 (w2176, w2079, IN50[4], w2177, w2178);
  FullAdder U197 (w2178, w2081, IN51[2], w2179, w2180);
  FullAdder U198 (w2180, w2083, IN52[1], w2181, w2182);
  FullAdder U199 (w2182, w2084, IN53[0], w2183, w2184);
  HalfAdder U200 (w2087, IN5[5], Out1[5], w2186);
  FullAdder U201 (w2186, w2089, IN6[5], w2187, w2188);
  FullAdder U202 (w2188, w2091, IN7[5], w2189, w2190);
  FullAdder U203 (w2190, w2093, IN8[5], w2191, w2192);
  FullAdder U204 (w2192, w2095, IN9[5], w2193, w2194);
  FullAdder U205 (w2194, w2097, IN10[5], w2195, w2196);
  FullAdder U206 (w2196, w2099, IN11[5], w2197, w2198);
  FullAdder U207 (w2198, w2101, IN12[5], w2199, w2200);
  FullAdder U208 (w2200, w2103, IN13[5], w2201, w2202);
  FullAdder U209 (w2202, w2105, IN14[5], w2203, w2204);
  FullAdder U210 (w2204, w2107, IN15[5], w2205, w2206);
  FullAdder U211 (w2206, w2109, IN16[5], w2207, w2208);
  FullAdder U212 (w2208, w2111, IN17[5], w2209, w2210);
  FullAdder U213 (w2210, w2113, IN18[5], w2211, w2212);
  FullAdder U214 (w2212, w2115, IN19[5], w2213, w2214);
  FullAdder U215 (w2214, w2117, IN20[5], w2215, w2216);
  FullAdder U216 (w2216, w2119, IN21[5], w2217, w2218);
  FullAdder U217 (w2218, w2121, IN22[5], w2219, w2220);
  FullAdder U218 (w2220, w2123, IN23[5], w2221, w2222);
  FullAdder U219 (w2222, w2125, IN24[5], w2223, w2224);
  FullAdder U220 (w2224, w2127, IN25[5], w2225, w2226);
  FullAdder U221 (w2226, w2129, IN26[5], w2227, w2228);
  FullAdder U222 (w2228, w2131, IN27[5], w2229, w2230);
  FullAdder U223 (w2230, w2133, IN28[5], w2231, w2232);
  FullAdder U224 (w2232, w2135, IN29[5], w2233, w2234);
  FullAdder U225 (w2234, w2137, IN30[5], w2235, w2236);
  FullAdder U226 (w2236, w2139, IN31[5], w2237, w2238);
  FullAdder U227 (w2238, w2141, IN32[5], w2239, w2240);
  FullAdder U228 (w2240, w2143, IN33[5], w2241, w2242);
  FullAdder U229 (w2242, w2145, IN34[5], w2243, w2244);
  FullAdder U230 (w2244, w2147, IN35[5], w2245, w2246);
  FullAdder U231 (w2246, w2149, IN36[5], w2247, w2248);
  FullAdder U232 (w2248, w2151, IN37[5], w2249, w2250);
  FullAdder U233 (w2250, w2153, IN38[5], w2251, w2252);
  FullAdder U234 (w2252, w2155, IN39[5], w2253, w2254);
  FullAdder U235 (w2254, w2157, IN40[5], w2255, w2256);
  FullAdder U236 (w2256, w2159, IN41[5], w2257, w2258);
  FullAdder U237 (w2258, w2161, IN42[5], w2259, w2260);
  FullAdder U238 (w2260, w2163, IN43[5], w2261, w2262);
  FullAdder U239 (w2262, w2165, IN44[5], w2263, w2264);
  FullAdder U240 (w2264, w2167, IN45[5], w2265, w2266);
  FullAdder U241 (w2266, w2169, IN46[5], w2267, w2268);
  FullAdder U242 (w2268, w2171, IN47[5], w2269, w2270);
  FullAdder U243 (w2270, w2173, IN48[5], w2271, w2272);
  FullAdder U244 (w2272, w2175, IN49[5], w2273, w2274);
  FullAdder U245 (w2274, w2177, IN50[5], w2275, w2276);
  FullAdder U246 (w2276, w2179, IN51[3], w2277, w2278);
  FullAdder U247 (w2278, w2181, IN52[2], w2279, w2280);
  FullAdder U248 (w2280, w2183, IN53[1], w2281, w2282);
  FullAdder U249 (w2282, w2184, IN54[0], w2283, w2284);
  HalfAdder U250 (w2187, IN6[6], Out1[6], w2286);
  FullAdder U251 (w2286, w2189, IN7[6], w2287, w2288);
  FullAdder U252 (w2288, w2191, IN8[6], w2289, w2290);
  FullAdder U253 (w2290, w2193, IN9[6], w2291, w2292);
  FullAdder U254 (w2292, w2195, IN10[6], w2293, w2294);
  FullAdder U255 (w2294, w2197, IN11[6], w2295, w2296);
  FullAdder U256 (w2296, w2199, IN12[6], w2297, w2298);
  FullAdder U257 (w2298, w2201, IN13[6], w2299, w2300);
  FullAdder U258 (w2300, w2203, IN14[6], w2301, w2302);
  FullAdder U259 (w2302, w2205, IN15[6], w2303, w2304);
  FullAdder U260 (w2304, w2207, IN16[6], w2305, w2306);
  FullAdder U261 (w2306, w2209, IN17[6], w2307, w2308);
  FullAdder U262 (w2308, w2211, IN18[6], w2309, w2310);
  FullAdder U263 (w2310, w2213, IN19[6], w2311, w2312);
  FullAdder U264 (w2312, w2215, IN20[6], w2313, w2314);
  FullAdder U265 (w2314, w2217, IN21[6], w2315, w2316);
  FullAdder U266 (w2316, w2219, IN22[6], w2317, w2318);
  FullAdder U267 (w2318, w2221, IN23[6], w2319, w2320);
  FullAdder U268 (w2320, w2223, IN24[6], w2321, w2322);
  FullAdder U269 (w2322, w2225, IN25[6], w2323, w2324);
  FullAdder U270 (w2324, w2227, IN26[6], w2325, w2326);
  FullAdder U271 (w2326, w2229, IN27[6], w2327, w2328);
  FullAdder U272 (w2328, w2231, IN28[6], w2329, w2330);
  FullAdder U273 (w2330, w2233, IN29[6], w2331, w2332);
  FullAdder U274 (w2332, w2235, IN30[6], w2333, w2334);
  FullAdder U275 (w2334, w2237, IN31[6], w2335, w2336);
  FullAdder U276 (w2336, w2239, IN32[6], w2337, w2338);
  FullAdder U277 (w2338, w2241, IN33[6], w2339, w2340);
  FullAdder U278 (w2340, w2243, IN34[6], w2341, w2342);
  FullAdder U279 (w2342, w2245, IN35[6], w2343, w2344);
  FullAdder U280 (w2344, w2247, IN36[6], w2345, w2346);
  FullAdder U281 (w2346, w2249, IN37[6], w2347, w2348);
  FullAdder U282 (w2348, w2251, IN38[6], w2349, w2350);
  FullAdder U283 (w2350, w2253, IN39[6], w2351, w2352);
  FullAdder U284 (w2352, w2255, IN40[6], w2353, w2354);
  FullAdder U285 (w2354, w2257, IN41[6], w2355, w2356);
  FullAdder U286 (w2356, w2259, IN42[6], w2357, w2358);
  FullAdder U287 (w2358, w2261, IN43[6], w2359, w2360);
  FullAdder U288 (w2360, w2263, IN44[6], w2361, w2362);
  FullAdder U289 (w2362, w2265, IN45[6], w2363, w2364);
  FullAdder U290 (w2364, w2267, IN46[6], w2365, w2366);
  FullAdder U291 (w2366, w2269, IN47[6], w2367, w2368);
  FullAdder U292 (w2368, w2271, IN48[6], w2369, w2370);
  FullAdder U293 (w2370, w2273, IN49[6], w2371, w2372);
  FullAdder U294 (w2372, w2275, IN50[6], w2373, w2374);
  FullAdder U295 (w2374, w2277, IN51[4], w2375, w2376);
  FullAdder U296 (w2376, w2279, IN52[3], w2377, w2378);
  FullAdder U297 (w2378, w2281, IN53[2], w2379, w2380);
  FullAdder U298 (w2380, w2283, IN54[1], w2381, w2382);
  FullAdder U299 (w2382, w2284, IN55[0], w2383, w2384);
  HalfAdder U300 (w2287, IN7[7], Out1[7], w2386);
  FullAdder U301 (w2386, w2289, IN8[7], w2387, w2388);
  FullAdder U302 (w2388, w2291, IN9[7], w2389, w2390);
  FullAdder U303 (w2390, w2293, IN10[7], w2391, w2392);
  FullAdder U304 (w2392, w2295, IN11[7], w2393, w2394);
  FullAdder U305 (w2394, w2297, IN12[7], w2395, w2396);
  FullAdder U306 (w2396, w2299, IN13[7], w2397, w2398);
  FullAdder U307 (w2398, w2301, IN14[7], w2399, w2400);
  FullAdder U308 (w2400, w2303, IN15[7], w2401, w2402);
  FullAdder U309 (w2402, w2305, IN16[7], w2403, w2404);
  FullAdder U310 (w2404, w2307, IN17[7], w2405, w2406);
  FullAdder U311 (w2406, w2309, IN18[7], w2407, w2408);
  FullAdder U312 (w2408, w2311, IN19[7], w2409, w2410);
  FullAdder U313 (w2410, w2313, IN20[7], w2411, w2412);
  FullAdder U314 (w2412, w2315, IN21[7], w2413, w2414);
  FullAdder U315 (w2414, w2317, IN22[7], w2415, w2416);
  FullAdder U316 (w2416, w2319, IN23[7], w2417, w2418);
  FullAdder U317 (w2418, w2321, IN24[7], w2419, w2420);
  FullAdder U318 (w2420, w2323, IN25[7], w2421, w2422);
  FullAdder U319 (w2422, w2325, IN26[7], w2423, w2424);
  FullAdder U320 (w2424, w2327, IN27[7], w2425, w2426);
  FullAdder U321 (w2426, w2329, IN28[7], w2427, w2428);
  FullAdder U322 (w2428, w2331, IN29[7], w2429, w2430);
  FullAdder U323 (w2430, w2333, IN30[7], w2431, w2432);
  FullAdder U324 (w2432, w2335, IN31[7], w2433, w2434);
  FullAdder U325 (w2434, w2337, IN32[7], w2435, w2436);
  FullAdder U326 (w2436, w2339, IN33[7], w2437, w2438);
  FullAdder U327 (w2438, w2341, IN34[7], w2439, w2440);
  FullAdder U328 (w2440, w2343, IN35[7], w2441, w2442);
  FullAdder U329 (w2442, w2345, IN36[7], w2443, w2444);
  FullAdder U330 (w2444, w2347, IN37[7], w2445, w2446);
  FullAdder U331 (w2446, w2349, IN38[7], w2447, w2448);
  FullAdder U332 (w2448, w2351, IN39[7], w2449, w2450);
  FullAdder U333 (w2450, w2353, IN40[7], w2451, w2452);
  FullAdder U334 (w2452, w2355, IN41[7], w2453, w2454);
  FullAdder U335 (w2454, w2357, IN42[7], w2455, w2456);
  FullAdder U336 (w2456, w2359, IN43[7], w2457, w2458);
  FullAdder U337 (w2458, w2361, IN44[7], w2459, w2460);
  FullAdder U338 (w2460, w2363, IN45[7], w2461, w2462);
  FullAdder U339 (w2462, w2365, IN46[7], w2463, w2464);
  FullAdder U340 (w2464, w2367, IN47[7], w2465, w2466);
  FullAdder U341 (w2466, w2369, IN48[7], w2467, w2468);
  FullAdder U342 (w2468, w2371, IN49[7], w2469, w2470);
  FullAdder U343 (w2470, w2373, IN50[7], w2471, w2472);
  FullAdder U344 (w2472, w2375, IN51[5], w2473, w2474);
  FullAdder U345 (w2474, w2377, IN52[4], w2475, w2476);
  FullAdder U346 (w2476, w2379, IN53[3], w2477, w2478);
  FullAdder U347 (w2478, w2381, IN54[2], w2479, w2480);
  FullAdder U348 (w2480, w2383, IN55[1], w2481, w2482);
  FullAdder U349 (w2482, w2384, IN56[0], w2483, w2484);
  HalfAdder U350 (w2387, IN8[8], Out1[8], w2486);
  FullAdder U351 (w2486, w2389, IN9[8], w2487, w2488);
  FullAdder U352 (w2488, w2391, IN10[8], w2489, w2490);
  FullAdder U353 (w2490, w2393, IN11[8], w2491, w2492);
  FullAdder U354 (w2492, w2395, IN12[8], w2493, w2494);
  FullAdder U355 (w2494, w2397, IN13[8], w2495, w2496);
  FullAdder U356 (w2496, w2399, IN14[8], w2497, w2498);
  FullAdder U357 (w2498, w2401, IN15[8], w2499, w2500);
  FullAdder U358 (w2500, w2403, IN16[8], w2501, w2502);
  FullAdder U359 (w2502, w2405, IN17[8], w2503, w2504);
  FullAdder U360 (w2504, w2407, IN18[8], w2505, w2506);
  FullAdder U361 (w2506, w2409, IN19[8], w2507, w2508);
  FullAdder U362 (w2508, w2411, IN20[8], w2509, w2510);
  FullAdder U363 (w2510, w2413, IN21[8], w2511, w2512);
  FullAdder U364 (w2512, w2415, IN22[8], w2513, w2514);
  FullAdder U365 (w2514, w2417, IN23[8], w2515, w2516);
  FullAdder U366 (w2516, w2419, IN24[8], w2517, w2518);
  FullAdder U367 (w2518, w2421, IN25[8], w2519, w2520);
  FullAdder U368 (w2520, w2423, IN26[8], w2521, w2522);
  FullAdder U369 (w2522, w2425, IN27[8], w2523, w2524);
  FullAdder U370 (w2524, w2427, IN28[8], w2525, w2526);
  FullAdder U371 (w2526, w2429, IN29[8], w2527, w2528);
  FullAdder U372 (w2528, w2431, IN30[8], w2529, w2530);
  FullAdder U373 (w2530, w2433, IN31[8], w2531, w2532);
  FullAdder U374 (w2532, w2435, IN32[8], w2533, w2534);
  FullAdder U375 (w2534, w2437, IN33[8], w2535, w2536);
  FullAdder U376 (w2536, w2439, IN34[8], w2537, w2538);
  FullAdder U377 (w2538, w2441, IN35[8], w2539, w2540);
  FullAdder U378 (w2540, w2443, IN36[8], w2541, w2542);
  FullAdder U379 (w2542, w2445, IN37[8], w2543, w2544);
  FullAdder U380 (w2544, w2447, IN38[8], w2545, w2546);
  FullAdder U381 (w2546, w2449, IN39[8], w2547, w2548);
  FullAdder U382 (w2548, w2451, IN40[8], w2549, w2550);
  FullAdder U383 (w2550, w2453, IN41[8], w2551, w2552);
  FullAdder U384 (w2552, w2455, IN42[8], w2553, w2554);
  FullAdder U385 (w2554, w2457, IN43[8], w2555, w2556);
  FullAdder U386 (w2556, w2459, IN44[8], w2557, w2558);
  FullAdder U387 (w2558, w2461, IN45[8], w2559, w2560);
  FullAdder U388 (w2560, w2463, IN46[8], w2561, w2562);
  FullAdder U389 (w2562, w2465, IN47[8], w2563, w2564);
  FullAdder U390 (w2564, w2467, IN48[8], w2565, w2566);
  FullAdder U391 (w2566, w2469, IN49[8], w2567, w2568);
  FullAdder U392 (w2568, w2471, IN50[8], w2569, w2570);
  FullAdder U393 (w2570, w2473, IN51[6], w2571, w2572);
  FullAdder U394 (w2572, w2475, IN52[5], w2573, w2574);
  FullAdder U395 (w2574, w2477, IN53[4], w2575, w2576);
  FullAdder U396 (w2576, w2479, IN54[3], w2577, w2578);
  FullAdder U397 (w2578, w2481, IN55[2], w2579, w2580);
  FullAdder U398 (w2580, w2483, IN56[1], w2581, w2582);
  FullAdder U399 (w2582, w2484, IN57[0], w2583, w2584);
  HalfAdder U400 (w2487, IN9[9], Out1[9], w2586);
  FullAdder U401 (w2586, w2489, IN10[9], w2587, w2588);
  FullAdder U402 (w2588, w2491, IN11[9], w2589, w2590);
  FullAdder U403 (w2590, w2493, IN12[9], w2591, w2592);
  FullAdder U404 (w2592, w2495, IN13[9], w2593, w2594);
  FullAdder U405 (w2594, w2497, IN14[9], w2595, w2596);
  FullAdder U406 (w2596, w2499, IN15[9], w2597, w2598);
  FullAdder U407 (w2598, w2501, IN16[9], w2599, w2600);
  FullAdder U408 (w2600, w2503, IN17[9], w2601, w2602);
  FullAdder U409 (w2602, w2505, IN18[9], w2603, w2604);
  FullAdder U410 (w2604, w2507, IN19[9], w2605, w2606);
  FullAdder U411 (w2606, w2509, IN20[9], w2607, w2608);
  FullAdder U412 (w2608, w2511, IN21[9], w2609, w2610);
  FullAdder U413 (w2610, w2513, IN22[9], w2611, w2612);
  FullAdder U414 (w2612, w2515, IN23[9], w2613, w2614);
  FullAdder U415 (w2614, w2517, IN24[9], w2615, w2616);
  FullAdder U416 (w2616, w2519, IN25[9], w2617, w2618);
  FullAdder U417 (w2618, w2521, IN26[9], w2619, w2620);
  FullAdder U418 (w2620, w2523, IN27[9], w2621, w2622);
  FullAdder U419 (w2622, w2525, IN28[9], w2623, w2624);
  FullAdder U420 (w2624, w2527, IN29[9], w2625, w2626);
  FullAdder U421 (w2626, w2529, IN30[9], w2627, w2628);
  FullAdder U422 (w2628, w2531, IN31[9], w2629, w2630);
  FullAdder U423 (w2630, w2533, IN32[9], w2631, w2632);
  FullAdder U424 (w2632, w2535, IN33[9], w2633, w2634);
  FullAdder U425 (w2634, w2537, IN34[9], w2635, w2636);
  FullAdder U426 (w2636, w2539, IN35[9], w2637, w2638);
  FullAdder U427 (w2638, w2541, IN36[9], w2639, w2640);
  FullAdder U428 (w2640, w2543, IN37[9], w2641, w2642);
  FullAdder U429 (w2642, w2545, IN38[9], w2643, w2644);
  FullAdder U430 (w2644, w2547, IN39[9], w2645, w2646);
  FullAdder U431 (w2646, w2549, IN40[9], w2647, w2648);
  FullAdder U432 (w2648, w2551, IN41[9], w2649, w2650);
  FullAdder U433 (w2650, w2553, IN42[9], w2651, w2652);
  FullAdder U434 (w2652, w2555, IN43[9], w2653, w2654);
  FullAdder U435 (w2654, w2557, IN44[9], w2655, w2656);
  FullAdder U436 (w2656, w2559, IN45[9], w2657, w2658);
  FullAdder U437 (w2658, w2561, IN46[9], w2659, w2660);
  FullAdder U438 (w2660, w2563, IN47[9], w2661, w2662);
  FullAdder U439 (w2662, w2565, IN48[9], w2663, w2664);
  FullAdder U440 (w2664, w2567, IN49[9], w2665, w2666);
  FullAdder U441 (w2666, w2569, IN50[9], w2667, w2668);
  FullAdder U442 (w2668, w2571, IN51[7], w2669, w2670);
  FullAdder U443 (w2670, w2573, IN52[6], w2671, w2672);
  FullAdder U444 (w2672, w2575, IN53[5], w2673, w2674);
  FullAdder U445 (w2674, w2577, IN54[4], w2675, w2676);
  FullAdder U446 (w2676, w2579, IN55[3], w2677, w2678);
  FullAdder U447 (w2678, w2581, IN56[2], w2679, w2680);
  FullAdder U448 (w2680, w2583, IN57[1], w2681, w2682);
  FullAdder U449 (w2682, w2584, IN58[0], w2683, w2684);
  HalfAdder U450 (w2587, IN10[10], Out1[10], w2686);
  FullAdder U451 (w2686, w2589, IN11[10], w2687, w2688);
  FullAdder U452 (w2688, w2591, IN12[10], w2689, w2690);
  FullAdder U453 (w2690, w2593, IN13[10], w2691, w2692);
  FullAdder U454 (w2692, w2595, IN14[10], w2693, w2694);
  FullAdder U455 (w2694, w2597, IN15[10], w2695, w2696);
  FullAdder U456 (w2696, w2599, IN16[10], w2697, w2698);
  FullAdder U457 (w2698, w2601, IN17[10], w2699, w2700);
  FullAdder U458 (w2700, w2603, IN18[10], w2701, w2702);
  FullAdder U459 (w2702, w2605, IN19[10], w2703, w2704);
  FullAdder U460 (w2704, w2607, IN20[10], w2705, w2706);
  FullAdder U461 (w2706, w2609, IN21[10], w2707, w2708);
  FullAdder U462 (w2708, w2611, IN22[10], w2709, w2710);
  FullAdder U463 (w2710, w2613, IN23[10], w2711, w2712);
  FullAdder U464 (w2712, w2615, IN24[10], w2713, w2714);
  FullAdder U465 (w2714, w2617, IN25[10], w2715, w2716);
  FullAdder U466 (w2716, w2619, IN26[10], w2717, w2718);
  FullAdder U467 (w2718, w2621, IN27[10], w2719, w2720);
  FullAdder U468 (w2720, w2623, IN28[10], w2721, w2722);
  FullAdder U469 (w2722, w2625, IN29[10], w2723, w2724);
  FullAdder U470 (w2724, w2627, IN30[10], w2725, w2726);
  FullAdder U471 (w2726, w2629, IN31[10], w2727, w2728);
  FullAdder U472 (w2728, w2631, IN32[10], w2729, w2730);
  FullAdder U473 (w2730, w2633, IN33[10], w2731, w2732);
  FullAdder U474 (w2732, w2635, IN34[10], w2733, w2734);
  FullAdder U475 (w2734, w2637, IN35[10], w2735, w2736);
  FullAdder U476 (w2736, w2639, IN36[10], w2737, w2738);
  FullAdder U477 (w2738, w2641, IN37[10], w2739, w2740);
  FullAdder U478 (w2740, w2643, IN38[10], w2741, w2742);
  FullAdder U479 (w2742, w2645, IN39[10], w2743, w2744);
  FullAdder U480 (w2744, w2647, IN40[10], w2745, w2746);
  FullAdder U481 (w2746, w2649, IN41[10], w2747, w2748);
  FullAdder U482 (w2748, w2651, IN42[10], w2749, w2750);
  FullAdder U483 (w2750, w2653, IN43[10], w2751, w2752);
  FullAdder U484 (w2752, w2655, IN44[10], w2753, w2754);
  FullAdder U485 (w2754, w2657, IN45[10], w2755, w2756);
  FullAdder U486 (w2756, w2659, IN46[10], w2757, w2758);
  FullAdder U487 (w2758, w2661, IN47[10], w2759, w2760);
  FullAdder U488 (w2760, w2663, IN48[10], w2761, w2762);
  FullAdder U489 (w2762, w2665, IN49[10], w2763, w2764);
  FullAdder U490 (w2764, w2667, IN50[10], w2765, w2766);
  FullAdder U491 (w2766, w2669, IN51[8], w2767, w2768);
  FullAdder U492 (w2768, w2671, IN52[7], w2769, w2770);
  FullAdder U493 (w2770, w2673, IN53[6], w2771, w2772);
  FullAdder U494 (w2772, w2675, IN54[5], w2773, w2774);
  FullAdder U495 (w2774, w2677, IN55[4], w2775, w2776);
  FullAdder U496 (w2776, w2679, IN56[3], w2777, w2778);
  FullAdder U497 (w2778, w2681, IN57[2], w2779, w2780);
  FullAdder U498 (w2780, w2683, IN58[1], w2781, w2782);
  FullAdder U499 (w2782, w2684, IN59[0], w2783, w2784);
  HalfAdder U500 (w2687, IN11[11], Out1[11], w2786);
  FullAdder U501 (w2786, w2689, IN12[11], w2787, w2788);
  FullAdder U502 (w2788, w2691, IN13[11], w2789, w2790);
  FullAdder U503 (w2790, w2693, IN14[11], w2791, w2792);
  FullAdder U504 (w2792, w2695, IN15[11], w2793, w2794);
  FullAdder U505 (w2794, w2697, IN16[11], w2795, w2796);
  FullAdder U506 (w2796, w2699, IN17[11], w2797, w2798);
  FullAdder U507 (w2798, w2701, IN18[11], w2799, w2800);
  FullAdder U508 (w2800, w2703, IN19[11], w2801, w2802);
  FullAdder U509 (w2802, w2705, IN20[11], w2803, w2804);
  FullAdder U510 (w2804, w2707, IN21[11], w2805, w2806);
  FullAdder U511 (w2806, w2709, IN22[11], w2807, w2808);
  FullAdder U512 (w2808, w2711, IN23[11], w2809, w2810);
  FullAdder U513 (w2810, w2713, IN24[11], w2811, w2812);
  FullAdder U514 (w2812, w2715, IN25[11], w2813, w2814);
  FullAdder U515 (w2814, w2717, IN26[11], w2815, w2816);
  FullAdder U516 (w2816, w2719, IN27[11], w2817, w2818);
  FullAdder U517 (w2818, w2721, IN28[11], w2819, w2820);
  FullAdder U518 (w2820, w2723, IN29[11], w2821, w2822);
  FullAdder U519 (w2822, w2725, IN30[11], w2823, w2824);
  FullAdder U520 (w2824, w2727, IN31[11], w2825, w2826);
  FullAdder U521 (w2826, w2729, IN32[11], w2827, w2828);
  FullAdder U522 (w2828, w2731, IN33[11], w2829, w2830);
  FullAdder U523 (w2830, w2733, IN34[11], w2831, w2832);
  FullAdder U524 (w2832, w2735, IN35[11], w2833, w2834);
  FullAdder U525 (w2834, w2737, IN36[11], w2835, w2836);
  FullAdder U526 (w2836, w2739, IN37[11], w2837, w2838);
  FullAdder U527 (w2838, w2741, IN38[11], w2839, w2840);
  FullAdder U528 (w2840, w2743, IN39[11], w2841, w2842);
  FullAdder U529 (w2842, w2745, IN40[11], w2843, w2844);
  FullAdder U530 (w2844, w2747, IN41[11], w2845, w2846);
  FullAdder U531 (w2846, w2749, IN42[11], w2847, w2848);
  FullAdder U532 (w2848, w2751, IN43[11], w2849, w2850);
  FullAdder U533 (w2850, w2753, IN44[11], w2851, w2852);
  FullAdder U534 (w2852, w2755, IN45[11], w2853, w2854);
  FullAdder U535 (w2854, w2757, IN46[11], w2855, w2856);
  FullAdder U536 (w2856, w2759, IN47[11], w2857, w2858);
  FullAdder U537 (w2858, w2761, IN48[11], w2859, w2860);
  FullAdder U538 (w2860, w2763, IN49[11], w2861, w2862);
  FullAdder U539 (w2862, w2765, IN50[11], w2863, w2864);
  FullAdder U540 (w2864, w2767, IN51[9], w2865, w2866);
  FullAdder U541 (w2866, w2769, IN52[8], w2867, w2868);
  FullAdder U542 (w2868, w2771, IN53[7], w2869, w2870);
  FullAdder U543 (w2870, w2773, IN54[6], w2871, w2872);
  FullAdder U544 (w2872, w2775, IN55[5], w2873, w2874);
  FullAdder U545 (w2874, w2777, IN56[4], w2875, w2876);
  FullAdder U546 (w2876, w2779, IN57[3], w2877, w2878);
  FullAdder U547 (w2878, w2781, IN58[2], w2879, w2880);
  FullAdder U548 (w2880, w2783, IN59[1], w2881, w2882);
  FullAdder U549 (w2882, w2784, IN60[0], w2883, w2884);
  HalfAdder U550 (w2787, IN12[12], Out1[12], w2886);
  FullAdder U551 (w2886, w2789, IN13[12], w2887, w2888);
  FullAdder U552 (w2888, w2791, IN14[12], w2889, w2890);
  FullAdder U553 (w2890, w2793, IN15[12], w2891, w2892);
  FullAdder U554 (w2892, w2795, IN16[12], w2893, w2894);
  FullAdder U555 (w2894, w2797, IN17[12], w2895, w2896);
  FullAdder U556 (w2896, w2799, IN18[12], w2897, w2898);
  FullAdder U557 (w2898, w2801, IN19[12], w2899, w2900);
  FullAdder U558 (w2900, w2803, IN20[12], w2901, w2902);
  FullAdder U559 (w2902, w2805, IN21[12], w2903, w2904);
  FullAdder U560 (w2904, w2807, IN22[12], w2905, w2906);
  FullAdder U561 (w2906, w2809, IN23[12], w2907, w2908);
  FullAdder U562 (w2908, w2811, IN24[12], w2909, w2910);
  FullAdder U563 (w2910, w2813, IN25[12], w2911, w2912);
  FullAdder U564 (w2912, w2815, IN26[12], w2913, w2914);
  FullAdder U565 (w2914, w2817, IN27[12], w2915, w2916);
  FullAdder U566 (w2916, w2819, IN28[12], w2917, w2918);
  FullAdder U567 (w2918, w2821, IN29[12], w2919, w2920);
  FullAdder U568 (w2920, w2823, IN30[12], w2921, w2922);
  FullAdder U569 (w2922, w2825, IN31[12], w2923, w2924);
  FullAdder U570 (w2924, w2827, IN32[12], w2925, w2926);
  FullAdder U571 (w2926, w2829, IN33[12], w2927, w2928);
  FullAdder U572 (w2928, w2831, IN34[12], w2929, w2930);
  FullAdder U573 (w2930, w2833, IN35[12], w2931, w2932);
  FullAdder U574 (w2932, w2835, IN36[12], w2933, w2934);
  FullAdder U575 (w2934, w2837, IN37[12], w2935, w2936);
  FullAdder U576 (w2936, w2839, IN38[12], w2937, w2938);
  FullAdder U577 (w2938, w2841, IN39[12], w2939, w2940);
  FullAdder U578 (w2940, w2843, IN40[12], w2941, w2942);
  FullAdder U579 (w2942, w2845, IN41[12], w2943, w2944);
  FullAdder U580 (w2944, w2847, IN42[12], w2945, w2946);
  FullAdder U581 (w2946, w2849, IN43[12], w2947, w2948);
  FullAdder U582 (w2948, w2851, IN44[12], w2949, w2950);
  FullAdder U583 (w2950, w2853, IN45[12], w2951, w2952);
  FullAdder U584 (w2952, w2855, IN46[12], w2953, w2954);
  FullAdder U585 (w2954, w2857, IN47[12], w2955, w2956);
  FullAdder U586 (w2956, w2859, IN48[12], w2957, w2958);
  FullAdder U587 (w2958, w2861, IN49[12], w2959, w2960);
  FullAdder U588 (w2960, w2863, IN50[12], w2961, w2962);
  FullAdder U589 (w2962, w2865, IN51[10], w2963, w2964);
  FullAdder U590 (w2964, w2867, IN52[9], w2965, w2966);
  FullAdder U591 (w2966, w2869, IN53[8], w2967, w2968);
  FullAdder U592 (w2968, w2871, IN54[7], w2969, w2970);
  FullAdder U593 (w2970, w2873, IN55[6], w2971, w2972);
  FullAdder U594 (w2972, w2875, IN56[5], w2973, w2974);
  FullAdder U595 (w2974, w2877, IN57[4], w2975, w2976);
  FullAdder U596 (w2976, w2879, IN58[3], w2977, w2978);
  FullAdder U597 (w2978, w2881, IN59[2], w2979, w2980);
  FullAdder U598 (w2980, w2883, IN60[1], w2981, w2982);
  FullAdder U599 (w2982, w2884, IN61[0], w2983, w2984);
  HalfAdder U600 (w2887, IN13[13], Out1[13], w2986);
  FullAdder U601 (w2986, w2889, IN14[13], w2987, w2988);
  FullAdder U602 (w2988, w2891, IN15[13], w2989, w2990);
  FullAdder U603 (w2990, w2893, IN16[13], w2991, w2992);
  FullAdder U604 (w2992, w2895, IN17[13], w2993, w2994);
  FullAdder U605 (w2994, w2897, IN18[13], w2995, w2996);
  FullAdder U606 (w2996, w2899, IN19[13], w2997, w2998);
  FullAdder U607 (w2998, w2901, IN20[13], w2999, w3000);
  FullAdder U608 (w3000, w2903, IN21[13], w3001, w3002);
  FullAdder U609 (w3002, w2905, IN22[13], w3003, w3004);
  FullAdder U610 (w3004, w2907, IN23[13], w3005, w3006);
  FullAdder U611 (w3006, w2909, IN24[13], w3007, w3008);
  FullAdder U612 (w3008, w2911, IN25[13], w3009, w3010);
  FullAdder U613 (w3010, w2913, IN26[13], w3011, w3012);
  FullAdder U614 (w3012, w2915, IN27[13], w3013, w3014);
  FullAdder U615 (w3014, w2917, IN28[13], w3015, w3016);
  FullAdder U616 (w3016, w2919, IN29[13], w3017, w3018);
  FullAdder U617 (w3018, w2921, IN30[13], w3019, w3020);
  FullAdder U618 (w3020, w2923, IN31[13], w3021, w3022);
  FullAdder U619 (w3022, w2925, IN32[13], w3023, w3024);
  FullAdder U620 (w3024, w2927, IN33[13], w3025, w3026);
  FullAdder U621 (w3026, w2929, IN34[13], w3027, w3028);
  FullAdder U622 (w3028, w2931, IN35[13], w3029, w3030);
  FullAdder U623 (w3030, w2933, IN36[13], w3031, w3032);
  FullAdder U624 (w3032, w2935, IN37[13], w3033, w3034);
  FullAdder U625 (w3034, w2937, IN38[13], w3035, w3036);
  FullAdder U626 (w3036, w2939, IN39[13], w3037, w3038);
  FullAdder U627 (w3038, w2941, IN40[13], w3039, w3040);
  FullAdder U628 (w3040, w2943, IN41[13], w3041, w3042);
  FullAdder U629 (w3042, w2945, IN42[13], w3043, w3044);
  FullAdder U630 (w3044, w2947, IN43[13], w3045, w3046);
  FullAdder U631 (w3046, w2949, IN44[13], w3047, w3048);
  FullAdder U632 (w3048, w2951, IN45[13], w3049, w3050);
  FullAdder U633 (w3050, w2953, IN46[13], w3051, w3052);
  FullAdder U634 (w3052, w2955, IN47[13], w3053, w3054);
  FullAdder U635 (w3054, w2957, IN48[13], w3055, w3056);
  FullAdder U636 (w3056, w2959, IN49[13], w3057, w3058);
  FullAdder U637 (w3058, w2961, IN50[13], w3059, w3060);
  FullAdder U638 (w3060, w2963, IN51[11], w3061, w3062);
  FullAdder U639 (w3062, w2965, IN52[10], w3063, w3064);
  FullAdder U640 (w3064, w2967, IN53[9], w3065, w3066);
  FullAdder U641 (w3066, w2969, IN54[8], w3067, w3068);
  FullAdder U642 (w3068, w2971, IN55[7], w3069, w3070);
  FullAdder U643 (w3070, w2973, IN56[6], w3071, w3072);
  FullAdder U644 (w3072, w2975, IN57[5], w3073, w3074);
  FullAdder U645 (w3074, w2977, IN58[4], w3075, w3076);
  FullAdder U646 (w3076, w2979, IN59[3], w3077, w3078);
  FullAdder U647 (w3078, w2981, IN60[2], w3079, w3080);
  FullAdder U648 (w3080, w2983, IN61[1], w3081, w3082);
  FullAdder U649 (w3082, w2984, IN62[0], w3083, w3084);
  HalfAdder U650 (w2987, IN14[14], Out1[14], w3086);
  FullAdder U651 (w3086, w2989, IN15[14], w3087, w3088);
  FullAdder U652 (w3088, w2991, IN16[14], w3089, w3090);
  FullAdder U653 (w3090, w2993, IN17[14], w3091, w3092);
  FullAdder U654 (w3092, w2995, IN18[14], w3093, w3094);
  FullAdder U655 (w3094, w2997, IN19[14], w3095, w3096);
  FullAdder U656 (w3096, w2999, IN20[14], w3097, w3098);
  FullAdder U657 (w3098, w3001, IN21[14], w3099, w3100);
  FullAdder U658 (w3100, w3003, IN22[14], w3101, w3102);
  FullAdder U659 (w3102, w3005, IN23[14], w3103, w3104);
  FullAdder U660 (w3104, w3007, IN24[14], w3105, w3106);
  FullAdder U661 (w3106, w3009, IN25[14], w3107, w3108);
  FullAdder U662 (w3108, w3011, IN26[14], w3109, w3110);
  FullAdder U663 (w3110, w3013, IN27[14], w3111, w3112);
  FullAdder U664 (w3112, w3015, IN28[14], w3113, w3114);
  FullAdder U665 (w3114, w3017, IN29[14], w3115, w3116);
  FullAdder U666 (w3116, w3019, IN30[14], w3117, w3118);
  FullAdder U667 (w3118, w3021, IN31[14], w3119, w3120);
  FullAdder U668 (w3120, w3023, IN32[14], w3121, w3122);
  FullAdder U669 (w3122, w3025, IN33[14], w3123, w3124);
  FullAdder U670 (w3124, w3027, IN34[14], w3125, w3126);
  FullAdder U671 (w3126, w3029, IN35[14], w3127, w3128);
  FullAdder U672 (w3128, w3031, IN36[14], w3129, w3130);
  FullAdder U673 (w3130, w3033, IN37[14], w3131, w3132);
  FullAdder U674 (w3132, w3035, IN38[14], w3133, w3134);
  FullAdder U675 (w3134, w3037, IN39[14], w3135, w3136);
  FullAdder U676 (w3136, w3039, IN40[14], w3137, w3138);
  FullAdder U677 (w3138, w3041, IN41[14], w3139, w3140);
  FullAdder U678 (w3140, w3043, IN42[14], w3141, w3142);
  FullAdder U679 (w3142, w3045, IN43[14], w3143, w3144);
  FullAdder U680 (w3144, w3047, IN44[14], w3145, w3146);
  FullAdder U681 (w3146, w3049, IN45[14], w3147, w3148);
  FullAdder U682 (w3148, w3051, IN46[14], w3149, w3150);
  FullAdder U683 (w3150, w3053, IN47[14], w3151, w3152);
  FullAdder U684 (w3152, w3055, IN48[14], w3153, w3154);
  FullAdder U685 (w3154, w3057, IN49[14], w3155, w3156);
  FullAdder U686 (w3156, w3059, IN50[14], w3157, w3158);
  FullAdder U687 (w3158, w3061, IN51[12], w3159, w3160);
  FullAdder U688 (w3160, w3063, IN52[11], w3161, w3162);
  FullAdder U689 (w3162, w3065, IN53[10], w3163, w3164);
  FullAdder U690 (w3164, w3067, IN54[9], w3165, w3166);
  FullAdder U691 (w3166, w3069, IN55[8], w3167, w3168);
  FullAdder U692 (w3168, w3071, IN56[7], w3169, w3170);
  FullAdder U693 (w3170, w3073, IN57[6], w3171, w3172);
  FullAdder U694 (w3172, w3075, IN58[5], w3173, w3174);
  FullAdder U695 (w3174, w3077, IN59[4], w3175, w3176);
  FullAdder U696 (w3176, w3079, IN60[3], w3177, w3178);
  FullAdder U697 (w3178, w3081, IN61[2], w3179, w3180);
  FullAdder U698 (w3180, w3083, IN62[1], w3181, w3182);
  FullAdder U699 (w3182, w3084, IN63[0], w3183, w3184);
  HalfAdder U700 (w3087, IN15[15], Out1[15], w3186);
  FullAdder U701 (w3186, w3089, IN16[15], w3187, w3188);
  FullAdder U702 (w3188, w3091, IN17[15], w3189, w3190);
  FullAdder U703 (w3190, w3093, IN18[15], w3191, w3192);
  FullAdder U704 (w3192, w3095, IN19[15], w3193, w3194);
  FullAdder U705 (w3194, w3097, IN20[15], w3195, w3196);
  FullAdder U706 (w3196, w3099, IN21[15], w3197, w3198);
  FullAdder U707 (w3198, w3101, IN22[15], w3199, w3200);
  FullAdder U708 (w3200, w3103, IN23[15], w3201, w3202);
  FullAdder U709 (w3202, w3105, IN24[15], w3203, w3204);
  FullAdder U710 (w3204, w3107, IN25[15], w3205, w3206);
  FullAdder U711 (w3206, w3109, IN26[15], w3207, w3208);
  FullAdder U712 (w3208, w3111, IN27[15], w3209, w3210);
  FullAdder U713 (w3210, w3113, IN28[15], w3211, w3212);
  FullAdder U714 (w3212, w3115, IN29[15], w3213, w3214);
  FullAdder U715 (w3214, w3117, IN30[15], w3215, w3216);
  FullAdder U716 (w3216, w3119, IN31[15], w3217, w3218);
  FullAdder U717 (w3218, w3121, IN32[15], w3219, w3220);
  FullAdder U718 (w3220, w3123, IN33[15], w3221, w3222);
  FullAdder U719 (w3222, w3125, IN34[15], w3223, w3224);
  FullAdder U720 (w3224, w3127, IN35[15], w3225, w3226);
  FullAdder U721 (w3226, w3129, IN36[15], w3227, w3228);
  FullAdder U722 (w3228, w3131, IN37[15], w3229, w3230);
  FullAdder U723 (w3230, w3133, IN38[15], w3231, w3232);
  FullAdder U724 (w3232, w3135, IN39[15], w3233, w3234);
  FullAdder U725 (w3234, w3137, IN40[15], w3235, w3236);
  FullAdder U726 (w3236, w3139, IN41[15], w3237, w3238);
  FullAdder U727 (w3238, w3141, IN42[15], w3239, w3240);
  FullAdder U728 (w3240, w3143, IN43[15], w3241, w3242);
  FullAdder U729 (w3242, w3145, IN44[15], w3243, w3244);
  FullAdder U730 (w3244, w3147, IN45[15], w3245, w3246);
  FullAdder U731 (w3246, w3149, IN46[15], w3247, w3248);
  FullAdder U732 (w3248, w3151, IN47[15], w3249, w3250);
  FullAdder U733 (w3250, w3153, IN48[15], w3251, w3252);
  FullAdder U734 (w3252, w3155, IN49[15], w3253, w3254);
  FullAdder U735 (w3254, w3157, IN50[15], w3255, w3256);
  FullAdder U736 (w3256, w3159, IN51[13], w3257, w3258);
  FullAdder U737 (w3258, w3161, IN52[12], w3259, w3260);
  FullAdder U738 (w3260, w3163, IN53[11], w3261, w3262);
  FullAdder U739 (w3262, w3165, IN54[10], w3263, w3264);
  FullAdder U740 (w3264, w3167, IN55[9], w3265, w3266);
  FullAdder U741 (w3266, w3169, IN56[8], w3267, w3268);
  FullAdder U742 (w3268, w3171, IN57[7], w3269, w3270);
  FullAdder U743 (w3270, w3173, IN58[6], w3271, w3272);
  FullAdder U744 (w3272, w3175, IN59[5], w3273, w3274);
  FullAdder U745 (w3274, w3177, IN60[4], w3275, w3276);
  FullAdder U746 (w3276, w3179, IN61[3], w3277, w3278);
  FullAdder U747 (w3278, w3181, IN62[2], w3279, w3280);
  FullAdder U748 (w3280, w3183, IN63[1], w3281, w3282);
  FullAdder U749 (w3282, w3184, IN64[0], w3283, w3284);
  HalfAdder U750 (w3187, IN16[16], Out1[16], w3286);
  FullAdder U751 (w3286, w3189, IN17[16], w3287, w3288);
  FullAdder U752 (w3288, w3191, IN18[16], w3289, w3290);
  FullAdder U753 (w3290, w3193, IN19[16], w3291, w3292);
  FullAdder U754 (w3292, w3195, IN20[16], w3293, w3294);
  FullAdder U755 (w3294, w3197, IN21[16], w3295, w3296);
  FullAdder U756 (w3296, w3199, IN22[16], w3297, w3298);
  FullAdder U757 (w3298, w3201, IN23[16], w3299, w3300);
  FullAdder U758 (w3300, w3203, IN24[16], w3301, w3302);
  FullAdder U759 (w3302, w3205, IN25[16], w3303, w3304);
  FullAdder U760 (w3304, w3207, IN26[16], w3305, w3306);
  FullAdder U761 (w3306, w3209, IN27[16], w3307, w3308);
  FullAdder U762 (w3308, w3211, IN28[16], w3309, w3310);
  FullAdder U763 (w3310, w3213, IN29[16], w3311, w3312);
  FullAdder U764 (w3312, w3215, IN30[16], w3313, w3314);
  FullAdder U765 (w3314, w3217, IN31[16], w3315, w3316);
  FullAdder U766 (w3316, w3219, IN32[16], w3317, w3318);
  FullAdder U767 (w3318, w3221, IN33[16], w3319, w3320);
  FullAdder U768 (w3320, w3223, IN34[16], w3321, w3322);
  FullAdder U769 (w3322, w3225, IN35[16], w3323, w3324);
  FullAdder U770 (w3324, w3227, IN36[16], w3325, w3326);
  FullAdder U771 (w3326, w3229, IN37[16], w3327, w3328);
  FullAdder U772 (w3328, w3231, IN38[16], w3329, w3330);
  FullAdder U773 (w3330, w3233, IN39[16], w3331, w3332);
  FullAdder U774 (w3332, w3235, IN40[16], w3333, w3334);
  FullAdder U775 (w3334, w3237, IN41[16], w3335, w3336);
  FullAdder U776 (w3336, w3239, IN42[16], w3337, w3338);
  FullAdder U777 (w3338, w3241, IN43[16], w3339, w3340);
  FullAdder U778 (w3340, w3243, IN44[16], w3341, w3342);
  FullAdder U779 (w3342, w3245, IN45[16], w3343, w3344);
  FullAdder U780 (w3344, w3247, IN46[16], w3345, w3346);
  FullAdder U781 (w3346, w3249, IN47[16], w3347, w3348);
  FullAdder U782 (w3348, w3251, IN48[16], w3349, w3350);
  FullAdder U783 (w3350, w3253, IN49[16], w3351, w3352);
  FullAdder U784 (w3352, w3255, IN50[16], w3353, w3354);
  FullAdder U785 (w3354, w3257, IN51[14], w3355, w3356);
  FullAdder U786 (w3356, w3259, IN52[13], w3357, w3358);
  FullAdder U787 (w3358, w3261, IN53[12], w3359, w3360);
  FullAdder U788 (w3360, w3263, IN54[11], w3361, w3362);
  FullAdder U789 (w3362, w3265, IN55[10], w3363, w3364);
  FullAdder U790 (w3364, w3267, IN56[9], w3365, w3366);
  FullAdder U791 (w3366, w3269, IN57[8], w3367, w3368);
  FullAdder U792 (w3368, w3271, IN58[7], w3369, w3370);
  FullAdder U793 (w3370, w3273, IN59[6], w3371, w3372);
  FullAdder U794 (w3372, w3275, IN60[5], w3373, w3374);
  FullAdder U795 (w3374, w3277, IN61[4], w3375, w3376);
  FullAdder U796 (w3376, w3279, IN62[3], w3377, w3378);
  FullAdder U797 (w3378, w3281, IN63[2], w3379, w3380);
  FullAdder U798 (w3380, w3283, IN64[1], w3381, w3382);
  FullAdder U799 (w3382, w3284, IN65[0], w3383, w3384);
  HalfAdder U800 (w3287, IN17[17], Out1[17], w3386);
  FullAdder U801 (w3386, w3289, IN18[17], w3387, w3388);
  FullAdder U802 (w3388, w3291, IN19[17], w3389, w3390);
  FullAdder U803 (w3390, w3293, IN20[17], w3391, w3392);
  FullAdder U804 (w3392, w3295, IN21[17], w3393, w3394);
  FullAdder U805 (w3394, w3297, IN22[17], w3395, w3396);
  FullAdder U806 (w3396, w3299, IN23[17], w3397, w3398);
  FullAdder U807 (w3398, w3301, IN24[17], w3399, w3400);
  FullAdder U808 (w3400, w3303, IN25[17], w3401, w3402);
  FullAdder U809 (w3402, w3305, IN26[17], w3403, w3404);
  FullAdder U810 (w3404, w3307, IN27[17], w3405, w3406);
  FullAdder U811 (w3406, w3309, IN28[17], w3407, w3408);
  FullAdder U812 (w3408, w3311, IN29[17], w3409, w3410);
  FullAdder U813 (w3410, w3313, IN30[17], w3411, w3412);
  FullAdder U814 (w3412, w3315, IN31[17], w3413, w3414);
  FullAdder U815 (w3414, w3317, IN32[17], w3415, w3416);
  FullAdder U816 (w3416, w3319, IN33[17], w3417, w3418);
  FullAdder U817 (w3418, w3321, IN34[17], w3419, w3420);
  FullAdder U818 (w3420, w3323, IN35[17], w3421, w3422);
  FullAdder U819 (w3422, w3325, IN36[17], w3423, w3424);
  FullAdder U820 (w3424, w3327, IN37[17], w3425, w3426);
  FullAdder U821 (w3426, w3329, IN38[17], w3427, w3428);
  FullAdder U822 (w3428, w3331, IN39[17], w3429, w3430);
  FullAdder U823 (w3430, w3333, IN40[17], w3431, w3432);
  FullAdder U824 (w3432, w3335, IN41[17], w3433, w3434);
  FullAdder U825 (w3434, w3337, IN42[17], w3435, w3436);
  FullAdder U826 (w3436, w3339, IN43[17], w3437, w3438);
  FullAdder U827 (w3438, w3341, IN44[17], w3439, w3440);
  FullAdder U828 (w3440, w3343, IN45[17], w3441, w3442);
  FullAdder U829 (w3442, w3345, IN46[17], w3443, w3444);
  FullAdder U830 (w3444, w3347, IN47[17], w3445, w3446);
  FullAdder U831 (w3446, w3349, IN48[17], w3447, w3448);
  FullAdder U832 (w3448, w3351, IN49[17], w3449, w3450);
  FullAdder U833 (w3450, w3353, IN50[17], w3451, w3452);
  FullAdder U834 (w3452, w3355, IN51[15], w3453, w3454);
  FullAdder U835 (w3454, w3357, IN52[14], w3455, w3456);
  FullAdder U836 (w3456, w3359, IN53[13], w3457, w3458);
  FullAdder U837 (w3458, w3361, IN54[12], w3459, w3460);
  FullAdder U838 (w3460, w3363, IN55[11], w3461, w3462);
  FullAdder U839 (w3462, w3365, IN56[10], w3463, w3464);
  FullAdder U840 (w3464, w3367, IN57[9], w3465, w3466);
  FullAdder U841 (w3466, w3369, IN58[8], w3467, w3468);
  FullAdder U842 (w3468, w3371, IN59[7], w3469, w3470);
  FullAdder U843 (w3470, w3373, IN60[6], w3471, w3472);
  FullAdder U844 (w3472, w3375, IN61[5], w3473, w3474);
  FullAdder U845 (w3474, w3377, IN62[4], w3475, w3476);
  FullAdder U846 (w3476, w3379, IN63[3], w3477, w3478);
  FullAdder U847 (w3478, w3381, IN64[2], w3479, w3480);
  FullAdder U848 (w3480, w3383, IN65[1], w3481, w3482);
  FullAdder U849 (w3482, w3384, IN66[0], w3483, w3484);
  HalfAdder U850 (w3387, IN18[18], Out1[18], w3486);
  FullAdder U851 (w3486, w3389, IN19[18], w3487, w3488);
  FullAdder U852 (w3488, w3391, IN20[18], w3489, w3490);
  FullAdder U853 (w3490, w3393, IN21[18], w3491, w3492);
  FullAdder U854 (w3492, w3395, IN22[18], w3493, w3494);
  FullAdder U855 (w3494, w3397, IN23[18], w3495, w3496);
  FullAdder U856 (w3496, w3399, IN24[18], w3497, w3498);
  FullAdder U857 (w3498, w3401, IN25[18], w3499, w3500);
  FullAdder U858 (w3500, w3403, IN26[18], w3501, w3502);
  FullAdder U859 (w3502, w3405, IN27[18], w3503, w3504);
  FullAdder U860 (w3504, w3407, IN28[18], w3505, w3506);
  FullAdder U861 (w3506, w3409, IN29[18], w3507, w3508);
  FullAdder U862 (w3508, w3411, IN30[18], w3509, w3510);
  FullAdder U863 (w3510, w3413, IN31[18], w3511, w3512);
  FullAdder U864 (w3512, w3415, IN32[18], w3513, w3514);
  FullAdder U865 (w3514, w3417, IN33[18], w3515, w3516);
  FullAdder U866 (w3516, w3419, IN34[18], w3517, w3518);
  FullAdder U867 (w3518, w3421, IN35[18], w3519, w3520);
  FullAdder U868 (w3520, w3423, IN36[18], w3521, w3522);
  FullAdder U869 (w3522, w3425, IN37[18], w3523, w3524);
  FullAdder U870 (w3524, w3427, IN38[18], w3525, w3526);
  FullAdder U871 (w3526, w3429, IN39[18], w3527, w3528);
  FullAdder U872 (w3528, w3431, IN40[18], w3529, w3530);
  FullAdder U873 (w3530, w3433, IN41[18], w3531, w3532);
  FullAdder U874 (w3532, w3435, IN42[18], w3533, w3534);
  FullAdder U875 (w3534, w3437, IN43[18], w3535, w3536);
  FullAdder U876 (w3536, w3439, IN44[18], w3537, w3538);
  FullAdder U877 (w3538, w3441, IN45[18], w3539, w3540);
  FullAdder U878 (w3540, w3443, IN46[18], w3541, w3542);
  FullAdder U879 (w3542, w3445, IN47[18], w3543, w3544);
  FullAdder U880 (w3544, w3447, IN48[18], w3545, w3546);
  FullAdder U881 (w3546, w3449, IN49[18], w3547, w3548);
  FullAdder U882 (w3548, w3451, IN50[18], w3549, w3550);
  FullAdder U883 (w3550, w3453, IN51[16], w3551, w3552);
  FullAdder U884 (w3552, w3455, IN52[15], w3553, w3554);
  FullAdder U885 (w3554, w3457, IN53[14], w3555, w3556);
  FullAdder U886 (w3556, w3459, IN54[13], w3557, w3558);
  FullAdder U887 (w3558, w3461, IN55[12], w3559, w3560);
  FullAdder U888 (w3560, w3463, IN56[11], w3561, w3562);
  FullAdder U889 (w3562, w3465, IN57[10], w3563, w3564);
  FullAdder U890 (w3564, w3467, IN58[9], w3565, w3566);
  FullAdder U891 (w3566, w3469, IN59[8], w3567, w3568);
  FullAdder U892 (w3568, w3471, IN60[7], w3569, w3570);
  FullAdder U893 (w3570, w3473, IN61[6], w3571, w3572);
  FullAdder U894 (w3572, w3475, IN62[5], w3573, w3574);
  FullAdder U895 (w3574, w3477, IN63[4], w3575, w3576);
  FullAdder U896 (w3576, w3479, IN64[3], w3577, w3578);
  FullAdder U897 (w3578, w3481, IN65[2], w3579, w3580);
  FullAdder U898 (w3580, w3483, IN66[1], w3581, w3582);
  FullAdder U899 (w3582, w3484, IN67[0], w3583, w3584);
  HalfAdder U900 (w3487, IN19[19], Out1[19], w3586);
  FullAdder U901 (w3586, w3489, IN20[19], w3587, w3588);
  FullAdder U902 (w3588, w3491, IN21[19], w3589, w3590);
  FullAdder U903 (w3590, w3493, IN22[19], w3591, w3592);
  FullAdder U904 (w3592, w3495, IN23[19], w3593, w3594);
  FullAdder U905 (w3594, w3497, IN24[19], w3595, w3596);
  FullAdder U906 (w3596, w3499, IN25[19], w3597, w3598);
  FullAdder U907 (w3598, w3501, IN26[19], w3599, w3600);
  FullAdder U908 (w3600, w3503, IN27[19], w3601, w3602);
  FullAdder U909 (w3602, w3505, IN28[19], w3603, w3604);
  FullAdder U910 (w3604, w3507, IN29[19], w3605, w3606);
  FullAdder U911 (w3606, w3509, IN30[19], w3607, w3608);
  FullAdder U912 (w3608, w3511, IN31[19], w3609, w3610);
  FullAdder U913 (w3610, w3513, IN32[19], w3611, w3612);
  FullAdder U914 (w3612, w3515, IN33[19], w3613, w3614);
  FullAdder U915 (w3614, w3517, IN34[19], w3615, w3616);
  FullAdder U916 (w3616, w3519, IN35[19], w3617, w3618);
  FullAdder U917 (w3618, w3521, IN36[19], w3619, w3620);
  FullAdder U918 (w3620, w3523, IN37[19], w3621, w3622);
  FullAdder U919 (w3622, w3525, IN38[19], w3623, w3624);
  FullAdder U920 (w3624, w3527, IN39[19], w3625, w3626);
  FullAdder U921 (w3626, w3529, IN40[19], w3627, w3628);
  FullAdder U922 (w3628, w3531, IN41[19], w3629, w3630);
  FullAdder U923 (w3630, w3533, IN42[19], w3631, w3632);
  FullAdder U924 (w3632, w3535, IN43[19], w3633, w3634);
  FullAdder U925 (w3634, w3537, IN44[19], w3635, w3636);
  FullAdder U926 (w3636, w3539, IN45[19], w3637, w3638);
  FullAdder U927 (w3638, w3541, IN46[19], w3639, w3640);
  FullAdder U928 (w3640, w3543, IN47[19], w3641, w3642);
  FullAdder U929 (w3642, w3545, IN48[19], w3643, w3644);
  FullAdder U930 (w3644, w3547, IN49[19], w3645, w3646);
  FullAdder U931 (w3646, w3549, IN50[19], w3647, w3648);
  FullAdder U932 (w3648, w3551, IN51[17], w3649, w3650);
  FullAdder U933 (w3650, w3553, IN52[16], w3651, w3652);
  FullAdder U934 (w3652, w3555, IN53[15], w3653, w3654);
  FullAdder U935 (w3654, w3557, IN54[14], w3655, w3656);
  FullAdder U936 (w3656, w3559, IN55[13], w3657, w3658);
  FullAdder U937 (w3658, w3561, IN56[12], w3659, w3660);
  FullAdder U938 (w3660, w3563, IN57[11], w3661, w3662);
  FullAdder U939 (w3662, w3565, IN58[10], w3663, w3664);
  FullAdder U940 (w3664, w3567, IN59[9], w3665, w3666);
  FullAdder U941 (w3666, w3569, IN60[8], w3667, w3668);
  FullAdder U942 (w3668, w3571, IN61[7], w3669, w3670);
  FullAdder U943 (w3670, w3573, IN62[6], w3671, w3672);
  FullAdder U944 (w3672, w3575, IN63[5], w3673, w3674);
  FullAdder U945 (w3674, w3577, IN64[4], w3675, w3676);
  FullAdder U946 (w3676, w3579, IN65[3], w3677, w3678);
  FullAdder U947 (w3678, w3581, IN66[2], w3679, w3680);
  FullAdder U948 (w3680, w3583, IN67[1], w3681, w3682);
  FullAdder U949 (w3682, w3584, IN68[0], w3683, w3684);
  HalfAdder U950 (w3587, IN20[20], Out1[20], w3686);
  FullAdder U951 (w3686, w3589, IN21[20], w3687, w3688);
  FullAdder U952 (w3688, w3591, IN22[20], w3689, w3690);
  FullAdder U953 (w3690, w3593, IN23[20], w3691, w3692);
  FullAdder U954 (w3692, w3595, IN24[20], w3693, w3694);
  FullAdder U955 (w3694, w3597, IN25[20], w3695, w3696);
  FullAdder U956 (w3696, w3599, IN26[20], w3697, w3698);
  FullAdder U957 (w3698, w3601, IN27[20], w3699, w3700);
  FullAdder U958 (w3700, w3603, IN28[20], w3701, w3702);
  FullAdder U959 (w3702, w3605, IN29[20], w3703, w3704);
  FullAdder U960 (w3704, w3607, IN30[20], w3705, w3706);
  FullAdder U961 (w3706, w3609, IN31[20], w3707, w3708);
  FullAdder U962 (w3708, w3611, IN32[20], w3709, w3710);
  FullAdder U963 (w3710, w3613, IN33[20], w3711, w3712);
  FullAdder U964 (w3712, w3615, IN34[20], w3713, w3714);
  FullAdder U965 (w3714, w3617, IN35[20], w3715, w3716);
  FullAdder U966 (w3716, w3619, IN36[20], w3717, w3718);
  FullAdder U967 (w3718, w3621, IN37[20], w3719, w3720);
  FullAdder U968 (w3720, w3623, IN38[20], w3721, w3722);
  FullAdder U969 (w3722, w3625, IN39[20], w3723, w3724);
  FullAdder U970 (w3724, w3627, IN40[20], w3725, w3726);
  FullAdder U971 (w3726, w3629, IN41[20], w3727, w3728);
  FullAdder U972 (w3728, w3631, IN42[20], w3729, w3730);
  FullAdder U973 (w3730, w3633, IN43[20], w3731, w3732);
  FullAdder U974 (w3732, w3635, IN44[20], w3733, w3734);
  FullAdder U975 (w3734, w3637, IN45[20], w3735, w3736);
  FullAdder U976 (w3736, w3639, IN46[20], w3737, w3738);
  FullAdder U977 (w3738, w3641, IN47[20], w3739, w3740);
  FullAdder U978 (w3740, w3643, IN48[20], w3741, w3742);
  FullAdder U979 (w3742, w3645, IN49[20], w3743, w3744);
  FullAdder U980 (w3744, w3647, IN50[20], w3745, w3746);
  FullAdder U981 (w3746, w3649, IN51[18], w3747, w3748);
  FullAdder U982 (w3748, w3651, IN52[17], w3749, w3750);
  FullAdder U983 (w3750, w3653, IN53[16], w3751, w3752);
  FullAdder U984 (w3752, w3655, IN54[15], w3753, w3754);
  FullAdder U985 (w3754, w3657, IN55[14], w3755, w3756);
  FullAdder U986 (w3756, w3659, IN56[13], w3757, w3758);
  FullAdder U987 (w3758, w3661, IN57[12], w3759, w3760);
  FullAdder U988 (w3760, w3663, IN58[11], w3761, w3762);
  FullAdder U989 (w3762, w3665, IN59[10], w3763, w3764);
  FullAdder U990 (w3764, w3667, IN60[9], w3765, w3766);
  FullAdder U991 (w3766, w3669, IN61[8], w3767, w3768);
  FullAdder U992 (w3768, w3671, IN62[7], w3769, w3770);
  FullAdder U993 (w3770, w3673, IN63[6], w3771, w3772);
  FullAdder U994 (w3772, w3675, IN64[5], w3773, w3774);
  FullAdder U995 (w3774, w3677, IN65[4], w3775, w3776);
  FullAdder U996 (w3776, w3679, IN66[3], w3777, w3778);
  FullAdder U997 (w3778, w3681, IN67[2], w3779, w3780);
  FullAdder U998 (w3780, w3683, IN68[1], w3781, w3782);
  FullAdder U999 (w3782, w3684, IN69[0], w3783, w3784);
  HalfAdder U1000 (w3687, IN21[21], Out1[21], w3786);
  FullAdder U1001 (w3786, w3689, IN22[21], w3787, w3788);
  FullAdder U1002 (w3788, w3691, IN23[21], w3789, w3790);
  FullAdder U1003 (w3790, w3693, IN24[21], w3791, w3792);
  FullAdder U1004 (w3792, w3695, IN25[21], w3793, w3794);
  FullAdder U1005 (w3794, w3697, IN26[21], w3795, w3796);
  FullAdder U1006 (w3796, w3699, IN27[21], w3797, w3798);
  FullAdder U1007 (w3798, w3701, IN28[21], w3799, w3800);
  FullAdder U1008 (w3800, w3703, IN29[21], w3801, w3802);
  FullAdder U1009 (w3802, w3705, IN30[21], w3803, w3804);
  FullAdder U1010 (w3804, w3707, IN31[21], w3805, w3806);
  FullAdder U1011 (w3806, w3709, IN32[21], w3807, w3808);
  FullAdder U1012 (w3808, w3711, IN33[21], w3809, w3810);
  FullAdder U1013 (w3810, w3713, IN34[21], w3811, w3812);
  FullAdder U1014 (w3812, w3715, IN35[21], w3813, w3814);
  FullAdder U1015 (w3814, w3717, IN36[21], w3815, w3816);
  FullAdder U1016 (w3816, w3719, IN37[21], w3817, w3818);
  FullAdder U1017 (w3818, w3721, IN38[21], w3819, w3820);
  FullAdder U1018 (w3820, w3723, IN39[21], w3821, w3822);
  FullAdder U1019 (w3822, w3725, IN40[21], w3823, w3824);
  FullAdder U1020 (w3824, w3727, IN41[21], w3825, w3826);
  FullAdder U1021 (w3826, w3729, IN42[21], w3827, w3828);
  FullAdder U1022 (w3828, w3731, IN43[21], w3829, w3830);
  FullAdder U1023 (w3830, w3733, IN44[21], w3831, w3832);
  FullAdder U1024 (w3832, w3735, IN45[21], w3833, w3834);
  FullAdder U1025 (w3834, w3737, IN46[21], w3835, w3836);
  FullAdder U1026 (w3836, w3739, IN47[21], w3837, w3838);
  FullAdder U1027 (w3838, w3741, IN48[21], w3839, w3840);
  FullAdder U1028 (w3840, w3743, IN49[21], w3841, w3842);
  FullAdder U1029 (w3842, w3745, IN50[21], w3843, w3844);
  FullAdder U1030 (w3844, w3747, IN51[19], w3845, w3846);
  FullAdder U1031 (w3846, w3749, IN52[18], w3847, w3848);
  FullAdder U1032 (w3848, w3751, IN53[17], w3849, w3850);
  FullAdder U1033 (w3850, w3753, IN54[16], w3851, w3852);
  FullAdder U1034 (w3852, w3755, IN55[15], w3853, w3854);
  FullAdder U1035 (w3854, w3757, IN56[14], w3855, w3856);
  FullAdder U1036 (w3856, w3759, IN57[13], w3857, w3858);
  FullAdder U1037 (w3858, w3761, IN58[12], w3859, w3860);
  FullAdder U1038 (w3860, w3763, IN59[11], w3861, w3862);
  FullAdder U1039 (w3862, w3765, IN60[10], w3863, w3864);
  FullAdder U1040 (w3864, w3767, IN61[9], w3865, w3866);
  FullAdder U1041 (w3866, w3769, IN62[8], w3867, w3868);
  FullAdder U1042 (w3868, w3771, IN63[7], w3869, w3870);
  FullAdder U1043 (w3870, w3773, IN64[6], w3871, w3872);
  FullAdder U1044 (w3872, w3775, IN65[5], w3873, w3874);
  FullAdder U1045 (w3874, w3777, IN66[4], w3875, w3876);
  FullAdder U1046 (w3876, w3779, IN67[3], w3877, w3878);
  FullAdder U1047 (w3878, w3781, IN68[2], w3879, w3880);
  FullAdder U1048 (w3880, w3783, IN69[1], w3881, w3882);
  FullAdder U1049 (w3882, w3784, IN70[0], w3883, w3884);
  HalfAdder U1050 (w3787, IN22[22], Out1[22], w3886);
  FullAdder U1051 (w3886, w3789, IN23[22], w3887, w3888);
  FullAdder U1052 (w3888, w3791, IN24[22], w3889, w3890);
  FullAdder U1053 (w3890, w3793, IN25[22], w3891, w3892);
  FullAdder U1054 (w3892, w3795, IN26[22], w3893, w3894);
  FullAdder U1055 (w3894, w3797, IN27[22], w3895, w3896);
  FullAdder U1056 (w3896, w3799, IN28[22], w3897, w3898);
  FullAdder U1057 (w3898, w3801, IN29[22], w3899, w3900);
  FullAdder U1058 (w3900, w3803, IN30[22], w3901, w3902);
  FullAdder U1059 (w3902, w3805, IN31[22], w3903, w3904);
  FullAdder U1060 (w3904, w3807, IN32[22], w3905, w3906);
  FullAdder U1061 (w3906, w3809, IN33[22], w3907, w3908);
  FullAdder U1062 (w3908, w3811, IN34[22], w3909, w3910);
  FullAdder U1063 (w3910, w3813, IN35[22], w3911, w3912);
  FullAdder U1064 (w3912, w3815, IN36[22], w3913, w3914);
  FullAdder U1065 (w3914, w3817, IN37[22], w3915, w3916);
  FullAdder U1066 (w3916, w3819, IN38[22], w3917, w3918);
  FullAdder U1067 (w3918, w3821, IN39[22], w3919, w3920);
  FullAdder U1068 (w3920, w3823, IN40[22], w3921, w3922);
  FullAdder U1069 (w3922, w3825, IN41[22], w3923, w3924);
  FullAdder U1070 (w3924, w3827, IN42[22], w3925, w3926);
  FullAdder U1071 (w3926, w3829, IN43[22], w3927, w3928);
  FullAdder U1072 (w3928, w3831, IN44[22], w3929, w3930);
  FullAdder U1073 (w3930, w3833, IN45[22], w3931, w3932);
  FullAdder U1074 (w3932, w3835, IN46[22], w3933, w3934);
  FullAdder U1075 (w3934, w3837, IN47[22], w3935, w3936);
  FullAdder U1076 (w3936, w3839, IN48[22], w3937, w3938);
  FullAdder U1077 (w3938, w3841, IN49[22], w3939, w3940);
  FullAdder U1078 (w3940, w3843, IN50[22], w3941, w3942);
  FullAdder U1079 (w3942, w3845, IN51[20], w3943, w3944);
  FullAdder U1080 (w3944, w3847, IN52[19], w3945, w3946);
  FullAdder U1081 (w3946, w3849, IN53[18], w3947, w3948);
  FullAdder U1082 (w3948, w3851, IN54[17], w3949, w3950);
  FullAdder U1083 (w3950, w3853, IN55[16], w3951, w3952);
  FullAdder U1084 (w3952, w3855, IN56[15], w3953, w3954);
  FullAdder U1085 (w3954, w3857, IN57[14], w3955, w3956);
  FullAdder U1086 (w3956, w3859, IN58[13], w3957, w3958);
  FullAdder U1087 (w3958, w3861, IN59[12], w3959, w3960);
  FullAdder U1088 (w3960, w3863, IN60[11], w3961, w3962);
  FullAdder U1089 (w3962, w3865, IN61[10], w3963, w3964);
  FullAdder U1090 (w3964, w3867, IN62[9], w3965, w3966);
  FullAdder U1091 (w3966, w3869, IN63[8], w3967, w3968);
  FullAdder U1092 (w3968, w3871, IN64[7], w3969, w3970);
  FullAdder U1093 (w3970, w3873, IN65[6], w3971, w3972);
  FullAdder U1094 (w3972, w3875, IN66[5], w3973, w3974);
  FullAdder U1095 (w3974, w3877, IN67[4], w3975, w3976);
  FullAdder U1096 (w3976, w3879, IN68[3], w3977, w3978);
  FullAdder U1097 (w3978, w3881, IN69[2], w3979, w3980);
  FullAdder U1098 (w3980, w3883, IN70[1], w3981, w3982);
  FullAdder U1099 (w3982, w3884, IN71[0], w3983, w3984);
  HalfAdder U1100 (w3887, IN23[23], Out1[23], w3986);
  FullAdder U1101 (w3986, w3889, IN24[23], w3987, w3988);
  FullAdder U1102 (w3988, w3891, IN25[23], w3989, w3990);
  FullAdder U1103 (w3990, w3893, IN26[23], w3991, w3992);
  FullAdder U1104 (w3992, w3895, IN27[23], w3993, w3994);
  FullAdder U1105 (w3994, w3897, IN28[23], w3995, w3996);
  FullAdder U1106 (w3996, w3899, IN29[23], w3997, w3998);
  FullAdder U1107 (w3998, w3901, IN30[23], w3999, w4000);
  FullAdder U1108 (w4000, w3903, IN31[23], w4001, w4002);
  FullAdder U1109 (w4002, w3905, IN32[23], w4003, w4004);
  FullAdder U1110 (w4004, w3907, IN33[23], w4005, w4006);
  FullAdder U1111 (w4006, w3909, IN34[23], w4007, w4008);
  FullAdder U1112 (w4008, w3911, IN35[23], w4009, w4010);
  FullAdder U1113 (w4010, w3913, IN36[23], w4011, w4012);
  FullAdder U1114 (w4012, w3915, IN37[23], w4013, w4014);
  FullAdder U1115 (w4014, w3917, IN38[23], w4015, w4016);
  FullAdder U1116 (w4016, w3919, IN39[23], w4017, w4018);
  FullAdder U1117 (w4018, w3921, IN40[23], w4019, w4020);
  FullAdder U1118 (w4020, w3923, IN41[23], w4021, w4022);
  FullAdder U1119 (w4022, w3925, IN42[23], w4023, w4024);
  FullAdder U1120 (w4024, w3927, IN43[23], w4025, w4026);
  FullAdder U1121 (w4026, w3929, IN44[23], w4027, w4028);
  FullAdder U1122 (w4028, w3931, IN45[23], w4029, w4030);
  FullAdder U1123 (w4030, w3933, IN46[23], w4031, w4032);
  FullAdder U1124 (w4032, w3935, IN47[23], w4033, w4034);
  FullAdder U1125 (w4034, w3937, IN48[23], w4035, w4036);
  FullAdder U1126 (w4036, w3939, IN49[23], w4037, w4038);
  FullAdder U1127 (w4038, w3941, IN50[23], w4039, w4040);
  FullAdder U1128 (w4040, w3943, IN51[21], w4041, w4042);
  FullAdder U1129 (w4042, w3945, IN52[20], w4043, w4044);
  FullAdder U1130 (w4044, w3947, IN53[19], w4045, w4046);
  FullAdder U1131 (w4046, w3949, IN54[18], w4047, w4048);
  FullAdder U1132 (w4048, w3951, IN55[17], w4049, w4050);
  FullAdder U1133 (w4050, w3953, IN56[16], w4051, w4052);
  FullAdder U1134 (w4052, w3955, IN57[15], w4053, w4054);
  FullAdder U1135 (w4054, w3957, IN58[14], w4055, w4056);
  FullAdder U1136 (w4056, w3959, IN59[13], w4057, w4058);
  FullAdder U1137 (w4058, w3961, IN60[12], w4059, w4060);
  FullAdder U1138 (w4060, w3963, IN61[11], w4061, w4062);
  FullAdder U1139 (w4062, w3965, IN62[10], w4063, w4064);
  FullAdder U1140 (w4064, w3967, IN63[9], w4065, w4066);
  FullAdder U1141 (w4066, w3969, IN64[8], w4067, w4068);
  FullAdder U1142 (w4068, w3971, IN65[7], w4069, w4070);
  FullAdder U1143 (w4070, w3973, IN66[6], w4071, w4072);
  FullAdder U1144 (w4072, w3975, IN67[5], w4073, w4074);
  FullAdder U1145 (w4074, w3977, IN68[4], w4075, w4076);
  FullAdder U1146 (w4076, w3979, IN69[3], w4077, w4078);
  FullAdder U1147 (w4078, w3981, IN70[2], w4079, w4080);
  FullAdder U1148 (w4080, w3983, IN71[1], w4081, w4082);
  FullAdder U1149 (w4082, w3984, IN72[0], w4083, w4084);
  HalfAdder U1150 (w3987, IN24[24], Out1[24], w4086);
  FullAdder U1151 (w4086, w3989, IN25[24], w4087, w4088);
  FullAdder U1152 (w4088, w3991, IN26[24], w4089, w4090);
  FullAdder U1153 (w4090, w3993, IN27[24], w4091, w4092);
  FullAdder U1154 (w4092, w3995, IN28[24], w4093, w4094);
  FullAdder U1155 (w4094, w3997, IN29[24], w4095, w4096);
  FullAdder U1156 (w4096, w3999, IN30[24], w4097, w4098);
  FullAdder U1157 (w4098, w4001, IN31[24], w4099, w4100);
  FullAdder U1158 (w4100, w4003, IN32[24], w4101, w4102);
  FullAdder U1159 (w4102, w4005, IN33[24], w4103, w4104);
  FullAdder U1160 (w4104, w4007, IN34[24], w4105, w4106);
  FullAdder U1161 (w4106, w4009, IN35[24], w4107, w4108);
  FullAdder U1162 (w4108, w4011, IN36[24], w4109, w4110);
  FullAdder U1163 (w4110, w4013, IN37[24], w4111, w4112);
  FullAdder U1164 (w4112, w4015, IN38[24], w4113, w4114);
  FullAdder U1165 (w4114, w4017, IN39[24], w4115, w4116);
  FullAdder U1166 (w4116, w4019, IN40[24], w4117, w4118);
  FullAdder U1167 (w4118, w4021, IN41[24], w4119, w4120);
  FullAdder U1168 (w4120, w4023, IN42[24], w4121, w4122);
  FullAdder U1169 (w4122, w4025, IN43[24], w4123, w4124);
  FullAdder U1170 (w4124, w4027, IN44[24], w4125, w4126);
  FullAdder U1171 (w4126, w4029, IN45[24], w4127, w4128);
  FullAdder U1172 (w4128, w4031, IN46[24], w4129, w4130);
  FullAdder U1173 (w4130, w4033, IN47[24], w4131, w4132);
  FullAdder U1174 (w4132, w4035, IN48[24], w4133, w4134);
  FullAdder U1175 (w4134, w4037, IN49[24], w4135, w4136);
  FullAdder U1176 (w4136, w4039, IN50[24], w4137, w4138);
  FullAdder U1177 (w4138, w4041, IN51[22], w4139, w4140);
  FullAdder U1178 (w4140, w4043, IN52[21], w4141, w4142);
  FullAdder U1179 (w4142, w4045, IN53[20], w4143, w4144);
  FullAdder U1180 (w4144, w4047, IN54[19], w4145, w4146);
  FullAdder U1181 (w4146, w4049, IN55[18], w4147, w4148);
  FullAdder U1182 (w4148, w4051, IN56[17], w4149, w4150);
  FullAdder U1183 (w4150, w4053, IN57[16], w4151, w4152);
  FullAdder U1184 (w4152, w4055, IN58[15], w4153, w4154);
  FullAdder U1185 (w4154, w4057, IN59[14], w4155, w4156);
  FullAdder U1186 (w4156, w4059, IN60[13], w4157, w4158);
  FullAdder U1187 (w4158, w4061, IN61[12], w4159, w4160);
  FullAdder U1188 (w4160, w4063, IN62[11], w4161, w4162);
  FullAdder U1189 (w4162, w4065, IN63[10], w4163, w4164);
  FullAdder U1190 (w4164, w4067, IN64[9], w4165, w4166);
  FullAdder U1191 (w4166, w4069, IN65[8], w4167, w4168);
  FullAdder U1192 (w4168, w4071, IN66[7], w4169, w4170);
  FullAdder U1193 (w4170, w4073, IN67[6], w4171, w4172);
  FullAdder U1194 (w4172, w4075, IN68[5], w4173, w4174);
  FullAdder U1195 (w4174, w4077, IN69[4], w4175, w4176);
  FullAdder U1196 (w4176, w4079, IN70[3], w4177, w4178);
  FullAdder U1197 (w4178, w4081, IN71[2], w4179, w4180);
  FullAdder U1198 (w4180, w4083, IN72[1], w4181, w4182);
  FullAdder U1199 (w4182, w4084, IN73[0], w4183, w4184);
  HalfAdder U1200 (w4087, IN25[25], Out1[25], w4186);
  FullAdder U1201 (w4186, w4089, IN26[25], w4187, w4188);
  FullAdder U1202 (w4188, w4091, IN27[25], w4189, w4190);
  FullAdder U1203 (w4190, w4093, IN28[25], w4191, w4192);
  FullAdder U1204 (w4192, w4095, IN29[25], w4193, w4194);
  FullAdder U1205 (w4194, w4097, IN30[25], w4195, w4196);
  FullAdder U1206 (w4196, w4099, IN31[25], w4197, w4198);
  FullAdder U1207 (w4198, w4101, IN32[25], w4199, w4200);
  FullAdder U1208 (w4200, w4103, IN33[25], w4201, w4202);
  FullAdder U1209 (w4202, w4105, IN34[25], w4203, w4204);
  FullAdder U1210 (w4204, w4107, IN35[25], w4205, w4206);
  FullAdder U1211 (w4206, w4109, IN36[25], w4207, w4208);
  FullAdder U1212 (w4208, w4111, IN37[25], w4209, w4210);
  FullAdder U1213 (w4210, w4113, IN38[25], w4211, w4212);
  FullAdder U1214 (w4212, w4115, IN39[25], w4213, w4214);
  FullAdder U1215 (w4214, w4117, IN40[25], w4215, w4216);
  FullAdder U1216 (w4216, w4119, IN41[25], w4217, w4218);
  FullAdder U1217 (w4218, w4121, IN42[25], w4219, w4220);
  FullAdder U1218 (w4220, w4123, IN43[25], w4221, w4222);
  FullAdder U1219 (w4222, w4125, IN44[25], w4223, w4224);
  FullAdder U1220 (w4224, w4127, IN45[25], w4225, w4226);
  FullAdder U1221 (w4226, w4129, IN46[25], w4227, w4228);
  FullAdder U1222 (w4228, w4131, IN47[25], w4229, w4230);
  FullAdder U1223 (w4230, w4133, IN48[25], w4231, w4232);
  FullAdder U1224 (w4232, w4135, IN49[25], w4233, w4234);
  FullAdder U1225 (w4234, w4137, IN50[25], w4235, w4236);
  FullAdder U1226 (w4236, w4139, IN51[23], w4237, w4238);
  FullAdder U1227 (w4238, w4141, IN52[22], w4239, w4240);
  FullAdder U1228 (w4240, w4143, IN53[21], w4241, w4242);
  FullAdder U1229 (w4242, w4145, IN54[20], w4243, w4244);
  FullAdder U1230 (w4244, w4147, IN55[19], w4245, w4246);
  FullAdder U1231 (w4246, w4149, IN56[18], w4247, w4248);
  FullAdder U1232 (w4248, w4151, IN57[17], w4249, w4250);
  FullAdder U1233 (w4250, w4153, IN58[16], w4251, w4252);
  FullAdder U1234 (w4252, w4155, IN59[15], w4253, w4254);
  FullAdder U1235 (w4254, w4157, IN60[14], w4255, w4256);
  FullAdder U1236 (w4256, w4159, IN61[13], w4257, w4258);
  FullAdder U1237 (w4258, w4161, IN62[12], w4259, w4260);
  FullAdder U1238 (w4260, w4163, IN63[11], w4261, w4262);
  FullAdder U1239 (w4262, w4165, IN64[10], w4263, w4264);
  FullAdder U1240 (w4264, w4167, IN65[9], w4265, w4266);
  FullAdder U1241 (w4266, w4169, IN66[8], w4267, w4268);
  FullAdder U1242 (w4268, w4171, IN67[7], w4269, w4270);
  FullAdder U1243 (w4270, w4173, IN68[6], w4271, w4272);
  FullAdder U1244 (w4272, w4175, IN69[5], w4273, w4274);
  FullAdder U1245 (w4274, w4177, IN70[4], w4275, w4276);
  FullAdder U1246 (w4276, w4179, IN71[3], w4277, w4278);
  FullAdder U1247 (w4278, w4181, IN72[2], w4279, w4280);
  FullAdder U1248 (w4280, w4183, IN73[1], w4281, w4282);
  FullAdder U1249 (w4282, w4184, IN74[0], w4283, w4284);
  HalfAdder U1250 (w4187, IN26[26], Out1[26], w4286);
  FullAdder U1251 (w4286, w4189, IN27[26], w4287, w4288);
  FullAdder U1252 (w4288, w4191, IN28[26], w4289, w4290);
  FullAdder U1253 (w4290, w4193, IN29[26], w4291, w4292);
  FullAdder U1254 (w4292, w4195, IN30[26], w4293, w4294);
  FullAdder U1255 (w4294, w4197, IN31[26], w4295, w4296);
  FullAdder U1256 (w4296, w4199, IN32[26], w4297, w4298);
  FullAdder U1257 (w4298, w4201, IN33[26], w4299, w4300);
  FullAdder U1258 (w4300, w4203, IN34[26], w4301, w4302);
  FullAdder U1259 (w4302, w4205, IN35[26], w4303, w4304);
  FullAdder U1260 (w4304, w4207, IN36[26], w4305, w4306);
  FullAdder U1261 (w4306, w4209, IN37[26], w4307, w4308);
  FullAdder U1262 (w4308, w4211, IN38[26], w4309, w4310);
  FullAdder U1263 (w4310, w4213, IN39[26], w4311, w4312);
  FullAdder U1264 (w4312, w4215, IN40[26], w4313, w4314);
  FullAdder U1265 (w4314, w4217, IN41[26], w4315, w4316);
  FullAdder U1266 (w4316, w4219, IN42[26], w4317, w4318);
  FullAdder U1267 (w4318, w4221, IN43[26], w4319, w4320);
  FullAdder U1268 (w4320, w4223, IN44[26], w4321, w4322);
  FullAdder U1269 (w4322, w4225, IN45[26], w4323, w4324);
  FullAdder U1270 (w4324, w4227, IN46[26], w4325, w4326);
  FullAdder U1271 (w4326, w4229, IN47[26], w4327, w4328);
  FullAdder U1272 (w4328, w4231, IN48[26], w4329, w4330);
  FullAdder U1273 (w4330, w4233, IN49[26], w4331, w4332);
  FullAdder U1274 (w4332, w4235, IN50[26], w4333, w4334);
  FullAdder U1275 (w4334, w4237, IN51[24], w4335, w4336);
  FullAdder U1276 (w4336, w4239, IN52[23], w4337, w4338);
  FullAdder U1277 (w4338, w4241, IN53[22], w4339, w4340);
  FullAdder U1278 (w4340, w4243, IN54[21], w4341, w4342);
  FullAdder U1279 (w4342, w4245, IN55[20], w4343, w4344);
  FullAdder U1280 (w4344, w4247, IN56[19], w4345, w4346);
  FullAdder U1281 (w4346, w4249, IN57[18], w4347, w4348);
  FullAdder U1282 (w4348, w4251, IN58[17], w4349, w4350);
  FullAdder U1283 (w4350, w4253, IN59[16], w4351, w4352);
  FullAdder U1284 (w4352, w4255, IN60[15], w4353, w4354);
  FullAdder U1285 (w4354, w4257, IN61[14], w4355, w4356);
  FullAdder U1286 (w4356, w4259, IN62[13], w4357, w4358);
  FullAdder U1287 (w4358, w4261, IN63[12], w4359, w4360);
  FullAdder U1288 (w4360, w4263, IN64[11], w4361, w4362);
  FullAdder U1289 (w4362, w4265, IN65[10], w4363, w4364);
  FullAdder U1290 (w4364, w4267, IN66[9], w4365, w4366);
  FullAdder U1291 (w4366, w4269, IN67[8], w4367, w4368);
  FullAdder U1292 (w4368, w4271, IN68[7], w4369, w4370);
  FullAdder U1293 (w4370, w4273, IN69[6], w4371, w4372);
  FullAdder U1294 (w4372, w4275, IN70[5], w4373, w4374);
  FullAdder U1295 (w4374, w4277, IN71[4], w4375, w4376);
  FullAdder U1296 (w4376, w4279, IN72[3], w4377, w4378);
  FullAdder U1297 (w4378, w4281, IN73[2], w4379, w4380);
  FullAdder U1298 (w4380, w4283, IN74[1], w4381, w4382);
  FullAdder U1299 (w4382, w4284, IN75[0], w4383, w4384);
  HalfAdder U1300 (w4287, IN27[27], Out1[27], w4386);
  FullAdder U1301 (w4386, w4289, IN28[27], w4387, w4388);
  FullAdder U1302 (w4388, w4291, IN29[27], w4389, w4390);
  FullAdder U1303 (w4390, w4293, IN30[27], w4391, w4392);
  FullAdder U1304 (w4392, w4295, IN31[27], w4393, w4394);
  FullAdder U1305 (w4394, w4297, IN32[27], w4395, w4396);
  FullAdder U1306 (w4396, w4299, IN33[27], w4397, w4398);
  FullAdder U1307 (w4398, w4301, IN34[27], w4399, w4400);
  FullAdder U1308 (w4400, w4303, IN35[27], w4401, w4402);
  FullAdder U1309 (w4402, w4305, IN36[27], w4403, w4404);
  FullAdder U1310 (w4404, w4307, IN37[27], w4405, w4406);
  FullAdder U1311 (w4406, w4309, IN38[27], w4407, w4408);
  FullAdder U1312 (w4408, w4311, IN39[27], w4409, w4410);
  FullAdder U1313 (w4410, w4313, IN40[27], w4411, w4412);
  FullAdder U1314 (w4412, w4315, IN41[27], w4413, w4414);
  FullAdder U1315 (w4414, w4317, IN42[27], w4415, w4416);
  FullAdder U1316 (w4416, w4319, IN43[27], w4417, w4418);
  FullAdder U1317 (w4418, w4321, IN44[27], w4419, w4420);
  FullAdder U1318 (w4420, w4323, IN45[27], w4421, w4422);
  FullAdder U1319 (w4422, w4325, IN46[27], w4423, w4424);
  FullAdder U1320 (w4424, w4327, IN47[27], w4425, w4426);
  FullAdder U1321 (w4426, w4329, IN48[27], w4427, w4428);
  FullAdder U1322 (w4428, w4331, IN49[27], w4429, w4430);
  FullAdder U1323 (w4430, w4333, IN50[27], w4431, w4432);
  FullAdder U1324 (w4432, w4335, IN51[25], w4433, w4434);
  FullAdder U1325 (w4434, w4337, IN52[24], w4435, w4436);
  FullAdder U1326 (w4436, w4339, IN53[23], w4437, w4438);
  FullAdder U1327 (w4438, w4341, IN54[22], w4439, w4440);
  FullAdder U1328 (w4440, w4343, IN55[21], w4441, w4442);
  FullAdder U1329 (w4442, w4345, IN56[20], w4443, w4444);
  FullAdder U1330 (w4444, w4347, IN57[19], w4445, w4446);
  FullAdder U1331 (w4446, w4349, IN58[18], w4447, w4448);
  FullAdder U1332 (w4448, w4351, IN59[17], w4449, w4450);
  FullAdder U1333 (w4450, w4353, IN60[16], w4451, w4452);
  FullAdder U1334 (w4452, w4355, IN61[15], w4453, w4454);
  FullAdder U1335 (w4454, w4357, IN62[14], w4455, w4456);
  FullAdder U1336 (w4456, w4359, IN63[13], w4457, w4458);
  FullAdder U1337 (w4458, w4361, IN64[12], w4459, w4460);
  FullAdder U1338 (w4460, w4363, IN65[11], w4461, w4462);
  FullAdder U1339 (w4462, w4365, IN66[10], w4463, w4464);
  FullAdder U1340 (w4464, w4367, IN67[9], w4465, w4466);
  FullAdder U1341 (w4466, w4369, IN68[8], w4467, w4468);
  FullAdder U1342 (w4468, w4371, IN69[7], w4469, w4470);
  FullAdder U1343 (w4470, w4373, IN70[6], w4471, w4472);
  FullAdder U1344 (w4472, w4375, IN71[5], w4473, w4474);
  FullAdder U1345 (w4474, w4377, IN72[4], w4475, w4476);
  FullAdder U1346 (w4476, w4379, IN73[3], w4477, w4478);
  FullAdder U1347 (w4478, w4381, IN74[2], w4479, w4480);
  FullAdder U1348 (w4480, w4383, IN75[1], w4481, w4482);
  FullAdder U1349 (w4482, w4384, IN76[0], w4483, w4484);
  HalfAdder U1350 (w4387, IN28[28], Out1[28], w4486);
  FullAdder U1351 (w4486, w4389, IN29[28], w4487, w4488);
  FullAdder U1352 (w4488, w4391, IN30[28], w4489, w4490);
  FullAdder U1353 (w4490, w4393, IN31[28], w4491, w4492);
  FullAdder U1354 (w4492, w4395, IN32[28], w4493, w4494);
  FullAdder U1355 (w4494, w4397, IN33[28], w4495, w4496);
  FullAdder U1356 (w4496, w4399, IN34[28], w4497, w4498);
  FullAdder U1357 (w4498, w4401, IN35[28], w4499, w4500);
  FullAdder U1358 (w4500, w4403, IN36[28], w4501, w4502);
  FullAdder U1359 (w4502, w4405, IN37[28], w4503, w4504);
  FullAdder U1360 (w4504, w4407, IN38[28], w4505, w4506);
  FullAdder U1361 (w4506, w4409, IN39[28], w4507, w4508);
  FullAdder U1362 (w4508, w4411, IN40[28], w4509, w4510);
  FullAdder U1363 (w4510, w4413, IN41[28], w4511, w4512);
  FullAdder U1364 (w4512, w4415, IN42[28], w4513, w4514);
  FullAdder U1365 (w4514, w4417, IN43[28], w4515, w4516);
  FullAdder U1366 (w4516, w4419, IN44[28], w4517, w4518);
  FullAdder U1367 (w4518, w4421, IN45[28], w4519, w4520);
  FullAdder U1368 (w4520, w4423, IN46[28], w4521, w4522);
  FullAdder U1369 (w4522, w4425, IN47[28], w4523, w4524);
  FullAdder U1370 (w4524, w4427, IN48[28], w4525, w4526);
  FullAdder U1371 (w4526, w4429, IN49[28], w4527, w4528);
  FullAdder U1372 (w4528, w4431, IN50[28], w4529, w4530);
  FullAdder U1373 (w4530, w4433, IN51[26], w4531, w4532);
  FullAdder U1374 (w4532, w4435, IN52[25], w4533, w4534);
  FullAdder U1375 (w4534, w4437, IN53[24], w4535, w4536);
  FullAdder U1376 (w4536, w4439, IN54[23], w4537, w4538);
  FullAdder U1377 (w4538, w4441, IN55[22], w4539, w4540);
  FullAdder U1378 (w4540, w4443, IN56[21], w4541, w4542);
  FullAdder U1379 (w4542, w4445, IN57[20], w4543, w4544);
  FullAdder U1380 (w4544, w4447, IN58[19], w4545, w4546);
  FullAdder U1381 (w4546, w4449, IN59[18], w4547, w4548);
  FullAdder U1382 (w4548, w4451, IN60[17], w4549, w4550);
  FullAdder U1383 (w4550, w4453, IN61[16], w4551, w4552);
  FullAdder U1384 (w4552, w4455, IN62[15], w4553, w4554);
  FullAdder U1385 (w4554, w4457, IN63[14], w4555, w4556);
  FullAdder U1386 (w4556, w4459, IN64[13], w4557, w4558);
  FullAdder U1387 (w4558, w4461, IN65[12], w4559, w4560);
  FullAdder U1388 (w4560, w4463, IN66[11], w4561, w4562);
  FullAdder U1389 (w4562, w4465, IN67[10], w4563, w4564);
  FullAdder U1390 (w4564, w4467, IN68[9], w4565, w4566);
  FullAdder U1391 (w4566, w4469, IN69[8], w4567, w4568);
  FullAdder U1392 (w4568, w4471, IN70[7], w4569, w4570);
  FullAdder U1393 (w4570, w4473, IN71[6], w4571, w4572);
  FullAdder U1394 (w4572, w4475, IN72[5], w4573, w4574);
  FullAdder U1395 (w4574, w4477, IN73[4], w4575, w4576);
  FullAdder U1396 (w4576, w4479, IN74[3], w4577, w4578);
  FullAdder U1397 (w4578, w4481, IN75[2], w4579, w4580);
  FullAdder U1398 (w4580, w4483, IN76[1], w4581, w4582);
  FullAdder U1399 (w4582, w4484, IN77[0], w4583, w4584);
  HalfAdder U1400 (w4487, IN29[29], Out1[29], w4586);
  FullAdder U1401 (w4586, w4489, IN30[29], w4587, w4588);
  FullAdder U1402 (w4588, w4491, IN31[29], w4589, w4590);
  FullAdder U1403 (w4590, w4493, IN32[29], w4591, w4592);
  FullAdder U1404 (w4592, w4495, IN33[29], w4593, w4594);
  FullAdder U1405 (w4594, w4497, IN34[29], w4595, w4596);
  FullAdder U1406 (w4596, w4499, IN35[29], w4597, w4598);
  FullAdder U1407 (w4598, w4501, IN36[29], w4599, w4600);
  FullAdder U1408 (w4600, w4503, IN37[29], w4601, w4602);
  FullAdder U1409 (w4602, w4505, IN38[29], w4603, w4604);
  FullAdder U1410 (w4604, w4507, IN39[29], w4605, w4606);
  FullAdder U1411 (w4606, w4509, IN40[29], w4607, w4608);
  FullAdder U1412 (w4608, w4511, IN41[29], w4609, w4610);
  FullAdder U1413 (w4610, w4513, IN42[29], w4611, w4612);
  FullAdder U1414 (w4612, w4515, IN43[29], w4613, w4614);
  FullAdder U1415 (w4614, w4517, IN44[29], w4615, w4616);
  FullAdder U1416 (w4616, w4519, IN45[29], w4617, w4618);
  FullAdder U1417 (w4618, w4521, IN46[29], w4619, w4620);
  FullAdder U1418 (w4620, w4523, IN47[29], w4621, w4622);
  FullAdder U1419 (w4622, w4525, IN48[29], w4623, w4624);
  FullAdder U1420 (w4624, w4527, IN49[29], w4625, w4626);
  FullAdder U1421 (w4626, w4529, IN50[29], w4627, w4628);
  FullAdder U1422 (w4628, w4531, IN51[27], w4629, w4630);
  FullAdder U1423 (w4630, w4533, IN52[26], w4631, w4632);
  FullAdder U1424 (w4632, w4535, IN53[25], w4633, w4634);
  FullAdder U1425 (w4634, w4537, IN54[24], w4635, w4636);
  FullAdder U1426 (w4636, w4539, IN55[23], w4637, w4638);
  FullAdder U1427 (w4638, w4541, IN56[22], w4639, w4640);
  FullAdder U1428 (w4640, w4543, IN57[21], w4641, w4642);
  FullAdder U1429 (w4642, w4545, IN58[20], w4643, w4644);
  FullAdder U1430 (w4644, w4547, IN59[19], w4645, w4646);
  FullAdder U1431 (w4646, w4549, IN60[18], w4647, w4648);
  FullAdder U1432 (w4648, w4551, IN61[17], w4649, w4650);
  FullAdder U1433 (w4650, w4553, IN62[16], w4651, w4652);
  FullAdder U1434 (w4652, w4555, IN63[15], w4653, w4654);
  FullAdder U1435 (w4654, w4557, IN64[14], w4655, w4656);
  FullAdder U1436 (w4656, w4559, IN65[13], w4657, w4658);
  FullAdder U1437 (w4658, w4561, IN66[12], w4659, w4660);
  FullAdder U1438 (w4660, w4563, IN67[11], w4661, w4662);
  FullAdder U1439 (w4662, w4565, IN68[10], w4663, w4664);
  FullAdder U1440 (w4664, w4567, IN69[9], w4665, w4666);
  FullAdder U1441 (w4666, w4569, IN70[8], w4667, w4668);
  FullAdder U1442 (w4668, w4571, IN71[7], w4669, w4670);
  FullAdder U1443 (w4670, w4573, IN72[6], w4671, w4672);
  FullAdder U1444 (w4672, w4575, IN73[5], w4673, w4674);
  FullAdder U1445 (w4674, w4577, IN74[4], w4675, w4676);
  FullAdder U1446 (w4676, w4579, IN75[3], w4677, w4678);
  FullAdder U1447 (w4678, w4581, IN76[2], w4679, w4680);
  FullAdder U1448 (w4680, w4583, IN77[1], w4681, w4682);
  FullAdder U1449 (w4682, w4584, IN78[0], w4683, w4684);
  HalfAdder U1450 (w4587, IN30[30], Out1[30], w4686);
  FullAdder U1451 (w4686, w4589, IN31[30], w4687, w4688);
  FullAdder U1452 (w4688, w4591, IN32[30], w4689, w4690);
  FullAdder U1453 (w4690, w4593, IN33[30], w4691, w4692);
  FullAdder U1454 (w4692, w4595, IN34[30], w4693, w4694);
  FullAdder U1455 (w4694, w4597, IN35[30], w4695, w4696);
  FullAdder U1456 (w4696, w4599, IN36[30], w4697, w4698);
  FullAdder U1457 (w4698, w4601, IN37[30], w4699, w4700);
  FullAdder U1458 (w4700, w4603, IN38[30], w4701, w4702);
  FullAdder U1459 (w4702, w4605, IN39[30], w4703, w4704);
  FullAdder U1460 (w4704, w4607, IN40[30], w4705, w4706);
  FullAdder U1461 (w4706, w4609, IN41[30], w4707, w4708);
  FullAdder U1462 (w4708, w4611, IN42[30], w4709, w4710);
  FullAdder U1463 (w4710, w4613, IN43[30], w4711, w4712);
  FullAdder U1464 (w4712, w4615, IN44[30], w4713, w4714);
  FullAdder U1465 (w4714, w4617, IN45[30], w4715, w4716);
  FullAdder U1466 (w4716, w4619, IN46[30], w4717, w4718);
  FullAdder U1467 (w4718, w4621, IN47[30], w4719, w4720);
  FullAdder U1468 (w4720, w4623, IN48[30], w4721, w4722);
  FullAdder U1469 (w4722, w4625, IN49[30], w4723, w4724);
  FullAdder U1470 (w4724, w4627, IN50[30], w4725, w4726);
  FullAdder U1471 (w4726, w4629, IN51[28], w4727, w4728);
  FullAdder U1472 (w4728, w4631, IN52[27], w4729, w4730);
  FullAdder U1473 (w4730, w4633, IN53[26], w4731, w4732);
  FullAdder U1474 (w4732, w4635, IN54[25], w4733, w4734);
  FullAdder U1475 (w4734, w4637, IN55[24], w4735, w4736);
  FullAdder U1476 (w4736, w4639, IN56[23], w4737, w4738);
  FullAdder U1477 (w4738, w4641, IN57[22], w4739, w4740);
  FullAdder U1478 (w4740, w4643, IN58[21], w4741, w4742);
  FullAdder U1479 (w4742, w4645, IN59[20], w4743, w4744);
  FullAdder U1480 (w4744, w4647, IN60[19], w4745, w4746);
  FullAdder U1481 (w4746, w4649, IN61[18], w4747, w4748);
  FullAdder U1482 (w4748, w4651, IN62[17], w4749, w4750);
  FullAdder U1483 (w4750, w4653, IN63[16], w4751, w4752);
  FullAdder U1484 (w4752, w4655, IN64[15], w4753, w4754);
  FullAdder U1485 (w4754, w4657, IN65[14], w4755, w4756);
  FullAdder U1486 (w4756, w4659, IN66[13], w4757, w4758);
  FullAdder U1487 (w4758, w4661, IN67[12], w4759, w4760);
  FullAdder U1488 (w4760, w4663, IN68[11], w4761, w4762);
  FullAdder U1489 (w4762, w4665, IN69[10], w4763, w4764);
  FullAdder U1490 (w4764, w4667, IN70[9], w4765, w4766);
  FullAdder U1491 (w4766, w4669, IN71[8], w4767, w4768);
  FullAdder U1492 (w4768, w4671, IN72[7], w4769, w4770);
  FullAdder U1493 (w4770, w4673, IN73[6], w4771, w4772);
  FullAdder U1494 (w4772, w4675, IN74[5], w4773, w4774);
  FullAdder U1495 (w4774, w4677, IN75[4], w4775, w4776);
  FullAdder U1496 (w4776, w4679, IN76[3], w4777, w4778);
  FullAdder U1497 (w4778, w4681, IN77[2], w4779, w4780);
  FullAdder U1498 (w4780, w4683, IN78[1], w4781, w4782);
  FullAdder U1499 (w4782, w4684, IN79[0], w4783, w4784);
  HalfAdder U1500 (w4687, IN31[31], Out1[31], w4786);
  FullAdder U1501 (w4786, w4689, IN32[31], w4787, w4788);
  FullAdder U1502 (w4788, w4691, IN33[31], w4789, w4790);
  FullAdder U1503 (w4790, w4693, IN34[31], w4791, w4792);
  FullAdder U1504 (w4792, w4695, IN35[31], w4793, w4794);
  FullAdder U1505 (w4794, w4697, IN36[31], w4795, w4796);
  FullAdder U1506 (w4796, w4699, IN37[31], w4797, w4798);
  FullAdder U1507 (w4798, w4701, IN38[31], w4799, w4800);
  FullAdder U1508 (w4800, w4703, IN39[31], w4801, w4802);
  FullAdder U1509 (w4802, w4705, IN40[31], w4803, w4804);
  FullAdder U1510 (w4804, w4707, IN41[31], w4805, w4806);
  FullAdder U1511 (w4806, w4709, IN42[31], w4807, w4808);
  FullAdder U1512 (w4808, w4711, IN43[31], w4809, w4810);
  FullAdder U1513 (w4810, w4713, IN44[31], w4811, w4812);
  FullAdder U1514 (w4812, w4715, IN45[31], w4813, w4814);
  FullAdder U1515 (w4814, w4717, IN46[31], w4815, w4816);
  FullAdder U1516 (w4816, w4719, IN47[31], w4817, w4818);
  FullAdder U1517 (w4818, w4721, IN48[31], w4819, w4820);
  FullAdder U1518 (w4820, w4723, IN49[31], w4821, w4822);
  FullAdder U1519 (w4822, w4725, IN50[31], w4823, w4824);
  FullAdder U1520 (w4824, w4727, IN51[29], w4825, w4826);
  FullAdder U1521 (w4826, w4729, IN52[28], w4827, w4828);
  FullAdder U1522 (w4828, w4731, IN53[27], w4829, w4830);
  FullAdder U1523 (w4830, w4733, IN54[26], w4831, w4832);
  FullAdder U1524 (w4832, w4735, IN55[25], w4833, w4834);
  FullAdder U1525 (w4834, w4737, IN56[24], w4835, w4836);
  FullAdder U1526 (w4836, w4739, IN57[23], w4837, w4838);
  FullAdder U1527 (w4838, w4741, IN58[22], w4839, w4840);
  FullAdder U1528 (w4840, w4743, IN59[21], w4841, w4842);
  FullAdder U1529 (w4842, w4745, IN60[20], w4843, w4844);
  FullAdder U1530 (w4844, w4747, IN61[19], w4845, w4846);
  FullAdder U1531 (w4846, w4749, IN62[18], w4847, w4848);
  FullAdder U1532 (w4848, w4751, IN63[17], w4849, w4850);
  FullAdder U1533 (w4850, w4753, IN64[16], w4851, w4852);
  FullAdder U1534 (w4852, w4755, IN65[15], w4853, w4854);
  FullAdder U1535 (w4854, w4757, IN66[14], w4855, w4856);
  FullAdder U1536 (w4856, w4759, IN67[13], w4857, w4858);
  FullAdder U1537 (w4858, w4761, IN68[12], w4859, w4860);
  FullAdder U1538 (w4860, w4763, IN69[11], w4861, w4862);
  FullAdder U1539 (w4862, w4765, IN70[10], w4863, w4864);
  FullAdder U1540 (w4864, w4767, IN71[9], w4865, w4866);
  FullAdder U1541 (w4866, w4769, IN72[8], w4867, w4868);
  FullAdder U1542 (w4868, w4771, IN73[7], w4869, w4870);
  FullAdder U1543 (w4870, w4773, IN74[6], w4871, w4872);
  FullAdder U1544 (w4872, w4775, IN75[5], w4873, w4874);
  FullAdder U1545 (w4874, w4777, IN76[4], w4875, w4876);
  FullAdder U1546 (w4876, w4779, IN77[3], w4877, w4878);
  FullAdder U1547 (w4878, w4781, IN78[2], w4879, w4880);
  FullAdder U1548 (w4880, w4783, IN79[1], w4881, w4882);
  FullAdder U1549 (w4882, w4784, IN80[0], w4883, w4884);
  HalfAdder U1550 (w4787, IN32[32], Out1[32], w4886);
  FullAdder U1551 (w4886, w4789, IN33[32], w4887, w4888);
  FullAdder U1552 (w4888, w4791, IN34[32], w4889, w4890);
  FullAdder U1553 (w4890, w4793, IN35[32], w4891, w4892);
  FullAdder U1554 (w4892, w4795, IN36[32], w4893, w4894);
  FullAdder U1555 (w4894, w4797, IN37[32], w4895, w4896);
  FullAdder U1556 (w4896, w4799, IN38[32], w4897, w4898);
  FullAdder U1557 (w4898, w4801, IN39[32], w4899, w4900);
  FullAdder U1558 (w4900, w4803, IN40[32], w4901, w4902);
  FullAdder U1559 (w4902, w4805, IN41[32], w4903, w4904);
  FullAdder U1560 (w4904, w4807, IN42[32], w4905, w4906);
  FullAdder U1561 (w4906, w4809, IN43[32], w4907, w4908);
  FullAdder U1562 (w4908, w4811, IN44[32], w4909, w4910);
  FullAdder U1563 (w4910, w4813, IN45[32], w4911, w4912);
  FullAdder U1564 (w4912, w4815, IN46[32], w4913, w4914);
  FullAdder U1565 (w4914, w4817, IN47[32], w4915, w4916);
  FullAdder U1566 (w4916, w4819, IN48[32], w4917, w4918);
  FullAdder U1567 (w4918, w4821, IN49[32], w4919, w4920);
  FullAdder U1568 (w4920, w4823, IN50[32], w4921, w4922);
  FullAdder U1569 (w4922, w4825, IN51[30], w4923, w4924);
  FullAdder U1570 (w4924, w4827, IN52[29], w4925, w4926);
  FullAdder U1571 (w4926, w4829, IN53[28], w4927, w4928);
  FullAdder U1572 (w4928, w4831, IN54[27], w4929, w4930);
  FullAdder U1573 (w4930, w4833, IN55[26], w4931, w4932);
  FullAdder U1574 (w4932, w4835, IN56[25], w4933, w4934);
  FullAdder U1575 (w4934, w4837, IN57[24], w4935, w4936);
  FullAdder U1576 (w4936, w4839, IN58[23], w4937, w4938);
  FullAdder U1577 (w4938, w4841, IN59[22], w4939, w4940);
  FullAdder U1578 (w4940, w4843, IN60[21], w4941, w4942);
  FullAdder U1579 (w4942, w4845, IN61[20], w4943, w4944);
  FullAdder U1580 (w4944, w4847, IN62[19], w4945, w4946);
  FullAdder U1581 (w4946, w4849, IN63[18], w4947, w4948);
  FullAdder U1582 (w4948, w4851, IN64[17], w4949, w4950);
  FullAdder U1583 (w4950, w4853, IN65[16], w4951, w4952);
  FullAdder U1584 (w4952, w4855, IN66[15], w4953, w4954);
  FullAdder U1585 (w4954, w4857, IN67[14], w4955, w4956);
  FullAdder U1586 (w4956, w4859, IN68[13], w4957, w4958);
  FullAdder U1587 (w4958, w4861, IN69[12], w4959, w4960);
  FullAdder U1588 (w4960, w4863, IN70[11], w4961, w4962);
  FullAdder U1589 (w4962, w4865, IN71[10], w4963, w4964);
  FullAdder U1590 (w4964, w4867, IN72[9], w4965, w4966);
  FullAdder U1591 (w4966, w4869, IN73[8], w4967, w4968);
  FullAdder U1592 (w4968, w4871, IN74[7], w4969, w4970);
  FullAdder U1593 (w4970, w4873, IN75[6], w4971, w4972);
  FullAdder U1594 (w4972, w4875, IN76[5], w4973, w4974);
  FullAdder U1595 (w4974, w4877, IN77[4], w4975, w4976);
  FullAdder U1596 (w4976, w4879, IN78[3], w4977, w4978);
  FullAdder U1597 (w4978, w4881, IN79[2], w4979, w4980);
  FullAdder U1598 (w4980, w4883, IN80[1], w4981, w4982);
  FullAdder U1599 (w4982, w4884, IN81[0], w4983, w4984);
  HalfAdder U1600 (w4887, IN33[33], Out1[33], w4986);
  FullAdder U1601 (w4986, w4889, IN34[33], w4987, w4988);
  FullAdder U1602 (w4988, w4891, IN35[33], w4989, w4990);
  FullAdder U1603 (w4990, w4893, IN36[33], w4991, w4992);
  FullAdder U1604 (w4992, w4895, IN37[33], w4993, w4994);
  FullAdder U1605 (w4994, w4897, IN38[33], w4995, w4996);
  FullAdder U1606 (w4996, w4899, IN39[33], w4997, w4998);
  FullAdder U1607 (w4998, w4901, IN40[33], w4999, w5000);
  FullAdder U1608 (w5000, w4903, IN41[33], w5001, w5002);
  FullAdder U1609 (w5002, w4905, IN42[33], w5003, w5004);
  FullAdder U1610 (w5004, w4907, IN43[33], w5005, w5006);
  FullAdder U1611 (w5006, w4909, IN44[33], w5007, w5008);
  FullAdder U1612 (w5008, w4911, IN45[33], w5009, w5010);
  FullAdder U1613 (w5010, w4913, IN46[33], w5011, w5012);
  FullAdder U1614 (w5012, w4915, IN47[33], w5013, w5014);
  FullAdder U1615 (w5014, w4917, IN48[33], w5015, w5016);
  FullAdder U1616 (w5016, w4919, IN49[33], w5017, w5018);
  FullAdder U1617 (w5018, w4921, IN50[33], w5019, w5020);
  FullAdder U1618 (w5020, w4923, IN51[31], w5021, w5022);
  FullAdder U1619 (w5022, w4925, IN52[30], w5023, w5024);
  FullAdder U1620 (w5024, w4927, IN53[29], w5025, w5026);
  FullAdder U1621 (w5026, w4929, IN54[28], w5027, w5028);
  FullAdder U1622 (w5028, w4931, IN55[27], w5029, w5030);
  FullAdder U1623 (w5030, w4933, IN56[26], w5031, w5032);
  FullAdder U1624 (w5032, w4935, IN57[25], w5033, w5034);
  FullAdder U1625 (w5034, w4937, IN58[24], w5035, w5036);
  FullAdder U1626 (w5036, w4939, IN59[23], w5037, w5038);
  FullAdder U1627 (w5038, w4941, IN60[22], w5039, w5040);
  FullAdder U1628 (w5040, w4943, IN61[21], w5041, w5042);
  FullAdder U1629 (w5042, w4945, IN62[20], w5043, w5044);
  FullAdder U1630 (w5044, w4947, IN63[19], w5045, w5046);
  FullAdder U1631 (w5046, w4949, IN64[18], w5047, w5048);
  FullAdder U1632 (w5048, w4951, IN65[17], w5049, w5050);
  FullAdder U1633 (w5050, w4953, IN66[16], w5051, w5052);
  FullAdder U1634 (w5052, w4955, IN67[15], w5053, w5054);
  FullAdder U1635 (w5054, w4957, IN68[14], w5055, w5056);
  FullAdder U1636 (w5056, w4959, IN69[13], w5057, w5058);
  FullAdder U1637 (w5058, w4961, IN70[12], w5059, w5060);
  FullAdder U1638 (w5060, w4963, IN71[11], w5061, w5062);
  FullAdder U1639 (w5062, w4965, IN72[10], w5063, w5064);
  FullAdder U1640 (w5064, w4967, IN73[9], w5065, w5066);
  FullAdder U1641 (w5066, w4969, IN74[8], w5067, w5068);
  FullAdder U1642 (w5068, w4971, IN75[7], w5069, w5070);
  FullAdder U1643 (w5070, w4973, IN76[6], w5071, w5072);
  FullAdder U1644 (w5072, w4975, IN77[5], w5073, w5074);
  FullAdder U1645 (w5074, w4977, IN78[4], w5075, w5076);
  FullAdder U1646 (w5076, w4979, IN79[3], w5077, w5078);
  FullAdder U1647 (w5078, w4981, IN80[2], w5079, w5080);
  FullAdder U1648 (w5080, w4983, IN81[1], w5081, w5082);
  FullAdder U1649 (w5082, w4984, IN82[0], w5083, w5084);
  HalfAdder U1650 (w4987, IN34[34], Out1[34], w5086);
  FullAdder U1651 (w5086, w4989, IN35[34], Out1[35], w5088);
  FullAdder U1652 (w5088, w4991, IN36[34], Out1[36], w5090);
  FullAdder U1653 (w5090, w4993, IN37[34], Out1[37], w5092);
  FullAdder U1654 (w5092, w4995, IN38[34], Out1[38], w5094);
  FullAdder U1655 (w5094, w4997, IN39[34], Out1[39], w5096);
  FullAdder U1656 (w5096, w4999, IN40[34], Out1[40], w5098);
  FullAdder U1657 (w5098, w5001, IN41[34], Out1[41], w5100);
  FullAdder U1658 (w5100, w5003, IN42[34], Out1[42], w5102);
  FullAdder U1659 (w5102, w5005, IN43[34], Out1[43], w5104);
  FullAdder U1660 (w5104, w5007, IN44[34], Out1[44], w5106);
  FullAdder U1661 (w5106, w5009, IN45[34], Out1[45], w5108);
  FullAdder U1662 (w5108, w5011, IN46[34], Out1[46], w5110);
  FullAdder U1663 (w5110, w5013, IN47[34], Out1[47], w5112);
  FullAdder U1664 (w5112, w5015, IN48[34], Out1[48], w5114);
  FullAdder U1665 (w5114, w5017, IN49[34], Out1[49], w5116);
  FullAdder U1666 (w5116, w5019, IN50[34], Out1[50], w5118);
  FullAdder U1667 (w5118, w5021, IN51[32], Out1[51], w5120);
  FullAdder U1668 (w5120, w5023, IN52[31], Out1[52], w5122);
  FullAdder U1669 (w5122, w5025, IN53[30], Out1[53], w5124);
  FullAdder U1670 (w5124, w5027, IN54[29], Out1[54], w5126);
  FullAdder U1671 (w5126, w5029, IN55[28], Out1[55], w5128);
  FullAdder U1672 (w5128, w5031, IN56[27], Out1[56], w5130);
  FullAdder U1673 (w5130, w5033, IN57[26], Out1[57], w5132);
  FullAdder U1674 (w5132, w5035, IN58[25], Out1[58], w5134);
  FullAdder U1675 (w5134, w5037, IN59[24], Out1[59], w5136);
  FullAdder U1676 (w5136, w5039, IN60[23], Out1[60], w5138);
  FullAdder U1677 (w5138, w5041, IN61[22], Out1[61], w5140);
  FullAdder U1678 (w5140, w5043, IN62[21], Out1[62], w5142);
  FullAdder U1679 (w5142, w5045, IN63[20], Out1[63], w5144);
  FullAdder U1680 (w5144, w5047, IN64[19], Out1[64], w5146);
  FullAdder U1681 (w5146, w5049, IN65[18], Out1[65], w5148);
  FullAdder U1682 (w5148, w5051, IN66[17], Out1[66], w5150);
  FullAdder U1683 (w5150, w5053, IN67[16], Out1[67], w5152);
  FullAdder U1684 (w5152, w5055, IN68[15], Out1[68], w5154);
  FullAdder U1685 (w5154, w5057, IN69[14], Out1[69], w5156);
  FullAdder U1686 (w5156, w5059, IN70[13], Out1[70], w5158);
  FullAdder U1687 (w5158, w5061, IN71[12], Out1[71], w5160);
  FullAdder U1688 (w5160, w5063, IN72[11], Out1[72], w5162);
  FullAdder U1689 (w5162, w5065, IN73[10], Out1[73], w5164);
  FullAdder U1690 (w5164, w5067, IN74[9], Out1[74], w5166);
  FullAdder U1691 (w5166, w5069, IN75[8], Out1[75], w5168);
  FullAdder U1692 (w5168, w5071, IN76[7], Out1[76], w5170);
  FullAdder U1693 (w5170, w5073, IN77[6], Out1[77], w5172);
  FullAdder U1694 (w5172, w5075, IN78[5], Out1[78], w5174);
  FullAdder U1695 (w5174, w5077, IN79[4], Out1[79], w5176);
  FullAdder U1696 (w5176, w5079, IN80[3], Out1[80], w5178);
  FullAdder U1697 (w5178, w5081, IN81[2], Out1[81], w5180);
  FullAdder U1698 (w5180, w5083, IN82[1], Out1[82], w5182);
  FullAdder U1699 (w5182, w5084, IN83[0], Out1[83], Out1[84]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN51[33];
  assign Out2[1] = IN52[32];
  assign Out2[2] = IN53[31];
  assign Out2[3] = IN54[30];
  assign Out2[4] = IN55[29];
  assign Out2[5] = IN56[28];
  assign Out2[6] = IN57[27];
  assign Out2[7] = IN58[26];
  assign Out2[8] = IN59[25];
  assign Out2[9] = IN60[24];
  assign Out2[10] = IN61[23];
  assign Out2[11] = IN62[22];
  assign Out2[12] = IN63[21];
  assign Out2[13] = IN64[20];
  assign Out2[14] = IN65[19];
  assign Out2[15] = IN66[18];
  assign Out2[16] = IN67[17];
  assign Out2[17] = IN68[16];
  assign Out2[18] = IN69[15];
  assign Out2[19] = IN70[14];
  assign Out2[20] = IN71[13];
  assign Out2[21] = IN72[12];
  assign Out2[22] = IN73[11];
  assign Out2[23] = IN74[10];
  assign Out2[24] = IN75[9];
  assign Out2[25] = IN76[8];
  assign Out2[26] = IN77[7];
  assign Out2[27] = IN78[6];
  assign Out2[28] = IN79[5];
  assign Out2[29] = IN80[4];
  assign Out2[30] = IN81[3];
  assign Out2[31] = IN82[2];
  assign Out2[32] = IN83[1];
  assign Out2[33] = IN84[0];

endmodule
module RC_34_34(IN1, IN2, Out);
  input [33:0] IN1;
  input [33:0] IN2;
  output [34:0] Out;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w69);
  FullAdder U1 (IN1[1], IN2[1], w69, Out[1], w71);
  FullAdder U2 (IN1[2], IN2[2], w71, Out[2], w73);
  FullAdder U3 (IN1[3], IN2[3], w73, Out[3], w75);
  FullAdder U4 (IN1[4], IN2[4], w75, Out[4], w77);
  FullAdder U5 (IN1[5], IN2[5], w77, Out[5], w79);
  FullAdder U6 (IN1[6], IN2[6], w79, Out[6], w81);
  FullAdder U7 (IN1[7], IN2[7], w81, Out[7], w83);
  FullAdder U8 (IN1[8], IN2[8], w83, Out[8], w85);
  FullAdder U9 (IN1[9], IN2[9], w85, Out[9], w87);
  FullAdder U10 (IN1[10], IN2[10], w87, Out[10], w89);
  FullAdder U11 (IN1[11], IN2[11], w89, Out[11], w91);
  FullAdder U12 (IN1[12], IN2[12], w91, Out[12], w93);
  FullAdder U13 (IN1[13], IN2[13], w93, Out[13], w95);
  FullAdder U14 (IN1[14], IN2[14], w95, Out[14], w97);
  FullAdder U15 (IN1[15], IN2[15], w97, Out[15], w99);
  FullAdder U16 (IN1[16], IN2[16], w99, Out[16], w101);
  FullAdder U17 (IN1[17], IN2[17], w101, Out[17], w103);
  FullAdder U18 (IN1[18], IN2[18], w103, Out[18], w105);
  FullAdder U19 (IN1[19], IN2[19], w105, Out[19], w107);
  FullAdder U20 (IN1[20], IN2[20], w107, Out[20], w109);
  FullAdder U21 (IN1[21], IN2[21], w109, Out[21], w111);
  FullAdder U22 (IN1[22], IN2[22], w111, Out[22], w113);
  FullAdder U23 (IN1[23], IN2[23], w113, Out[23], w115);
  FullAdder U24 (IN1[24], IN2[24], w115, Out[24], w117);
  FullAdder U25 (IN1[25], IN2[25], w117, Out[25], w119);
  FullAdder U26 (IN1[26], IN2[26], w119, Out[26], w121);
  FullAdder U27 (IN1[27], IN2[27], w121, Out[27], w123);
  FullAdder U28 (IN1[28], IN2[28], w123, Out[28], w125);
  FullAdder U29 (IN1[29], IN2[29], w125, Out[29], w127);
  FullAdder U30 (IN1[30], IN2[30], w127, Out[30], w129);
  FullAdder U31 (IN1[31], IN2[31], w129, Out[31], w131);
  FullAdder U32 (IN1[32], IN2[32], w131, Out[32], w133);
  FullAdder U33 (IN1[33], IN2[33], w133, Out[33], Out[34]);

endmodule
module NR_51_35(IN1, IN2, Out);
  input [50:0] IN1;
  input [34:0] IN2;
  output [85:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [29:0] P29;
  wire [30:0] P30;
  wire [31:0] P31;
  wire [32:0] P32;
  wire [33:0] P33;
  wire [34:0] P34;
  wire [34:0] P35;
  wire [34:0] P36;
  wire [34:0] P37;
  wire [34:0] P38;
  wire [34:0] P39;
  wire [34:0] P40;
  wire [34:0] P41;
  wire [34:0] P42;
  wire [34:0] P43;
  wire [34:0] P44;
  wire [34:0] P45;
  wire [34:0] P46;
  wire [34:0] P47;
  wire [34:0] P48;
  wire [34:0] P49;
  wire [34:0] P50;
  wire [33:0] P51;
  wire [32:0] P52;
  wire [31:0] P53;
  wire [30:0] P54;
  wire [29:0] P55;
  wire [28:0] P56;
  wire [27:0] P57;
  wire [26:0] P58;
  wire [25:0] P59;
  wire [24:0] P60;
  wire [23:0] P61;
  wire [22:0] P62;
  wire [21:0] P63;
  wire [20:0] P64;
  wire [19:0] P65;
  wire [18:0] P66;
  wire [17:0] P67;
  wire [16:0] P68;
  wire [15:0] P69;
  wire [14:0] P70;
  wire [13:0] P71;
  wire [12:0] P72;
  wire [11:0] P73;
  wire [10:0] P74;
  wire [9:0] P75;
  wire [8:0] P76;
  wire [7:0] P77;
  wire [6:0] P78;
  wire [5:0] P79;
  wire [4:0] P80;
  wire [3:0] P81;
  wire [2:0] P82;
  wire [1:0] P83;
  wire [0:0] P84;
  wire [84:0] R1;
  wire [33:0] R2;
  wire [85:0] aOut;
  U_SP_51_35 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, R1, R2);
  RC_34_34 S2 (R1[84:51], R2, aOut[85:51]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign Out = aOut[85:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
