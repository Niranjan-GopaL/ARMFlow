//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 15
  second input length: 35
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_15_35(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48);
  input [14:0] IN1;
  input [34:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [14:0] P15;
  output [14:0] P16;
  output [14:0] P17;
  output [14:0] P18;
  output [14:0] P19;
  output [14:0] P20;
  output [14:0] P21;
  output [14:0] P22;
  output [14:0] P23;
  output [14:0] P24;
  output [14:0] P25;
  output [14:0] P26;
  output [14:0] P27;
  output [14:0] P28;
  output [14:0] P29;
  output [14:0] P30;
  output [14:0] P31;
  output [14:0] P32;
  output [14:0] P33;
  output [14:0] P34;
  output [13:0] P35;
  output [12:0] P36;
  output [11:0] P37;
  output [10:0] P38;
  output [9:0] P39;
  output [8:0] P40;
  output [7:0] P41;
  output [6:0] P42;
  output [5:0] P43;
  output [4:0] P44;
  output [3:0] P45;
  output [2:0] P46;
  output [1:0] P47;
  output [0:0] P48;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[0] = IN1[1]&IN2[34];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[1] = IN1[2]&IN2[33];
  assign P36[0] = IN1[2]&IN2[34];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[2] = IN1[3]&IN2[32];
  assign P36[1] = IN1[3]&IN2[33];
  assign P37[0] = IN1[3]&IN2[34];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[3] = IN1[4]&IN2[31];
  assign P36[2] = IN1[4]&IN2[32];
  assign P37[1] = IN1[4]&IN2[33];
  assign P38[0] = IN1[4]&IN2[34];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[4] = IN1[5]&IN2[30];
  assign P36[3] = IN1[5]&IN2[31];
  assign P37[2] = IN1[5]&IN2[32];
  assign P38[1] = IN1[5]&IN2[33];
  assign P39[0] = IN1[5]&IN2[34];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[5] = IN1[6]&IN2[29];
  assign P36[4] = IN1[6]&IN2[30];
  assign P37[3] = IN1[6]&IN2[31];
  assign P38[2] = IN1[6]&IN2[32];
  assign P39[1] = IN1[6]&IN2[33];
  assign P40[0] = IN1[6]&IN2[34];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[6] = IN1[7]&IN2[28];
  assign P36[5] = IN1[7]&IN2[29];
  assign P37[4] = IN1[7]&IN2[30];
  assign P38[3] = IN1[7]&IN2[31];
  assign P39[2] = IN1[7]&IN2[32];
  assign P40[1] = IN1[7]&IN2[33];
  assign P41[0] = IN1[7]&IN2[34];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[7] = IN1[8]&IN2[27];
  assign P36[6] = IN1[8]&IN2[28];
  assign P37[5] = IN1[8]&IN2[29];
  assign P38[4] = IN1[8]&IN2[30];
  assign P39[3] = IN1[8]&IN2[31];
  assign P40[2] = IN1[8]&IN2[32];
  assign P41[1] = IN1[8]&IN2[33];
  assign P42[0] = IN1[8]&IN2[34];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[8] = IN1[9]&IN2[26];
  assign P36[7] = IN1[9]&IN2[27];
  assign P37[6] = IN1[9]&IN2[28];
  assign P38[5] = IN1[9]&IN2[29];
  assign P39[4] = IN1[9]&IN2[30];
  assign P40[3] = IN1[9]&IN2[31];
  assign P41[2] = IN1[9]&IN2[32];
  assign P42[1] = IN1[9]&IN2[33];
  assign P43[0] = IN1[9]&IN2[34];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[9] = IN1[10]&IN2[25];
  assign P36[8] = IN1[10]&IN2[26];
  assign P37[7] = IN1[10]&IN2[27];
  assign P38[6] = IN1[10]&IN2[28];
  assign P39[5] = IN1[10]&IN2[29];
  assign P40[4] = IN1[10]&IN2[30];
  assign P41[3] = IN1[10]&IN2[31];
  assign P42[2] = IN1[10]&IN2[32];
  assign P43[1] = IN1[10]&IN2[33];
  assign P44[0] = IN1[10]&IN2[34];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[10] = IN1[11]&IN2[24];
  assign P36[9] = IN1[11]&IN2[25];
  assign P37[8] = IN1[11]&IN2[26];
  assign P38[7] = IN1[11]&IN2[27];
  assign P39[6] = IN1[11]&IN2[28];
  assign P40[5] = IN1[11]&IN2[29];
  assign P41[4] = IN1[11]&IN2[30];
  assign P42[3] = IN1[11]&IN2[31];
  assign P43[2] = IN1[11]&IN2[32];
  assign P44[1] = IN1[11]&IN2[33];
  assign P45[0] = IN1[11]&IN2[34];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[11] = IN1[12]&IN2[23];
  assign P36[10] = IN1[12]&IN2[24];
  assign P37[9] = IN1[12]&IN2[25];
  assign P38[8] = IN1[12]&IN2[26];
  assign P39[7] = IN1[12]&IN2[27];
  assign P40[6] = IN1[12]&IN2[28];
  assign P41[5] = IN1[12]&IN2[29];
  assign P42[4] = IN1[12]&IN2[30];
  assign P43[3] = IN1[12]&IN2[31];
  assign P44[2] = IN1[12]&IN2[32];
  assign P45[1] = IN1[12]&IN2[33];
  assign P46[0] = IN1[12]&IN2[34];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[12] = IN1[13]&IN2[22];
  assign P36[11] = IN1[13]&IN2[23];
  assign P37[10] = IN1[13]&IN2[24];
  assign P38[9] = IN1[13]&IN2[25];
  assign P39[8] = IN1[13]&IN2[26];
  assign P40[7] = IN1[13]&IN2[27];
  assign P41[6] = IN1[13]&IN2[28];
  assign P42[5] = IN1[13]&IN2[29];
  assign P43[4] = IN1[13]&IN2[30];
  assign P44[3] = IN1[13]&IN2[31];
  assign P45[2] = IN1[13]&IN2[32];
  assign P46[1] = IN1[13]&IN2[33];
  assign P47[0] = IN1[13]&IN2[34];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[13] = IN1[14]&IN2[21];
  assign P36[12] = IN1[14]&IN2[22];
  assign P37[11] = IN1[14]&IN2[23];
  assign P38[10] = IN1[14]&IN2[24];
  assign P39[9] = IN1[14]&IN2[25];
  assign P40[8] = IN1[14]&IN2[26];
  assign P41[7] = IN1[14]&IN2[27];
  assign P42[6] = IN1[14]&IN2[28];
  assign P43[5] = IN1[14]&IN2[29];
  assign P44[4] = IN1[14]&IN2[30];
  assign P45[3] = IN1[14]&IN2[31];
  assign P46[2] = IN1[14]&IN2[32];
  assign P47[1] = IN1[14]&IN2[33];
  assign P48[0] = IN1[14]&IN2[34];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [14:0] IN15;
  input [14:0] IN16;
  input [14:0] IN17;
  input [14:0] IN18;
  input [14:0] IN19;
  input [14:0] IN20;
  input [14:0] IN21;
  input [14:0] IN22;
  input [14:0] IN23;
  input [14:0] IN24;
  input [14:0] IN25;
  input [14:0] IN26;
  input [14:0] IN27;
  input [14:0] IN28;
  input [14:0] IN29;
  input [14:0] IN30;
  input [14:0] IN31;
  input [14:0] IN32;
  input [14:0] IN33;
  input [14:0] IN34;
  input [13:0] IN35;
  input [12:0] IN36;
  input [11:0] IN37;
  input [10:0] IN38;
  input [9:0] IN39;
  input [8:0] IN40;
  input [7:0] IN41;
  input [6:0] IN42;
  input [5:0] IN43;
  input [4:0] IN44;
  input [3:0] IN45;
  input [2:0] IN46;
  input [1:0] IN47;
  input [0:0] IN48;
  output [48:0] Out1;
  output [33:0] Out2;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1450;
  wire w1452;
  wire w1454;
  wire w1456;
  wire w1458;
  wire w1460;
  wire w1462;
  wire w1464;
  wire w1466;
  wire w1468;
  wire w1470;
  wire w1472;
  wire w1474;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w526);
  FullAdder U1 (w526, IN2[0], IN2[1], w527, w528);
  FullAdder U2 (w528, IN3[0], IN3[1], w529, w530);
  FullAdder U3 (w530, IN4[0], IN4[1], w531, w532);
  FullAdder U4 (w532, IN5[0], IN5[1], w533, w534);
  FullAdder U5 (w534, IN6[0], IN6[1], w535, w536);
  FullAdder U6 (w536, IN7[0], IN7[1], w537, w538);
  FullAdder U7 (w538, IN8[0], IN8[1], w539, w540);
  FullAdder U8 (w540, IN9[0], IN9[1], w541, w542);
  FullAdder U9 (w542, IN10[0], IN10[1], w543, w544);
  FullAdder U10 (w544, IN11[0], IN11[1], w545, w546);
  FullAdder U11 (w546, IN12[0], IN12[1], w547, w548);
  FullAdder U12 (w548, IN13[0], IN13[1], w549, w550);
  FullAdder U13 (w550, IN14[0], IN14[1], w551, w552);
  HalfAdder U14 (w527, IN2[2], Out1[2], w554);
  FullAdder U15 (w554, w529, IN3[2], w555, w556);
  FullAdder U16 (w556, w531, IN4[2], w557, w558);
  FullAdder U17 (w558, w533, IN5[2], w559, w560);
  FullAdder U18 (w560, w535, IN6[2], w561, w562);
  FullAdder U19 (w562, w537, IN7[2], w563, w564);
  FullAdder U20 (w564, w539, IN8[2], w565, w566);
  FullAdder U21 (w566, w541, IN9[2], w567, w568);
  FullAdder U22 (w568, w543, IN10[2], w569, w570);
  FullAdder U23 (w570, w545, IN11[2], w571, w572);
  FullAdder U24 (w572, w547, IN12[2], w573, w574);
  FullAdder U25 (w574, w549, IN13[2], w575, w576);
  FullAdder U26 (w576, w551, IN14[2], w577, w578);
  FullAdder U27 (w578, w552, IN15[0], w579, w580);
  HalfAdder U28 (w555, IN3[3], Out1[3], w582);
  FullAdder U29 (w582, w557, IN4[3], w583, w584);
  FullAdder U30 (w584, w559, IN5[3], w585, w586);
  FullAdder U31 (w586, w561, IN6[3], w587, w588);
  FullAdder U32 (w588, w563, IN7[3], w589, w590);
  FullAdder U33 (w590, w565, IN8[3], w591, w592);
  FullAdder U34 (w592, w567, IN9[3], w593, w594);
  FullAdder U35 (w594, w569, IN10[3], w595, w596);
  FullAdder U36 (w596, w571, IN11[3], w597, w598);
  FullAdder U37 (w598, w573, IN12[3], w599, w600);
  FullAdder U38 (w600, w575, IN13[3], w601, w602);
  FullAdder U39 (w602, w577, IN14[3], w603, w604);
  FullAdder U40 (w604, w579, IN15[1], w605, w606);
  FullAdder U41 (w606, w580, IN16[0], w607, w608);
  HalfAdder U42 (w583, IN4[4], Out1[4], w610);
  FullAdder U43 (w610, w585, IN5[4], w611, w612);
  FullAdder U44 (w612, w587, IN6[4], w613, w614);
  FullAdder U45 (w614, w589, IN7[4], w615, w616);
  FullAdder U46 (w616, w591, IN8[4], w617, w618);
  FullAdder U47 (w618, w593, IN9[4], w619, w620);
  FullAdder U48 (w620, w595, IN10[4], w621, w622);
  FullAdder U49 (w622, w597, IN11[4], w623, w624);
  FullAdder U50 (w624, w599, IN12[4], w625, w626);
  FullAdder U51 (w626, w601, IN13[4], w627, w628);
  FullAdder U52 (w628, w603, IN14[4], w629, w630);
  FullAdder U53 (w630, w605, IN15[2], w631, w632);
  FullAdder U54 (w632, w607, IN16[1], w633, w634);
  FullAdder U55 (w634, w608, IN17[0], w635, w636);
  HalfAdder U56 (w611, IN5[5], Out1[5], w638);
  FullAdder U57 (w638, w613, IN6[5], w639, w640);
  FullAdder U58 (w640, w615, IN7[5], w641, w642);
  FullAdder U59 (w642, w617, IN8[5], w643, w644);
  FullAdder U60 (w644, w619, IN9[5], w645, w646);
  FullAdder U61 (w646, w621, IN10[5], w647, w648);
  FullAdder U62 (w648, w623, IN11[5], w649, w650);
  FullAdder U63 (w650, w625, IN12[5], w651, w652);
  FullAdder U64 (w652, w627, IN13[5], w653, w654);
  FullAdder U65 (w654, w629, IN14[5], w655, w656);
  FullAdder U66 (w656, w631, IN15[3], w657, w658);
  FullAdder U67 (w658, w633, IN16[2], w659, w660);
  FullAdder U68 (w660, w635, IN17[1], w661, w662);
  FullAdder U69 (w662, w636, IN18[0], w663, w664);
  HalfAdder U70 (w639, IN6[6], Out1[6], w666);
  FullAdder U71 (w666, w641, IN7[6], w667, w668);
  FullAdder U72 (w668, w643, IN8[6], w669, w670);
  FullAdder U73 (w670, w645, IN9[6], w671, w672);
  FullAdder U74 (w672, w647, IN10[6], w673, w674);
  FullAdder U75 (w674, w649, IN11[6], w675, w676);
  FullAdder U76 (w676, w651, IN12[6], w677, w678);
  FullAdder U77 (w678, w653, IN13[6], w679, w680);
  FullAdder U78 (w680, w655, IN14[6], w681, w682);
  FullAdder U79 (w682, w657, IN15[4], w683, w684);
  FullAdder U80 (w684, w659, IN16[3], w685, w686);
  FullAdder U81 (w686, w661, IN17[2], w687, w688);
  FullAdder U82 (w688, w663, IN18[1], w689, w690);
  FullAdder U83 (w690, w664, IN19[0], w691, w692);
  HalfAdder U84 (w667, IN7[7], Out1[7], w694);
  FullAdder U85 (w694, w669, IN8[7], w695, w696);
  FullAdder U86 (w696, w671, IN9[7], w697, w698);
  FullAdder U87 (w698, w673, IN10[7], w699, w700);
  FullAdder U88 (w700, w675, IN11[7], w701, w702);
  FullAdder U89 (w702, w677, IN12[7], w703, w704);
  FullAdder U90 (w704, w679, IN13[7], w705, w706);
  FullAdder U91 (w706, w681, IN14[7], w707, w708);
  FullAdder U92 (w708, w683, IN15[5], w709, w710);
  FullAdder U93 (w710, w685, IN16[4], w711, w712);
  FullAdder U94 (w712, w687, IN17[3], w713, w714);
  FullAdder U95 (w714, w689, IN18[2], w715, w716);
  FullAdder U96 (w716, w691, IN19[1], w717, w718);
  FullAdder U97 (w718, w692, IN20[0], w719, w720);
  HalfAdder U98 (w695, IN8[8], Out1[8], w722);
  FullAdder U99 (w722, w697, IN9[8], w723, w724);
  FullAdder U100 (w724, w699, IN10[8], w725, w726);
  FullAdder U101 (w726, w701, IN11[8], w727, w728);
  FullAdder U102 (w728, w703, IN12[8], w729, w730);
  FullAdder U103 (w730, w705, IN13[8], w731, w732);
  FullAdder U104 (w732, w707, IN14[8], w733, w734);
  FullAdder U105 (w734, w709, IN15[6], w735, w736);
  FullAdder U106 (w736, w711, IN16[5], w737, w738);
  FullAdder U107 (w738, w713, IN17[4], w739, w740);
  FullAdder U108 (w740, w715, IN18[3], w741, w742);
  FullAdder U109 (w742, w717, IN19[2], w743, w744);
  FullAdder U110 (w744, w719, IN20[1], w745, w746);
  FullAdder U111 (w746, w720, IN21[0], w747, w748);
  HalfAdder U112 (w723, IN9[9], Out1[9], w750);
  FullAdder U113 (w750, w725, IN10[9], w751, w752);
  FullAdder U114 (w752, w727, IN11[9], w753, w754);
  FullAdder U115 (w754, w729, IN12[9], w755, w756);
  FullAdder U116 (w756, w731, IN13[9], w757, w758);
  FullAdder U117 (w758, w733, IN14[9], w759, w760);
  FullAdder U118 (w760, w735, IN15[7], w761, w762);
  FullAdder U119 (w762, w737, IN16[6], w763, w764);
  FullAdder U120 (w764, w739, IN17[5], w765, w766);
  FullAdder U121 (w766, w741, IN18[4], w767, w768);
  FullAdder U122 (w768, w743, IN19[3], w769, w770);
  FullAdder U123 (w770, w745, IN20[2], w771, w772);
  FullAdder U124 (w772, w747, IN21[1], w773, w774);
  FullAdder U125 (w774, w748, IN22[0], w775, w776);
  HalfAdder U126 (w751, IN10[10], Out1[10], w778);
  FullAdder U127 (w778, w753, IN11[10], w779, w780);
  FullAdder U128 (w780, w755, IN12[10], w781, w782);
  FullAdder U129 (w782, w757, IN13[10], w783, w784);
  FullAdder U130 (w784, w759, IN14[10], w785, w786);
  FullAdder U131 (w786, w761, IN15[8], w787, w788);
  FullAdder U132 (w788, w763, IN16[7], w789, w790);
  FullAdder U133 (w790, w765, IN17[6], w791, w792);
  FullAdder U134 (w792, w767, IN18[5], w793, w794);
  FullAdder U135 (w794, w769, IN19[4], w795, w796);
  FullAdder U136 (w796, w771, IN20[3], w797, w798);
  FullAdder U137 (w798, w773, IN21[2], w799, w800);
  FullAdder U138 (w800, w775, IN22[1], w801, w802);
  FullAdder U139 (w802, w776, IN23[0], w803, w804);
  HalfAdder U140 (w779, IN11[11], Out1[11], w806);
  FullAdder U141 (w806, w781, IN12[11], w807, w808);
  FullAdder U142 (w808, w783, IN13[11], w809, w810);
  FullAdder U143 (w810, w785, IN14[11], w811, w812);
  FullAdder U144 (w812, w787, IN15[9], w813, w814);
  FullAdder U145 (w814, w789, IN16[8], w815, w816);
  FullAdder U146 (w816, w791, IN17[7], w817, w818);
  FullAdder U147 (w818, w793, IN18[6], w819, w820);
  FullAdder U148 (w820, w795, IN19[5], w821, w822);
  FullAdder U149 (w822, w797, IN20[4], w823, w824);
  FullAdder U150 (w824, w799, IN21[3], w825, w826);
  FullAdder U151 (w826, w801, IN22[2], w827, w828);
  FullAdder U152 (w828, w803, IN23[1], w829, w830);
  FullAdder U153 (w830, w804, IN24[0], w831, w832);
  HalfAdder U154 (w807, IN12[12], Out1[12], w834);
  FullAdder U155 (w834, w809, IN13[12], w835, w836);
  FullAdder U156 (w836, w811, IN14[12], w837, w838);
  FullAdder U157 (w838, w813, IN15[10], w839, w840);
  FullAdder U158 (w840, w815, IN16[9], w841, w842);
  FullAdder U159 (w842, w817, IN17[8], w843, w844);
  FullAdder U160 (w844, w819, IN18[7], w845, w846);
  FullAdder U161 (w846, w821, IN19[6], w847, w848);
  FullAdder U162 (w848, w823, IN20[5], w849, w850);
  FullAdder U163 (w850, w825, IN21[4], w851, w852);
  FullAdder U164 (w852, w827, IN22[3], w853, w854);
  FullAdder U165 (w854, w829, IN23[2], w855, w856);
  FullAdder U166 (w856, w831, IN24[1], w857, w858);
  FullAdder U167 (w858, w832, IN25[0], w859, w860);
  HalfAdder U168 (w835, IN13[13], Out1[13], w862);
  FullAdder U169 (w862, w837, IN14[13], w863, w864);
  FullAdder U170 (w864, w839, IN15[11], w865, w866);
  FullAdder U171 (w866, w841, IN16[10], w867, w868);
  FullAdder U172 (w868, w843, IN17[9], w869, w870);
  FullAdder U173 (w870, w845, IN18[8], w871, w872);
  FullAdder U174 (w872, w847, IN19[7], w873, w874);
  FullAdder U175 (w874, w849, IN20[6], w875, w876);
  FullAdder U176 (w876, w851, IN21[5], w877, w878);
  FullAdder U177 (w878, w853, IN22[4], w879, w880);
  FullAdder U178 (w880, w855, IN23[3], w881, w882);
  FullAdder U179 (w882, w857, IN24[2], w883, w884);
  FullAdder U180 (w884, w859, IN25[1], w885, w886);
  FullAdder U181 (w886, w860, IN26[0], w887, w888);
  HalfAdder U182 (w863, IN14[14], Out1[14], w890);
  FullAdder U183 (w890, w865, IN15[12], w891, w892);
  FullAdder U184 (w892, w867, IN16[11], w893, w894);
  FullAdder U185 (w894, w869, IN17[10], w895, w896);
  FullAdder U186 (w896, w871, IN18[9], w897, w898);
  FullAdder U187 (w898, w873, IN19[8], w899, w900);
  FullAdder U188 (w900, w875, IN20[7], w901, w902);
  FullAdder U189 (w902, w877, IN21[6], w903, w904);
  FullAdder U190 (w904, w879, IN22[5], w905, w906);
  FullAdder U191 (w906, w881, IN23[4], w907, w908);
  FullAdder U192 (w908, w883, IN24[3], w909, w910);
  FullAdder U193 (w910, w885, IN25[2], w911, w912);
  FullAdder U194 (w912, w887, IN26[1], w913, w914);
  FullAdder U195 (w914, w888, IN27[0], w915, w916);
  HalfAdder U196 (w891, IN15[13], Out1[15], w918);
  FullAdder U197 (w918, w893, IN16[12], w919, w920);
  FullAdder U198 (w920, w895, IN17[11], w921, w922);
  FullAdder U199 (w922, w897, IN18[10], w923, w924);
  FullAdder U200 (w924, w899, IN19[9], w925, w926);
  FullAdder U201 (w926, w901, IN20[8], w927, w928);
  FullAdder U202 (w928, w903, IN21[7], w929, w930);
  FullAdder U203 (w930, w905, IN22[6], w931, w932);
  FullAdder U204 (w932, w907, IN23[5], w933, w934);
  FullAdder U205 (w934, w909, IN24[4], w935, w936);
  FullAdder U206 (w936, w911, IN25[3], w937, w938);
  FullAdder U207 (w938, w913, IN26[2], w939, w940);
  FullAdder U208 (w940, w915, IN27[1], w941, w942);
  FullAdder U209 (w942, w916, IN28[0], w943, w944);
  HalfAdder U210 (w919, IN16[13], Out1[16], w946);
  FullAdder U211 (w946, w921, IN17[12], w947, w948);
  FullAdder U212 (w948, w923, IN18[11], w949, w950);
  FullAdder U213 (w950, w925, IN19[10], w951, w952);
  FullAdder U214 (w952, w927, IN20[9], w953, w954);
  FullAdder U215 (w954, w929, IN21[8], w955, w956);
  FullAdder U216 (w956, w931, IN22[7], w957, w958);
  FullAdder U217 (w958, w933, IN23[6], w959, w960);
  FullAdder U218 (w960, w935, IN24[5], w961, w962);
  FullAdder U219 (w962, w937, IN25[4], w963, w964);
  FullAdder U220 (w964, w939, IN26[3], w965, w966);
  FullAdder U221 (w966, w941, IN27[2], w967, w968);
  FullAdder U222 (w968, w943, IN28[1], w969, w970);
  FullAdder U223 (w970, w944, IN29[0], w971, w972);
  HalfAdder U224 (w947, IN17[13], Out1[17], w974);
  FullAdder U225 (w974, w949, IN18[12], w975, w976);
  FullAdder U226 (w976, w951, IN19[11], w977, w978);
  FullAdder U227 (w978, w953, IN20[10], w979, w980);
  FullAdder U228 (w980, w955, IN21[9], w981, w982);
  FullAdder U229 (w982, w957, IN22[8], w983, w984);
  FullAdder U230 (w984, w959, IN23[7], w985, w986);
  FullAdder U231 (w986, w961, IN24[6], w987, w988);
  FullAdder U232 (w988, w963, IN25[5], w989, w990);
  FullAdder U233 (w990, w965, IN26[4], w991, w992);
  FullAdder U234 (w992, w967, IN27[3], w993, w994);
  FullAdder U235 (w994, w969, IN28[2], w995, w996);
  FullAdder U236 (w996, w971, IN29[1], w997, w998);
  FullAdder U237 (w998, w972, IN30[0], w999, w1000);
  HalfAdder U238 (w975, IN18[13], Out1[18], w1002);
  FullAdder U239 (w1002, w977, IN19[12], w1003, w1004);
  FullAdder U240 (w1004, w979, IN20[11], w1005, w1006);
  FullAdder U241 (w1006, w981, IN21[10], w1007, w1008);
  FullAdder U242 (w1008, w983, IN22[9], w1009, w1010);
  FullAdder U243 (w1010, w985, IN23[8], w1011, w1012);
  FullAdder U244 (w1012, w987, IN24[7], w1013, w1014);
  FullAdder U245 (w1014, w989, IN25[6], w1015, w1016);
  FullAdder U246 (w1016, w991, IN26[5], w1017, w1018);
  FullAdder U247 (w1018, w993, IN27[4], w1019, w1020);
  FullAdder U248 (w1020, w995, IN28[3], w1021, w1022);
  FullAdder U249 (w1022, w997, IN29[2], w1023, w1024);
  FullAdder U250 (w1024, w999, IN30[1], w1025, w1026);
  FullAdder U251 (w1026, w1000, IN31[0], w1027, w1028);
  HalfAdder U252 (w1003, IN19[13], Out1[19], w1030);
  FullAdder U253 (w1030, w1005, IN20[12], w1031, w1032);
  FullAdder U254 (w1032, w1007, IN21[11], w1033, w1034);
  FullAdder U255 (w1034, w1009, IN22[10], w1035, w1036);
  FullAdder U256 (w1036, w1011, IN23[9], w1037, w1038);
  FullAdder U257 (w1038, w1013, IN24[8], w1039, w1040);
  FullAdder U258 (w1040, w1015, IN25[7], w1041, w1042);
  FullAdder U259 (w1042, w1017, IN26[6], w1043, w1044);
  FullAdder U260 (w1044, w1019, IN27[5], w1045, w1046);
  FullAdder U261 (w1046, w1021, IN28[4], w1047, w1048);
  FullAdder U262 (w1048, w1023, IN29[3], w1049, w1050);
  FullAdder U263 (w1050, w1025, IN30[2], w1051, w1052);
  FullAdder U264 (w1052, w1027, IN31[1], w1053, w1054);
  FullAdder U265 (w1054, w1028, IN32[0], w1055, w1056);
  HalfAdder U266 (w1031, IN20[13], Out1[20], w1058);
  FullAdder U267 (w1058, w1033, IN21[12], w1059, w1060);
  FullAdder U268 (w1060, w1035, IN22[11], w1061, w1062);
  FullAdder U269 (w1062, w1037, IN23[10], w1063, w1064);
  FullAdder U270 (w1064, w1039, IN24[9], w1065, w1066);
  FullAdder U271 (w1066, w1041, IN25[8], w1067, w1068);
  FullAdder U272 (w1068, w1043, IN26[7], w1069, w1070);
  FullAdder U273 (w1070, w1045, IN27[6], w1071, w1072);
  FullAdder U274 (w1072, w1047, IN28[5], w1073, w1074);
  FullAdder U275 (w1074, w1049, IN29[4], w1075, w1076);
  FullAdder U276 (w1076, w1051, IN30[3], w1077, w1078);
  FullAdder U277 (w1078, w1053, IN31[2], w1079, w1080);
  FullAdder U278 (w1080, w1055, IN32[1], w1081, w1082);
  FullAdder U279 (w1082, w1056, IN33[0], w1083, w1084);
  HalfAdder U280 (w1059, IN21[13], Out1[21], w1086);
  FullAdder U281 (w1086, w1061, IN22[12], w1087, w1088);
  FullAdder U282 (w1088, w1063, IN23[11], w1089, w1090);
  FullAdder U283 (w1090, w1065, IN24[10], w1091, w1092);
  FullAdder U284 (w1092, w1067, IN25[9], w1093, w1094);
  FullAdder U285 (w1094, w1069, IN26[8], w1095, w1096);
  FullAdder U286 (w1096, w1071, IN27[7], w1097, w1098);
  FullAdder U287 (w1098, w1073, IN28[6], w1099, w1100);
  FullAdder U288 (w1100, w1075, IN29[5], w1101, w1102);
  FullAdder U289 (w1102, w1077, IN30[4], w1103, w1104);
  FullAdder U290 (w1104, w1079, IN31[3], w1105, w1106);
  FullAdder U291 (w1106, w1081, IN32[2], w1107, w1108);
  FullAdder U292 (w1108, w1083, IN33[1], w1109, w1110);
  FullAdder U293 (w1110, w1084, IN34[0], w1111, w1112);
  HalfAdder U294 (w1087, IN22[13], Out1[22], w1114);
  FullAdder U295 (w1114, w1089, IN23[12], w1115, w1116);
  FullAdder U296 (w1116, w1091, IN24[11], w1117, w1118);
  FullAdder U297 (w1118, w1093, IN25[10], w1119, w1120);
  FullAdder U298 (w1120, w1095, IN26[9], w1121, w1122);
  FullAdder U299 (w1122, w1097, IN27[8], w1123, w1124);
  FullAdder U300 (w1124, w1099, IN28[7], w1125, w1126);
  FullAdder U301 (w1126, w1101, IN29[6], w1127, w1128);
  FullAdder U302 (w1128, w1103, IN30[5], w1129, w1130);
  FullAdder U303 (w1130, w1105, IN31[4], w1131, w1132);
  FullAdder U304 (w1132, w1107, IN32[3], w1133, w1134);
  FullAdder U305 (w1134, w1109, IN33[2], w1135, w1136);
  FullAdder U306 (w1136, w1111, IN34[1], w1137, w1138);
  FullAdder U307 (w1138, w1112, IN35[0], w1139, w1140);
  HalfAdder U308 (w1115, IN23[13], Out1[23], w1142);
  FullAdder U309 (w1142, w1117, IN24[12], w1143, w1144);
  FullAdder U310 (w1144, w1119, IN25[11], w1145, w1146);
  FullAdder U311 (w1146, w1121, IN26[10], w1147, w1148);
  FullAdder U312 (w1148, w1123, IN27[9], w1149, w1150);
  FullAdder U313 (w1150, w1125, IN28[8], w1151, w1152);
  FullAdder U314 (w1152, w1127, IN29[7], w1153, w1154);
  FullAdder U315 (w1154, w1129, IN30[6], w1155, w1156);
  FullAdder U316 (w1156, w1131, IN31[5], w1157, w1158);
  FullAdder U317 (w1158, w1133, IN32[4], w1159, w1160);
  FullAdder U318 (w1160, w1135, IN33[3], w1161, w1162);
  FullAdder U319 (w1162, w1137, IN34[2], w1163, w1164);
  FullAdder U320 (w1164, w1139, IN35[1], w1165, w1166);
  FullAdder U321 (w1166, w1140, IN36[0], w1167, w1168);
  HalfAdder U322 (w1143, IN24[13], Out1[24], w1170);
  FullAdder U323 (w1170, w1145, IN25[12], w1171, w1172);
  FullAdder U324 (w1172, w1147, IN26[11], w1173, w1174);
  FullAdder U325 (w1174, w1149, IN27[10], w1175, w1176);
  FullAdder U326 (w1176, w1151, IN28[9], w1177, w1178);
  FullAdder U327 (w1178, w1153, IN29[8], w1179, w1180);
  FullAdder U328 (w1180, w1155, IN30[7], w1181, w1182);
  FullAdder U329 (w1182, w1157, IN31[6], w1183, w1184);
  FullAdder U330 (w1184, w1159, IN32[5], w1185, w1186);
  FullAdder U331 (w1186, w1161, IN33[4], w1187, w1188);
  FullAdder U332 (w1188, w1163, IN34[3], w1189, w1190);
  FullAdder U333 (w1190, w1165, IN35[2], w1191, w1192);
  FullAdder U334 (w1192, w1167, IN36[1], w1193, w1194);
  FullAdder U335 (w1194, w1168, IN37[0], w1195, w1196);
  HalfAdder U336 (w1171, IN25[13], Out1[25], w1198);
  FullAdder U337 (w1198, w1173, IN26[12], w1199, w1200);
  FullAdder U338 (w1200, w1175, IN27[11], w1201, w1202);
  FullAdder U339 (w1202, w1177, IN28[10], w1203, w1204);
  FullAdder U340 (w1204, w1179, IN29[9], w1205, w1206);
  FullAdder U341 (w1206, w1181, IN30[8], w1207, w1208);
  FullAdder U342 (w1208, w1183, IN31[7], w1209, w1210);
  FullAdder U343 (w1210, w1185, IN32[6], w1211, w1212);
  FullAdder U344 (w1212, w1187, IN33[5], w1213, w1214);
  FullAdder U345 (w1214, w1189, IN34[4], w1215, w1216);
  FullAdder U346 (w1216, w1191, IN35[3], w1217, w1218);
  FullAdder U347 (w1218, w1193, IN36[2], w1219, w1220);
  FullAdder U348 (w1220, w1195, IN37[1], w1221, w1222);
  FullAdder U349 (w1222, w1196, IN38[0], w1223, w1224);
  HalfAdder U350 (w1199, IN26[13], Out1[26], w1226);
  FullAdder U351 (w1226, w1201, IN27[12], w1227, w1228);
  FullAdder U352 (w1228, w1203, IN28[11], w1229, w1230);
  FullAdder U353 (w1230, w1205, IN29[10], w1231, w1232);
  FullAdder U354 (w1232, w1207, IN30[9], w1233, w1234);
  FullAdder U355 (w1234, w1209, IN31[8], w1235, w1236);
  FullAdder U356 (w1236, w1211, IN32[7], w1237, w1238);
  FullAdder U357 (w1238, w1213, IN33[6], w1239, w1240);
  FullAdder U358 (w1240, w1215, IN34[5], w1241, w1242);
  FullAdder U359 (w1242, w1217, IN35[4], w1243, w1244);
  FullAdder U360 (w1244, w1219, IN36[3], w1245, w1246);
  FullAdder U361 (w1246, w1221, IN37[2], w1247, w1248);
  FullAdder U362 (w1248, w1223, IN38[1], w1249, w1250);
  FullAdder U363 (w1250, w1224, IN39[0], w1251, w1252);
  HalfAdder U364 (w1227, IN27[13], Out1[27], w1254);
  FullAdder U365 (w1254, w1229, IN28[12], w1255, w1256);
  FullAdder U366 (w1256, w1231, IN29[11], w1257, w1258);
  FullAdder U367 (w1258, w1233, IN30[10], w1259, w1260);
  FullAdder U368 (w1260, w1235, IN31[9], w1261, w1262);
  FullAdder U369 (w1262, w1237, IN32[8], w1263, w1264);
  FullAdder U370 (w1264, w1239, IN33[7], w1265, w1266);
  FullAdder U371 (w1266, w1241, IN34[6], w1267, w1268);
  FullAdder U372 (w1268, w1243, IN35[5], w1269, w1270);
  FullAdder U373 (w1270, w1245, IN36[4], w1271, w1272);
  FullAdder U374 (w1272, w1247, IN37[3], w1273, w1274);
  FullAdder U375 (w1274, w1249, IN38[2], w1275, w1276);
  FullAdder U376 (w1276, w1251, IN39[1], w1277, w1278);
  FullAdder U377 (w1278, w1252, IN40[0], w1279, w1280);
  HalfAdder U378 (w1255, IN28[13], Out1[28], w1282);
  FullAdder U379 (w1282, w1257, IN29[12], w1283, w1284);
  FullAdder U380 (w1284, w1259, IN30[11], w1285, w1286);
  FullAdder U381 (w1286, w1261, IN31[10], w1287, w1288);
  FullAdder U382 (w1288, w1263, IN32[9], w1289, w1290);
  FullAdder U383 (w1290, w1265, IN33[8], w1291, w1292);
  FullAdder U384 (w1292, w1267, IN34[7], w1293, w1294);
  FullAdder U385 (w1294, w1269, IN35[6], w1295, w1296);
  FullAdder U386 (w1296, w1271, IN36[5], w1297, w1298);
  FullAdder U387 (w1298, w1273, IN37[4], w1299, w1300);
  FullAdder U388 (w1300, w1275, IN38[3], w1301, w1302);
  FullAdder U389 (w1302, w1277, IN39[2], w1303, w1304);
  FullAdder U390 (w1304, w1279, IN40[1], w1305, w1306);
  FullAdder U391 (w1306, w1280, IN41[0], w1307, w1308);
  HalfAdder U392 (w1283, IN29[13], Out1[29], w1310);
  FullAdder U393 (w1310, w1285, IN30[12], w1311, w1312);
  FullAdder U394 (w1312, w1287, IN31[11], w1313, w1314);
  FullAdder U395 (w1314, w1289, IN32[10], w1315, w1316);
  FullAdder U396 (w1316, w1291, IN33[9], w1317, w1318);
  FullAdder U397 (w1318, w1293, IN34[8], w1319, w1320);
  FullAdder U398 (w1320, w1295, IN35[7], w1321, w1322);
  FullAdder U399 (w1322, w1297, IN36[6], w1323, w1324);
  FullAdder U400 (w1324, w1299, IN37[5], w1325, w1326);
  FullAdder U401 (w1326, w1301, IN38[4], w1327, w1328);
  FullAdder U402 (w1328, w1303, IN39[3], w1329, w1330);
  FullAdder U403 (w1330, w1305, IN40[2], w1331, w1332);
  FullAdder U404 (w1332, w1307, IN41[1], w1333, w1334);
  FullAdder U405 (w1334, w1308, IN42[0], w1335, w1336);
  HalfAdder U406 (w1311, IN30[13], Out1[30], w1338);
  FullAdder U407 (w1338, w1313, IN31[12], w1339, w1340);
  FullAdder U408 (w1340, w1315, IN32[11], w1341, w1342);
  FullAdder U409 (w1342, w1317, IN33[10], w1343, w1344);
  FullAdder U410 (w1344, w1319, IN34[9], w1345, w1346);
  FullAdder U411 (w1346, w1321, IN35[8], w1347, w1348);
  FullAdder U412 (w1348, w1323, IN36[7], w1349, w1350);
  FullAdder U413 (w1350, w1325, IN37[6], w1351, w1352);
  FullAdder U414 (w1352, w1327, IN38[5], w1353, w1354);
  FullAdder U415 (w1354, w1329, IN39[4], w1355, w1356);
  FullAdder U416 (w1356, w1331, IN40[3], w1357, w1358);
  FullAdder U417 (w1358, w1333, IN41[2], w1359, w1360);
  FullAdder U418 (w1360, w1335, IN42[1], w1361, w1362);
  FullAdder U419 (w1362, w1336, IN43[0], w1363, w1364);
  HalfAdder U420 (w1339, IN31[13], Out1[31], w1366);
  FullAdder U421 (w1366, w1341, IN32[12], w1367, w1368);
  FullAdder U422 (w1368, w1343, IN33[11], w1369, w1370);
  FullAdder U423 (w1370, w1345, IN34[10], w1371, w1372);
  FullAdder U424 (w1372, w1347, IN35[9], w1373, w1374);
  FullAdder U425 (w1374, w1349, IN36[8], w1375, w1376);
  FullAdder U426 (w1376, w1351, IN37[7], w1377, w1378);
  FullAdder U427 (w1378, w1353, IN38[6], w1379, w1380);
  FullAdder U428 (w1380, w1355, IN39[5], w1381, w1382);
  FullAdder U429 (w1382, w1357, IN40[4], w1383, w1384);
  FullAdder U430 (w1384, w1359, IN41[3], w1385, w1386);
  FullAdder U431 (w1386, w1361, IN42[2], w1387, w1388);
  FullAdder U432 (w1388, w1363, IN43[1], w1389, w1390);
  FullAdder U433 (w1390, w1364, IN44[0], w1391, w1392);
  HalfAdder U434 (w1367, IN32[13], Out1[32], w1394);
  FullAdder U435 (w1394, w1369, IN33[12], w1395, w1396);
  FullAdder U436 (w1396, w1371, IN34[11], w1397, w1398);
  FullAdder U437 (w1398, w1373, IN35[10], w1399, w1400);
  FullAdder U438 (w1400, w1375, IN36[9], w1401, w1402);
  FullAdder U439 (w1402, w1377, IN37[8], w1403, w1404);
  FullAdder U440 (w1404, w1379, IN38[7], w1405, w1406);
  FullAdder U441 (w1406, w1381, IN39[6], w1407, w1408);
  FullAdder U442 (w1408, w1383, IN40[5], w1409, w1410);
  FullAdder U443 (w1410, w1385, IN41[4], w1411, w1412);
  FullAdder U444 (w1412, w1387, IN42[3], w1413, w1414);
  FullAdder U445 (w1414, w1389, IN43[2], w1415, w1416);
  FullAdder U446 (w1416, w1391, IN44[1], w1417, w1418);
  FullAdder U447 (w1418, w1392, IN45[0], w1419, w1420);
  HalfAdder U448 (w1395, IN33[13], Out1[33], w1422);
  FullAdder U449 (w1422, w1397, IN34[12], w1423, w1424);
  FullAdder U450 (w1424, w1399, IN35[11], w1425, w1426);
  FullAdder U451 (w1426, w1401, IN36[10], w1427, w1428);
  FullAdder U452 (w1428, w1403, IN37[9], w1429, w1430);
  FullAdder U453 (w1430, w1405, IN38[8], w1431, w1432);
  FullAdder U454 (w1432, w1407, IN39[7], w1433, w1434);
  FullAdder U455 (w1434, w1409, IN40[6], w1435, w1436);
  FullAdder U456 (w1436, w1411, IN41[5], w1437, w1438);
  FullAdder U457 (w1438, w1413, IN42[4], w1439, w1440);
  FullAdder U458 (w1440, w1415, IN43[3], w1441, w1442);
  FullAdder U459 (w1442, w1417, IN44[2], w1443, w1444);
  FullAdder U460 (w1444, w1419, IN45[1], w1445, w1446);
  FullAdder U461 (w1446, w1420, IN46[0], w1447, w1448);
  HalfAdder U462 (w1423, IN34[13], Out1[34], w1450);
  FullAdder U463 (w1450, w1425, IN35[12], Out1[35], w1452);
  FullAdder U464 (w1452, w1427, IN36[11], Out1[36], w1454);
  FullAdder U465 (w1454, w1429, IN37[10], Out1[37], w1456);
  FullAdder U466 (w1456, w1431, IN38[9], Out1[38], w1458);
  FullAdder U467 (w1458, w1433, IN39[8], Out1[39], w1460);
  FullAdder U468 (w1460, w1435, IN40[7], Out1[40], w1462);
  FullAdder U469 (w1462, w1437, IN41[6], Out1[41], w1464);
  FullAdder U470 (w1464, w1439, IN42[5], Out1[42], w1466);
  FullAdder U471 (w1466, w1441, IN43[4], Out1[43], w1468);
  FullAdder U472 (w1468, w1443, IN44[3], Out1[44], w1470);
  FullAdder U473 (w1470, w1445, IN45[2], Out1[45], w1472);
  FullAdder U474 (w1472, w1447, IN46[1], Out1[46], w1474);
  FullAdder U475 (w1474, w1448, IN47[0], Out1[47], Out1[48]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN15[14];
  assign Out2[1] = IN16[14];
  assign Out2[2] = IN17[14];
  assign Out2[3] = IN18[14];
  assign Out2[4] = IN19[14];
  assign Out2[5] = IN20[14];
  assign Out2[6] = IN21[14];
  assign Out2[7] = IN22[14];
  assign Out2[8] = IN23[14];
  assign Out2[9] = IN24[14];
  assign Out2[10] = IN25[14];
  assign Out2[11] = IN26[14];
  assign Out2[12] = IN27[14];
  assign Out2[13] = IN28[14];
  assign Out2[14] = IN29[14];
  assign Out2[15] = IN30[14];
  assign Out2[16] = IN31[14];
  assign Out2[17] = IN32[14];
  assign Out2[18] = IN33[14];
  assign Out2[19] = IN34[14];
  assign Out2[20] = IN35[13];
  assign Out2[21] = IN36[12];
  assign Out2[22] = IN37[11];
  assign Out2[23] = IN38[10];
  assign Out2[24] = IN39[9];
  assign Out2[25] = IN40[8];
  assign Out2[26] = IN41[7];
  assign Out2[27] = IN42[6];
  assign Out2[28] = IN43[5];
  assign Out2[29] = IN44[4];
  assign Out2[30] = IN45[3];
  assign Out2[31] = IN46[2];
  assign Out2[32] = IN47[1];
  assign Out2[33] = IN48[0];

endmodule
module RC_34_34(IN1, IN2, Out);
  input [33:0] IN1;
  input [33:0] IN2;
  output [34:0] Out;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w69);
  FullAdder U1 (IN1[1], IN2[1], w69, Out[1], w71);
  FullAdder U2 (IN1[2], IN2[2], w71, Out[2], w73);
  FullAdder U3 (IN1[3], IN2[3], w73, Out[3], w75);
  FullAdder U4 (IN1[4], IN2[4], w75, Out[4], w77);
  FullAdder U5 (IN1[5], IN2[5], w77, Out[5], w79);
  FullAdder U6 (IN1[6], IN2[6], w79, Out[6], w81);
  FullAdder U7 (IN1[7], IN2[7], w81, Out[7], w83);
  FullAdder U8 (IN1[8], IN2[8], w83, Out[8], w85);
  FullAdder U9 (IN1[9], IN2[9], w85, Out[9], w87);
  FullAdder U10 (IN1[10], IN2[10], w87, Out[10], w89);
  FullAdder U11 (IN1[11], IN2[11], w89, Out[11], w91);
  FullAdder U12 (IN1[12], IN2[12], w91, Out[12], w93);
  FullAdder U13 (IN1[13], IN2[13], w93, Out[13], w95);
  FullAdder U14 (IN1[14], IN2[14], w95, Out[14], w97);
  FullAdder U15 (IN1[15], IN2[15], w97, Out[15], w99);
  FullAdder U16 (IN1[16], IN2[16], w99, Out[16], w101);
  FullAdder U17 (IN1[17], IN2[17], w101, Out[17], w103);
  FullAdder U18 (IN1[18], IN2[18], w103, Out[18], w105);
  FullAdder U19 (IN1[19], IN2[19], w105, Out[19], w107);
  FullAdder U20 (IN1[20], IN2[20], w107, Out[20], w109);
  FullAdder U21 (IN1[21], IN2[21], w109, Out[21], w111);
  FullAdder U22 (IN1[22], IN2[22], w111, Out[22], w113);
  FullAdder U23 (IN1[23], IN2[23], w113, Out[23], w115);
  FullAdder U24 (IN1[24], IN2[24], w115, Out[24], w117);
  FullAdder U25 (IN1[25], IN2[25], w117, Out[25], w119);
  FullAdder U26 (IN1[26], IN2[26], w119, Out[26], w121);
  FullAdder U27 (IN1[27], IN2[27], w121, Out[27], w123);
  FullAdder U28 (IN1[28], IN2[28], w123, Out[28], w125);
  FullAdder U29 (IN1[29], IN2[29], w125, Out[29], w127);
  FullAdder U30 (IN1[30], IN2[30], w127, Out[30], w129);
  FullAdder U31 (IN1[31], IN2[31], w129, Out[31], w131);
  FullAdder U32 (IN1[32], IN2[32], w131, Out[32], w133);
  FullAdder U33 (IN1[33], IN2[33], w133, Out[33], Out[34]);

endmodule
module NR_15_35(IN1, IN2, Out);
  input [14:0] IN1;
  input [34:0] IN2;
  output [49:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [14:0] P15;
  wire [14:0] P16;
  wire [14:0] P17;
  wire [14:0] P18;
  wire [14:0] P19;
  wire [14:0] P20;
  wire [14:0] P21;
  wire [14:0] P22;
  wire [14:0] P23;
  wire [14:0] P24;
  wire [14:0] P25;
  wire [14:0] P26;
  wire [14:0] P27;
  wire [14:0] P28;
  wire [14:0] P29;
  wire [14:0] P30;
  wire [14:0] P31;
  wire [14:0] P32;
  wire [14:0] P33;
  wire [14:0] P34;
  wire [13:0] P35;
  wire [12:0] P36;
  wire [11:0] P37;
  wire [10:0] P38;
  wire [9:0] P39;
  wire [8:0] P40;
  wire [7:0] P41;
  wire [6:0] P42;
  wire [5:0] P43;
  wire [4:0] P44;
  wire [3:0] P45;
  wire [2:0] P46;
  wire [1:0] P47;
  wire [0:0] P48;
  wire [48:0] R1;
  wire [33:0] R2;
  wire [49:0] aOut;
  U_SP_15_35 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, R1, R2);
  RC_34_34 S2 (R1[48:15], R2, aOut[49:15]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign Out = aOut[49:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
