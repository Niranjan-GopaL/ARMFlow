//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 9
  second input length: 33
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_9_33(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40);
  input [8:0] IN1;
  input [32:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [8:0] P9;
  output [8:0] P10;
  output [8:0] P11;
  output [8:0] P12;
  output [8:0] P13;
  output [8:0] P14;
  output [8:0] P15;
  output [8:0] P16;
  output [8:0] P17;
  output [8:0] P18;
  output [8:0] P19;
  output [8:0] P20;
  output [8:0] P21;
  output [8:0] P22;
  output [8:0] P23;
  output [8:0] P24;
  output [8:0] P25;
  output [8:0] P26;
  output [8:0] P27;
  output [8:0] P28;
  output [8:0] P29;
  output [8:0] P30;
  output [8:0] P31;
  output [8:0] P32;
  output [7:0] P33;
  output [6:0] P34;
  output [5:0] P35;
  output [4:0] P36;
  output [3:0] P37;
  output [2:0] P38;
  output [1:0] P39;
  output [0:0] P40;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[0] = IN1[1]&IN2[32];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[1] = IN1[2]&IN2[31];
  assign P34[0] = IN1[2]&IN2[32];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[2] = IN1[3]&IN2[30];
  assign P34[1] = IN1[3]&IN2[31];
  assign P35[0] = IN1[3]&IN2[32];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[3] = IN1[4]&IN2[29];
  assign P34[2] = IN1[4]&IN2[30];
  assign P35[1] = IN1[4]&IN2[31];
  assign P36[0] = IN1[4]&IN2[32];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[4] = IN1[5]&IN2[28];
  assign P34[3] = IN1[5]&IN2[29];
  assign P35[2] = IN1[5]&IN2[30];
  assign P36[1] = IN1[5]&IN2[31];
  assign P37[0] = IN1[5]&IN2[32];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[5] = IN1[6]&IN2[27];
  assign P34[4] = IN1[6]&IN2[28];
  assign P35[3] = IN1[6]&IN2[29];
  assign P36[2] = IN1[6]&IN2[30];
  assign P37[1] = IN1[6]&IN2[31];
  assign P38[0] = IN1[6]&IN2[32];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[6] = IN1[7]&IN2[26];
  assign P34[5] = IN1[7]&IN2[27];
  assign P35[4] = IN1[7]&IN2[28];
  assign P36[3] = IN1[7]&IN2[29];
  assign P37[2] = IN1[7]&IN2[30];
  assign P38[1] = IN1[7]&IN2[31];
  assign P39[0] = IN1[7]&IN2[32];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[7] = IN1[8]&IN2[25];
  assign P34[6] = IN1[8]&IN2[26];
  assign P35[5] = IN1[8]&IN2[27];
  assign P36[4] = IN1[8]&IN2[28];
  assign P37[3] = IN1[8]&IN2[29];
  assign P38[2] = IN1[8]&IN2[30];
  assign P39[1] = IN1[8]&IN2[31];
  assign P40[0] = IN1[8]&IN2[32];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [8:0] IN9;
  input [8:0] IN10;
  input [8:0] IN11;
  input [8:0] IN12;
  input [8:0] IN13;
  input [8:0] IN14;
  input [8:0] IN15;
  input [8:0] IN16;
  input [8:0] IN17;
  input [8:0] IN18;
  input [8:0] IN19;
  input [8:0] IN20;
  input [8:0] IN21;
  input [8:0] IN22;
  input [8:0] IN23;
  input [8:0] IN24;
  input [8:0] IN25;
  input [8:0] IN26;
  input [8:0] IN27;
  input [8:0] IN28;
  input [8:0] IN29;
  input [8:0] IN30;
  input [8:0] IN31;
  input [8:0] IN32;
  input [7:0] IN33;
  input [6:0] IN34;
  input [5:0] IN35;
  input [4:0] IN36;
  input [3:0] IN37;
  input [2:0] IN38;
  input [1:0] IN39;
  input [0:0] IN40;
  output [40:0] Out1;
  output [31:0] Out2;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w794;
  wire w796;
  wire w798;
  wire w800;
  wire w802;
  wire w804;
  wire w806;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w298);
  FullAdder U1 (w298, IN2[0], IN2[1], w299, w300);
  FullAdder U2 (w300, IN3[0], IN3[1], w301, w302);
  FullAdder U3 (w302, IN4[0], IN4[1], w303, w304);
  FullAdder U4 (w304, IN5[0], IN5[1], w305, w306);
  FullAdder U5 (w306, IN6[0], IN6[1], w307, w308);
  FullAdder U6 (w308, IN7[0], IN7[1], w309, w310);
  FullAdder U7 (w310, IN8[0], IN8[1], w311, w312);
  HalfAdder U8 (w299, IN2[2], Out1[2], w314);
  FullAdder U9 (w314, w301, IN3[2], w315, w316);
  FullAdder U10 (w316, w303, IN4[2], w317, w318);
  FullAdder U11 (w318, w305, IN5[2], w319, w320);
  FullAdder U12 (w320, w307, IN6[2], w321, w322);
  FullAdder U13 (w322, w309, IN7[2], w323, w324);
  FullAdder U14 (w324, w311, IN8[2], w325, w326);
  FullAdder U15 (w326, w312, IN9[0], w327, w328);
  HalfAdder U16 (w315, IN3[3], Out1[3], w330);
  FullAdder U17 (w330, w317, IN4[3], w331, w332);
  FullAdder U18 (w332, w319, IN5[3], w333, w334);
  FullAdder U19 (w334, w321, IN6[3], w335, w336);
  FullAdder U20 (w336, w323, IN7[3], w337, w338);
  FullAdder U21 (w338, w325, IN8[3], w339, w340);
  FullAdder U22 (w340, w327, IN9[1], w341, w342);
  FullAdder U23 (w342, w328, IN10[0], w343, w344);
  HalfAdder U24 (w331, IN4[4], Out1[4], w346);
  FullAdder U25 (w346, w333, IN5[4], w347, w348);
  FullAdder U26 (w348, w335, IN6[4], w349, w350);
  FullAdder U27 (w350, w337, IN7[4], w351, w352);
  FullAdder U28 (w352, w339, IN8[4], w353, w354);
  FullAdder U29 (w354, w341, IN9[2], w355, w356);
  FullAdder U30 (w356, w343, IN10[1], w357, w358);
  FullAdder U31 (w358, w344, IN11[0], w359, w360);
  HalfAdder U32 (w347, IN5[5], Out1[5], w362);
  FullAdder U33 (w362, w349, IN6[5], w363, w364);
  FullAdder U34 (w364, w351, IN7[5], w365, w366);
  FullAdder U35 (w366, w353, IN8[5], w367, w368);
  FullAdder U36 (w368, w355, IN9[3], w369, w370);
  FullAdder U37 (w370, w357, IN10[2], w371, w372);
  FullAdder U38 (w372, w359, IN11[1], w373, w374);
  FullAdder U39 (w374, w360, IN12[0], w375, w376);
  HalfAdder U40 (w363, IN6[6], Out1[6], w378);
  FullAdder U41 (w378, w365, IN7[6], w379, w380);
  FullAdder U42 (w380, w367, IN8[6], w381, w382);
  FullAdder U43 (w382, w369, IN9[4], w383, w384);
  FullAdder U44 (w384, w371, IN10[3], w385, w386);
  FullAdder U45 (w386, w373, IN11[2], w387, w388);
  FullAdder U46 (w388, w375, IN12[1], w389, w390);
  FullAdder U47 (w390, w376, IN13[0], w391, w392);
  HalfAdder U48 (w379, IN7[7], Out1[7], w394);
  FullAdder U49 (w394, w381, IN8[7], w395, w396);
  FullAdder U50 (w396, w383, IN9[5], w397, w398);
  FullAdder U51 (w398, w385, IN10[4], w399, w400);
  FullAdder U52 (w400, w387, IN11[3], w401, w402);
  FullAdder U53 (w402, w389, IN12[2], w403, w404);
  FullAdder U54 (w404, w391, IN13[1], w405, w406);
  FullAdder U55 (w406, w392, IN14[0], w407, w408);
  HalfAdder U56 (w395, IN8[8], Out1[8], w410);
  FullAdder U57 (w410, w397, IN9[6], w411, w412);
  FullAdder U58 (w412, w399, IN10[5], w413, w414);
  FullAdder U59 (w414, w401, IN11[4], w415, w416);
  FullAdder U60 (w416, w403, IN12[3], w417, w418);
  FullAdder U61 (w418, w405, IN13[2], w419, w420);
  FullAdder U62 (w420, w407, IN14[1], w421, w422);
  FullAdder U63 (w422, w408, IN15[0], w423, w424);
  HalfAdder U64 (w411, IN9[7], Out1[9], w426);
  FullAdder U65 (w426, w413, IN10[6], w427, w428);
  FullAdder U66 (w428, w415, IN11[5], w429, w430);
  FullAdder U67 (w430, w417, IN12[4], w431, w432);
  FullAdder U68 (w432, w419, IN13[3], w433, w434);
  FullAdder U69 (w434, w421, IN14[2], w435, w436);
  FullAdder U70 (w436, w423, IN15[1], w437, w438);
  FullAdder U71 (w438, w424, IN16[0], w439, w440);
  HalfAdder U72 (w427, IN10[7], Out1[10], w442);
  FullAdder U73 (w442, w429, IN11[6], w443, w444);
  FullAdder U74 (w444, w431, IN12[5], w445, w446);
  FullAdder U75 (w446, w433, IN13[4], w447, w448);
  FullAdder U76 (w448, w435, IN14[3], w449, w450);
  FullAdder U77 (w450, w437, IN15[2], w451, w452);
  FullAdder U78 (w452, w439, IN16[1], w453, w454);
  FullAdder U79 (w454, w440, IN17[0], w455, w456);
  HalfAdder U80 (w443, IN11[7], Out1[11], w458);
  FullAdder U81 (w458, w445, IN12[6], w459, w460);
  FullAdder U82 (w460, w447, IN13[5], w461, w462);
  FullAdder U83 (w462, w449, IN14[4], w463, w464);
  FullAdder U84 (w464, w451, IN15[3], w465, w466);
  FullAdder U85 (w466, w453, IN16[2], w467, w468);
  FullAdder U86 (w468, w455, IN17[1], w469, w470);
  FullAdder U87 (w470, w456, IN18[0], w471, w472);
  HalfAdder U88 (w459, IN12[7], Out1[12], w474);
  FullAdder U89 (w474, w461, IN13[6], w475, w476);
  FullAdder U90 (w476, w463, IN14[5], w477, w478);
  FullAdder U91 (w478, w465, IN15[4], w479, w480);
  FullAdder U92 (w480, w467, IN16[3], w481, w482);
  FullAdder U93 (w482, w469, IN17[2], w483, w484);
  FullAdder U94 (w484, w471, IN18[1], w485, w486);
  FullAdder U95 (w486, w472, IN19[0], w487, w488);
  HalfAdder U96 (w475, IN13[7], Out1[13], w490);
  FullAdder U97 (w490, w477, IN14[6], w491, w492);
  FullAdder U98 (w492, w479, IN15[5], w493, w494);
  FullAdder U99 (w494, w481, IN16[4], w495, w496);
  FullAdder U100 (w496, w483, IN17[3], w497, w498);
  FullAdder U101 (w498, w485, IN18[2], w499, w500);
  FullAdder U102 (w500, w487, IN19[1], w501, w502);
  FullAdder U103 (w502, w488, IN20[0], w503, w504);
  HalfAdder U104 (w491, IN14[7], Out1[14], w506);
  FullAdder U105 (w506, w493, IN15[6], w507, w508);
  FullAdder U106 (w508, w495, IN16[5], w509, w510);
  FullAdder U107 (w510, w497, IN17[4], w511, w512);
  FullAdder U108 (w512, w499, IN18[3], w513, w514);
  FullAdder U109 (w514, w501, IN19[2], w515, w516);
  FullAdder U110 (w516, w503, IN20[1], w517, w518);
  FullAdder U111 (w518, w504, IN21[0], w519, w520);
  HalfAdder U112 (w507, IN15[7], Out1[15], w522);
  FullAdder U113 (w522, w509, IN16[6], w523, w524);
  FullAdder U114 (w524, w511, IN17[5], w525, w526);
  FullAdder U115 (w526, w513, IN18[4], w527, w528);
  FullAdder U116 (w528, w515, IN19[3], w529, w530);
  FullAdder U117 (w530, w517, IN20[2], w531, w532);
  FullAdder U118 (w532, w519, IN21[1], w533, w534);
  FullAdder U119 (w534, w520, IN22[0], w535, w536);
  HalfAdder U120 (w523, IN16[7], Out1[16], w538);
  FullAdder U121 (w538, w525, IN17[6], w539, w540);
  FullAdder U122 (w540, w527, IN18[5], w541, w542);
  FullAdder U123 (w542, w529, IN19[4], w543, w544);
  FullAdder U124 (w544, w531, IN20[3], w545, w546);
  FullAdder U125 (w546, w533, IN21[2], w547, w548);
  FullAdder U126 (w548, w535, IN22[1], w549, w550);
  FullAdder U127 (w550, w536, IN23[0], w551, w552);
  HalfAdder U128 (w539, IN17[7], Out1[17], w554);
  FullAdder U129 (w554, w541, IN18[6], w555, w556);
  FullAdder U130 (w556, w543, IN19[5], w557, w558);
  FullAdder U131 (w558, w545, IN20[4], w559, w560);
  FullAdder U132 (w560, w547, IN21[3], w561, w562);
  FullAdder U133 (w562, w549, IN22[2], w563, w564);
  FullAdder U134 (w564, w551, IN23[1], w565, w566);
  FullAdder U135 (w566, w552, IN24[0], w567, w568);
  HalfAdder U136 (w555, IN18[7], Out1[18], w570);
  FullAdder U137 (w570, w557, IN19[6], w571, w572);
  FullAdder U138 (w572, w559, IN20[5], w573, w574);
  FullAdder U139 (w574, w561, IN21[4], w575, w576);
  FullAdder U140 (w576, w563, IN22[3], w577, w578);
  FullAdder U141 (w578, w565, IN23[2], w579, w580);
  FullAdder U142 (w580, w567, IN24[1], w581, w582);
  FullAdder U143 (w582, w568, IN25[0], w583, w584);
  HalfAdder U144 (w571, IN19[7], Out1[19], w586);
  FullAdder U145 (w586, w573, IN20[6], w587, w588);
  FullAdder U146 (w588, w575, IN21[5], w589, w590);
  FullAdder U147 (w590, w577, IN22[4], w591, w592);
  FullAdder U148 (w592, w579, IN23[3], w593, w594);
  FullAdder U149 (w594, w581, IN24[2], w595, w596);
  FullAdder U150 (w596, w583, IN25[1], w597, w598);
  FullAdder U151 (w598, w584, IN26[0], w599, w600);
  HalfAdder U152 (w587, IN20[7], Out1[20], w602);
  FullAdder U153 (w602, w589, IN21[6], w603, w604);
  FullAdder U154 (w604, w591, IN22[5], w605, w606);
  FullAdder U155 (w606, w593, IN23[4], w607, w608);
  FullAdder U156 (w608, w595, IN24[3], w609, w610);
  FullAdder U157 (w610, w597, IN25[2], w611, w612);
  FullAdder U158 (w612, w599, IN26[1], w613, w614);
  FullAdder U159 (w614, w600, IN27[0], w615, w616);
  HalfAdder U160 (w603, IN21[7], Out1[21], w618);
  FullAdder U161 (w618, w605, IN22[6], w619, w620);
  FullAdder U162 (w620, w607, IN23[5], w621, w622);
  FullAdder U163 (w622, w609, IN24[4], w623, w624);
  FullAdder U164 (w624, w611, IN25[3], w625, w626);
  FullAdder U165 (w626, w613, IN26[2], w627, w628);
  FullAdder U166 (w628, w615, IN27[1], w629, w630);
  FullAdder U167 (w630, w616, IN28[0], w631, w632);
  HalfAdder U168 (w619, IN22[7], Out1[22], w634);
  FullAdder U169 (w634, w621, IN23[6], w635, w636);
  FullAdder U170 (w636, w623, IN24[5], w637, w638);
  FullAdder U171 (w638, w625, IN25[4], w639, w640);
  FullAdder U172 (w640, w627, IN26[3], w641, w642);
  FullAdder U173 (w642, w629, IN27[2], w643, w644);
  FullAdder U174 (w644, w631, IN28[1], w645, w646);
  FullAdder U175 (w646, w632, IN29[0], w647, w648);
  HalfAdder U176 (w635, IN23[7], Out1[23], w650);
  FullAdder U177 (w650, w637, IN24[6], w651, w652);
  FullAdder U178 (w652, w639, IN25[5], w653, w654);
  FullAdder U179 (w654, w641, IN26[4], w655, w656);
  FullAdder U180 (w656, w643, IN27[3], w657, w658);
  FullAdder U181 (w658, w645, IN28[2], w659, w660);
  FullAdder U182 (w660, w647, IN29[1], w661, w662);
  FullAdder U183 (w662, w648, IN30[0], w663, w664);
  HalfAdder U184 (w651, IN24[7], Out1[24], w666);
  FullAdder U185 (w666, w653, IN25[6], w667, w668);
  FullAdder U186 (w668, w655, IN26[5], w669, w670);
  FullAdder U187 (w670, w657, IN27[4], w671, w672);
  FullAdder U188 (w672, w659, IN28[3], w673, w674);
  FullAdder U189 (w674, w661, IN29[2], w675, w676);
  FullAdder U190 (w676, w663, IN30[1], w677, w678);
  FullAdder U191 (w678, w664, IN31[0], w679, w680);
  HalfAdder U192 (w667, IN25[7], Out1[25], w682);
  FullAdder U193 (w682, w669, IN26[6], w683, w684);
  FullAdder U194 (w684, w671, IN27[5], w685, w686);
  FullAdder U195 (w686, w673, IN28[4], w687, w688);
  FullAdder U196 (w688, w675, IN29[3], w689, w690);
  FullAdder U197 (w690, w677, IN30[2], w691, w692);
  FullAdder U198 (w692, w679, IN31[1], w693, w694);
  FullAdder U199 (w694, w680, IN32[0], w695, w696);
  HalfAdder U200 (w683, IN26[7], Out1[26], w698);
  FullAdder U201 (w698, w685, IN27[6], w699, w700);
  FullAdder U202 (w700, w687, IN28[5], w701, w702);
  FullAdder U203 (w702, w689, IN29[4], w703, w704);
  FullAdder U204 (w704, w691, IN30[3], w705, w706);
  FullAdder U205 (w706, w693, IN31[2], w707, w708);
  FullAdder U206 (w708, w695, IN32[1], w709, w710);
  FullAdder U207 (w710, w696, IN33[0], w711, w712);
  HalfAdder U208 (w699, IN27[7], Out1[27], w714);
  FullAdder U209 (w714, w701, IN28[6], w715, w716);
  FullAdder U210 (w716, w703, IN29[5], w717, w718);
  FullAdder U211 (w718, w705, IN30[4], w719, w720);
  FullAdder U212 (w720, w707, IN31[3], w721, w722);
  FullAdder U213 (w722, w709, IN32[2], w723, w724);
  FullAdder U214 (w724, w711, IN33[1], w725, w726);
  FullAdder U215 (w726, w712, IN34[0], w727, w728);
  HalfAdder U216 (w715, IN28[7], Out1[28], w730);
  FullAdder U217 (w730, w717, IN29[6], w731, w732);
  FullAdder U218 (w732, w719, IN30[5], w733, w734);
  FullAdder U219 (w734, w721, IN31[4], w735, w736);
  FullAdder U220 (w736, w723, IN32[3], w737, w738);
  FullAdder U221 (w738, w725, IN33[2], w739, w740);
  FullAdder U222 (w740, w727, IN34[1], w741, w742);
  FullAdder U223 (w742, w728, IN35[0], w743, w744);
  HalfAdder U224 (w731, IN29[7], Out1[29], w746);
  FullAdder U225 (w746, w733, IN30[6], w747, w748);
  FullAdder U226 (w748, w735, IN31[5], w749, w750);
  FullAdder U227 (w750, w737, IN32[4], w751, w752);
  FullAdder U228 (w752, w739, IN33[3], w753, w754);
  FullAdder U229 (w754, w741, IN34[2], w755, w756);
  FullAdder U230 (w756, w743, IN35[1], w757, w758);
  FullAdder U231 (w758, w744, IN36[0], w759, w760);
  HalfAdder U232 (w747, IN30[7], Out1[30], w762);
  FullAdder U233 (w762, w749, IN31[6], w763, w764);
  FullAdder U234 (w764, w751, IN32[5], w765, w766);
  FullAdder U235 (w766, w753, IN33[4], w767, w768);
  FullAdder U236 (w768, w755, IN34[3], w769, w770);
  FullAdder U237 (w770, w757, IN35[2], w771, w772);
  FullAdder U238 (w772, w759, IN36[1], w773, w774);
  FullAdder U239 (w774, w760, IN37[0], w775, w776);
  HalfAdder U240 (w763, IN31[7], Out1[31], w778);
  FullAdder U241 (w778, w765, IN32[6], w779, w780);
  FullAdder U242 (w780, w767, IN33[5], w781, w782);
  FullAdder U243 (w782, w769, IN34[4], w783, w784);
  FullAdder U244 (w784, w771, IN35[3], w785, w786);
  FullAdder U245 (w786, w773, IN36[2], w787, w788);
  FullAdder U246 (w788, w775, IN37[1], w789, w790);
  FullAdder U247 (w790, w776, IN38[0], w791, w792);
  HalfAdder U248 (w779, IN32[7], Out1[32], w794);
  FullAdder U249 (w794, w781, IN33[6], Out1[33], w796);
  FullAdder U250 (w796, w783, IN34[5], Out1[34], w798);
  FullAdder U251 (w798, w785, IN35[4], Out1[35], w800);
  FullAdder U252 (w800, w787, IN36[3], Out1[36], w802);
  FullAdder U253 (w802, w789, IN37[2], Out1[37], w804);
  FullAdder U254 (w804, w791, IN38[1], Out1[38], w806);
  FullAdder U255 (w806, w792, IN39[0], Out1[39], Out1[40]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN9[8];
  assign Out2[1] = IN10[8];
  assign Out2[2] = IN11[8];
  assign Out2[3] = IN12[8];
  assign Out2[4] = IN13[8];
  assign Out2[5] = IN14[8];
  assign Out2[6] = IN15[8];
  assign Out2[7] = IN16[8];
  assign Out2[8] = IN17[8];
  assign Out2[9] = IN18[8];
  assign Out2[10] = IN19[8];
  assign Out2[11] = IN20[8];
  assign Out2[12] = IN21[8];
  assign Out2[13] = IN22[8];
  assign Out2[14] = IN23[8];
  assign Out2[15] = IN24[8];
  assign Out2[16] = IN25[8];
  assign Out2[17] = IN26[8];
  assign Out2[18] = IN27[8];
  assign Out2[19] = IN28[8];
  assign Out2[20] = IN29[8];
  assign Out2[21] = IN30[8];
  assign Out2[22] = IN31[8];
  assign Out2[23] = IN32[8];
  assign Out2[24] = IN33[7];
  assign Out2[25] = IN34[6];
  assign Out2[26] = IN35[5];
  assign Out2[27] = IN36[4];
  assign Out2[28] = IN37[3];
  assign Out2[29] = IN38[2];
  assign Out2[30] = IN39[1];
  assign Out2[31] = IN40[0];

endmodule
module RC_32_32(IN1, IN2, Out);
  input [31:0] IN1;
  input [31:0] IN2;
  output [32:0] Out;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w65);
  FullAdder U1 (IN1[1], IN2[1], w65, Out[1], w67);
  FullAdder U2 (IN1[2], IN2[2], w67, Out[2], w69);
  FullAdder U3 (IN1[3], IN2[3], w69, Out[3], w71);
  FullAdder U4 (IN1[4], IN2[4], w71, Out[4], w73);
  FullAdder U5 (IN1[5], IN2[5], w73, Out[5], w75);
  FullAdder U6 (IN1[6], IN2[6], w75, Out[6], w77);
  FullAdder U7 (IN1[7], IN2[7], w77, Out[7], w79);
  FullAdder U8 (IN1[8], IN2[8], w79, Out[8], w81);
  FullAdder U9 (IN1[9], IN2[9], w81, Out[9], w83);
  FullAdder U10 (IN1[10], IN2[10], w83, Out[10], w85);
  FullAdder U11 (IN1[11], IN2[11], w85, Out[11], w87);
  FullAdder U12 (IN1[12], IN2[12], w87, Out[12], w89);
  FullAdder U13 (IN1[13], IN2[13], w89, Out[13], w91);
  FullAdder U14 (IN1[14], IN2[14], w91, Out[14], w93);
  FullAdder U15 (IN1[15], IN2[15], w93, Out[15], w95);
  FullAdder U16 (IN1[16], IN2[16], w95, Out[16], w97);
  FullAdder U17 (IN1[17], IN2[17], w97, Out[17], w99);
  FullAdder U18 (IN1[18], IN2[18], w99, Out[18], w101);
  FullAdder U19 (IN1[19], IN2[19], w101, Out[19], w103);
  FullAdder U20 (IN1[20], IN2[20], w103, Out[20], w105);
  FullAdder U21 (IN1[21], IN2[21], w105, Out[21], w107);
  FullAdder U22 (IN1[22], IN2[22], w107, Out[22], w109);
  FullAdder U23 (IN1[23], IN2[23], w109, Out[23], w111);
  FullAdder U24 (IN1[24], IN2[24], w111, Out[24], w113);
  FullAdder U25 (IN1[25], IN2[25], w113, Out[25], w115);
  FullAdder U26 (IN1[26], IN2[26], w115, Out[26], w117);
  FullAdder U27 (IN1[27], IN2[27], w117, Out[27], w119);
  FullAdder U28 (IN1[28], IN2[28], w119, Out[28], w121);
  FullAdder U29 (IN1[29], IN2[29], w121, Out[29], w123);
  FullAdder U30 (IN1[30], IN2[30], w123, Out[30], w125);
  FullAdder U31 (IN1[31], IN2[31], w125, Out[31], Out[32]);

endmodule
module NR_9_33(IN1, IN2, Out);
  input [8:0] IN1;
  input [32:0] IN2;
  output [41:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [8:0] P9;
  wire [8:0] P10;
  wire [8:0] P11;
  wire [8:0] P12;
  wire [8:0] P13;
  wire [8:0] P14;
  wire [8:0] P15;
  wire [8:0] P16;
  wire [8:0] P17;
  wire [8:0] P18;
  wire [8:0] P19;
  wire [8:0] P20;
  wire [8:0] P21;
  wire [8:0] P22;
  wire [8:0] P23;
  wire [8:0] P24;
  wire [8:0] P25;
  wire [8:0] P26;
  wire [8:0] P27;
  wire [8:0] P28;
  wire [8:0] P29;
  wire [8:0] P30;
  wire [8:0] P31;
  wire [8:0] P32;
  wire [7:0] P33;
  wire [6:0] P34;
  wire [5:0] P35;
  wire [4:0] P36;
  wire [3:0] P37;
  wire [2:0] P38;
  wire [1:0] P39;
  wire [0:0] P40;
  wire [40:0] R1;
  wire [31:0] R2;
  wire [41:0] aOut;
  U_SP_9_33 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, R1, R2);
  RC_32_32 S2 (R1[40:9], R2, aOut[41:9]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign Out = aOut[41:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
