
module customAdder53_0(
    input [52 : 0] A,
    input [52 : 0] B,
    output [53 : 0] Sum
);

    assign Sum = A+B;

endmodule
