
module NR_54_1(
    input [53:0]IN1,
    input [0:0]IN2,
    output [53:0]Out
);
    assign Out = IN2;
endmodule
