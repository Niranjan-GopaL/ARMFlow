
module customAdder45_0(
    input [44 : 0] A,
    input [44 : 0] B,
    output [45 : 0] Sum
);

    assign Sum = A+B;

endmodule
