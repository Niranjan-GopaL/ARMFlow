//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 5
  second input length: 40
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_5_40(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43);
  input [4:0] IN1;
  input [39:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [4:0] P5;
  output [4:0] P6;
  output [4:0] P7;
  output [4:0] P8;
  output [4:0] P9;
  output [4:0] P10;
  output [4:0] P11;
  output [4:0] P12;
  output [4:0] P13;
  output [4:0] P14;
  output [4:0] P15;
  output [4:0] P16;
  output [4:0] P17;
  output [4:0] P18;
  output [4:0] P19;
  output [4:0] P20;
  output [4:0] P21;
  output [4:0] P22;
  output [4:0] P23;
  output [4:0] P24;
  output [4:0] P25;
  output [4:0] P26;
  output [4:0] P27;
  output [4:0] P28;
  output [4:0] P29;
  output [4:0] P30;
  output [4:0] P31;
  output [4:0] P32;
  output [4:0] P33;
  output [4:0] P34;
  output [4:0] P35;
  output [4:0] P36;
  output [4:0] P37;
  output [4:0] P38;
  output [4:0] P39;
  output [3:0] P40;
  output [2:0] P41;
  output [1:0] P42;
  output [0:0] P43;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[0] = IN1[1]&IN2[39];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[1] = IN1[2]&IN2[38];
  assign P41[0] = IN1[2]&IN2[39];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[2] = IN1[3]&IN2[37];
  assign P41[1] = IN1[3]&IN2[38];
  assign P42[0] = IN1[3]&IN2[39];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[3] = IN1[4]&IN2[36];
  assign P41[2] = IN1[4]&IN2[37];
  assign P42[1] = IN1[4]&IN2[38];
  assign P43[0] = IN1[4]&IN2[39];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [4:0] IN5;
  input [4:0] IN6;
  input [4:0] IN7;
  input [4:0] IN8;
  input [4:0] IN9;
  input [4:0] IN10;
  input [4:0] IN11;
  input [4:0] IN12;
  input [4:0] IN13;
  input [4:0] IN14;
  input [4:0] IN15;
  input [4:0] IN16;
  input [4:0] IN17;
  input [4:0] IN18;
  input [4:0] IN19;
  input [4:0] IN20;
  input [4:0] IN21;
  input [4:0] IN22;
  input [4:0] IN23;
  input [4:0] IN24;
  input [4:0] IN25;
  input [4:0] IN26;
  input [4:0] IN27;
  input [4:0] IN28;
  input [4:0] IN29;
  input [4:0] IN30;
  input [4:0] IN31;
  input [4:0] IN32;
  input [4:0] IN33;
  input [4:0] IN34;
  input [4:0] IN35;
  input [4:0] IN36;
  input [4:0] IN37;
  input [4:0] IN38;
  input [4:0] IN39;
  input [3:0] IN40;
  input [2:0] IN41;
  input [1:0] IN42;
  input [0:0] IN43;
  output [43:0] Out1;
  output [38:0] Out2;
  wire w201;
  wire w202;
  wire w203;
  wire w204;
  wire w205;
  wire w206;
  wire w207;
  wire w209;
  wire w210;
  wire w211;
  wire w212;
  wire w213;
  wire w214;
  wire w215;
  wire w217;
  wire w218;
  wire w219;
  wire w220;
  wire w221;
  wire w222;
  wire w223;
  wire w225;
  wire w226;
  wire w227;
  wire w228;
  wire w229;
  wire w230;
  wire w231;
  wire w233;
  wire w234;
  wire w235;
  wire w236;
  wire w237;
  wire w238;
  wire w239;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w246;
  wire w247;
  wire w249;
  wire w250;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w505;
  wire w507;
  wire w509;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w201);
  FullAdder U1 (w201, IN2[0], IN2[1], w202, w203);
  FullAdder U2 (w203, IN3[0], IN3[1], w204, w205);
  FullAdder U3 (w205, IN4[0], IN4[1], w206, w207);
  HalfAdder U4 (w202, IN2[2], Out1[2], w209);
  FullAdder U5 (w209, w204, IN3[2], w210, w211);
  FullAdder U6 (w211, w206, IN4[2], w212, w213);
  FullAdder U7 (w213, w207, IN5[0], w214, w215);
  HalfAdder U8 (w210, IN3[3], Out1[3], w217);
  FullAdder U9 (w217, w212, IN4[3], w218, w219);
  FullAdder U10 (w219, w214, IN5[1], w220, w221);
  FullAdder U11 (w221, w215, IN6[0], w222, w223);
  HalfAdder U12 (w218, IN4[4], Out1[4], w225);
  FullAdder U13 (w225, w220, IN5[2], w226, w227);
  FullAdder U14 (w227, w222, IN6[1], w228, w229);
  FullAdder U15 (w229, w223, IN7[0], w230, w231);
  HalfAdder U16 (w226, IN5[3], Out1[5], w233);
  FullAdder U17 (w233, w228, IN6[2], w234, w235);
  FullAdder U18 (w235, w230, IN7[1], w236, w237);
  FullAdder U19 (w237, w231, IN8[0], w238, w239);
  HalfAdder U20 (w234, IN6[3], Out1[6], w241);
  FullAdder U21 (w241, w236, IN7[2], w242, w243);
  FullAdder U22 (w243, w238, IN8[1], w244, w245);
  FullAdder U23 (w245, w239, IN9[0], w246, w247);
  HalfAdder U24 (w242, IN7[3], Out1[7], w249);
  FullAdder U25 (w249, w244, IN8[2], w250, w251);
  FullAdder U26 (w251, w246, IN9[1], w252, w253);
  FullAdder U27 (w253, w247, IN10[0], w254, w255);
  HalfAdder U28 (w250, IN8[3], Out1[8], w257);
  FullAdder U29 (w257, w252, IN9[2], w258, w259);
  FullAdder U30 (w259, w254, IN10[1], w260, w261);
  FullAdder U31 (w261, w255, IN11[0], w262, w263);
  HalfAdder U32 (w258, IN9[3], Out1[9], w265);
  FullAdder U33 (w265, w260, IN10[2], w266, w267);
  FullAdder U34 (w267, w262, IN11[1], w268, w269);
  FullAdder U35 (w269, w263, IN12[0], w270, w271);
  HalfAdder U36 (w266, IN10[3], Out1[10], w273);
  FullAdder U37 (w273, w268, IN11[2], w274, w275);
  FullAdder U38 (w275, w270, IN12[1], w276, w277);
  FullAdder U39 (w277, w271, IN13[0], w278, w279);
  HalfAdder U40 (w274, IN11[3], Out1[11], w281);
  FullAdder U41 (w281, w276, IN12[2], w282, w283);
  FullAdder U42 (w283, w278, IN13[1], w284, w285);
  FullAdder U43 (w285, w279, IN14[0], w286, w287);
  HalfAdder U44 (w282, IN12[3], Out1[12], w289);
  FullAdder U45 (w289, w284, IN13[2], w290, w291);
  FullAdder U46 (w291, w286, IN14[1], w292, w293);
  FullAdder U47 (w293, w287, IN15[0], w294, w295);
  HalfAdder U48 (w290, IN13[3], Out1[13], w297);
  FullAdder U49 (w297, w292, IN14[2], w298, w299);
  FullAdder U50 (w299, w294, IN15[1], w300, w301);
  FullAdder U51 (w301, w295, IN16[0], w302, w303);
  HalfAdder U52 (w298, IN14[3], Out1[14], w305);
  FullAdder U53 (w305, w300, IN15[2], w306, w307);
  FullAdder U54 (w307, w302, IN16[1], w308, w309);
  FullAdder U55 (w309, w303, IN17[0], w310, w311);
  HalfAdder U56 (w306, IN15[3], Out1[15], w313);
  FullAdder U57 (w313, w308, IN16[2], w314, w315);
  FullAdder U58 (w315, w310, IN17[1], w316, w317);
  FullAdder U59 (w317, w311, IN18[0], w318, w319);
  HalfAdder U60 (w314, IN16[3], Out1[16], w321);
  FullAdder U61 (w321, w316, IN17[2], w322, w323);
  FullAdder U62 (w323, w318, IN18[1], w324, w325);
  FullAdder U63 (w325, w319, IN19[0], w326, w327);
  HalfAdder U64 (w322, IN17[3], Out1[17], w329);
  FullAdder U65 (w329, w324, IN18[2], w330, w331);
  FullAdder U66 (w331, w326, IN19[1], w332, w333);
  FullAdder U67 (w333, w327, IN20[0], w334, w335);
  HalfAdder U68 (w330, IN18[3], Out1[18], w337);
  FullAdder U69 (w337, w332, IN19[2], w338, w339);
  FullAdder U70 (w339, w334, IN20[1], w340, w341);
  FullAdder U71 (w341, w335, IN21[0], w342, w343);
  HalfAdder U72 (w338, IN19[3], Out1[19], w345);
  FullAdder U73 (w345, w340, IN20[2], w346, w347);
  FullAdder U74 (w347, w342, IN21[1], w348, w349);
  FullAdder U75 (w349, w343, IN22[0], w350, w351);
  HalfAdder U76 (w346, IN20[3], Out1[20], w353);
  FullAdder U77 (w353, w348, IN21[2], w354, w355);
  FullAdder U78 (w355, w350, IN22[1], w356, w357);
  FullAdder U79 (w357, w351, IN23[0], w358, w359);
  HalfAdder U80 (w354, IN21[3], Out1[21], w361);
  FullAdder U81 (w361, w356, IN22[2], w362, w363);
  FullAdder U82 (w363, w358, IN23[1], w364, w365);
  FullAdder U83 (w365, w359, IN24[0], w366, w367);
  HalfAdder U84 (w362, IN22[3], Out1[22], w369);
  FullAdder U85 (w369, w364, IN23[2], w370, w371);
  FullAdder U86 (w371, w366, IN24[1], w372, w373);
  FullAdder U87 (w373, w367, IN25[0], w374, w375);
  HalfAdder U88 (w370, IN23[3], Out1[23], w377);
  FullAdder U89 (w377, w372, IN24[2], w378, w379);
  FullAdder U90 (w379, w374, IN25[1], w380, w381);
  FullAdder U91 (w381, w375, IN26[0], w382, w383);
  HalfAdder U92 (w378, IN24[3], Out1[24], w385);
  FullAdder U93 (w385, w380, IN25[2], w386, w387);
  FullAdder U94 (w387, w382, IN26[1], w388, w389);
  FullAdder U95 (w389, w383, IN27[0], w390, w391);
  HalfAdder U96 (w386, IN25[3], Out1[25], w393);
  FullAdder U97 (w393, w388, IN26[2], w394, w395);
  FullAdder U98 (w395, w390, IN27[1], w396, w397);
  FullAdder U99 (w397, w391, IN28[0], w398, w399);
  HalfAdder U100 (w394, IN26[3], Out1[26], w401);
  FullAdder U101 (w401, w396, IN27[2], w402, w403);
  FullAdder U102 (w403, w398, IN28[1], w404, w405);
  FullAdder U103 (w405, w399, IN29[0], w406, w407);
  HalfAdder U104 (w402, IN27[3], Out1[27], w409);
  FullAdder U105 (w409, w404, IN28[2], w410, w411);
  FullAdder U106 (w411, w406, IN29[1], w412, w413);
  FullAdder U107 (w413, w407, IN30[0], w414, w415);
  HalfAdder U108 (w410, IN28[3], Out1[28], w417);
  FullAdder U109 (w417, w412, IN29[2], w418, w419);
  FullAdder U110 (w419, w414, IN30[1], w420, w421);
  FullAdder U111 (w421, w415, IN31[0], w422, w423);
  HalfAdder U112 (w418, IN29[3], Out1[29], w425);
  FullAdder U113 (w425, w420, IN30[2], w426, w427);
  FullAdder U114 (w427, w422, IN31[1], w428, w429);
  FullAdder U115 (w429, w423, IN32[0], w430, w431);
  HalfAdder U116 (w426, IN30[3], Out1[30], w433);
  FullAdder U117 (w433, w428, IN31[2], w434, w435);
  FullAdder U118 (w435, w430, IN32[1], w436, w437);
  FullAdder U119 (w437, w431, IN33[0], w438, w439);
  HalfAdder U120 (w434, IN31[3], Out1[31], w441);
  FullAdder U121 (w441, w436, IN32[2], w442, w443);
  FullAdder U122 (w443, w438, IN33[1], w444, w445);
  FullAdder U123 (w445, w439, IN34[0], w446, w447);
  HalfAdder U124 (w442, IN32[3], Out1[32], w449);
  FullAdder U125 (w449, w444, IN33[2], w450, w451);
  FullAdder U126 (w451, w446, IN34[1], w452, w453);
  FullAdder U127 (w453, w447, IN35[0], w454, w455);
  HalfAdder U128 (w450, IN33[3], Out1[33], w457);
  FullAdder U129 (w457, w452, IN34[2], w458, w459);
  FullAdder U130 (w459, w454, IN35[1], w460, w461);
  FullAdder U131 (w461, w455, IN36[0], w462, w463);
  HalfAdder U132 (w458, IN34[3], Out1[34], w465);
  FullAdder U133 (w465, w460, IN35[2], w466, w467);
  FullAdder U134 (w467, w462, IN36[1], w468, w469);
  FullAdder U135 (w469, w463, IN37[0], w470, w471);
  HalfAdder U136 (w466, IN35[3], Out1[35], w473);
  FullAdder U137 (w473, w468, IN36[2], w474, w475);
  FullAdder U138 (w475, w470, IN37[1], w476, w477);
  FullAdder U139 (w477, w471, IN38[0], w478, w479);
  HalfAdder U140 (w474, IN36[3], Out1[36], w481);
  FullAdder U141 (w481, w476, IN37[2], w482, w483);
  FullAdder U142 (w483, w478, IN38[1], w484, w485);
  FullAdder U143 (w485, w479, IN39[0], w486, w487);
  HalfAdder U144 (w482, IN37[3], Out1[37], w489);
  FullAdder U145 (w489, w484, IN38[2], w490, w491);
  FullAdder U146 (w491, w486, IN39[1], w492, w493);
  FullAdder U147 (w493, w487, IN40[0], w494, w495);
  HalfAdder U148 (w490, IN38[3], Out1[38], w497);
  FullAdder U149 (w497, w492, IN39[2], w498, w499);
  FullAdder U150 (w499, w494, IN40[1], w500, w501);
  FullAdder U151 (w501, w495, IN41[0], w502, w503);
  HalfAdder U152 (w498, IN39[3], Out1[39], w505);
  FullAdder U153 (w505, w500, IN40[2], Out1[40], w507);
  FullAdder U154 (w507, w502, IN41[1], Out1[41], w509);
  FullAdder U155 (w509, w503, IN42[0], Out1[42], Out1[43]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN5[4];
  assign Out2[1] = IN6[4];
  assign Out2[2] = IN7[4];
  assign Out2[3] = IN8[4];
  assign Out2[4] = IN9[4];
  assign Out2[5] = IN10[4];
  assign Out2[6] = IN11[4];
  assign Out2[7] = IN12[4];
  assign Out2[8] = IN13[4];
  assign Out2[9] = IN14[4];
  assign Out2[10] = IN15[4];
  assign Out2[11] = IN16[4];
  assign Out2[12] = IN17[4];
  assign Out2[13] = IN18[4];
  assign Out2[14] = IN19[4];
  assign Out2[15] = IN20[4];
  assign Out2[16] = IN21[4];
  assign Out2[17] = IN22[4];
  assign Out2[18] = IN23[4];
  assign Out2[19] = IN24[4];
  assign Out2[20] = IN25[4];
  assign Out2[21] = IN26[4];
  assign Out2[22] = IN27[4];
  assign Out2[23] = IN28[4];
  assign Out2[24] = IN29[4];
  assign Out2[25] = IN30[4];
  assign Out2[26] = IN31[4];
  assign Out2[27] = IN32[4];
  assign Out2[28] = IN33[4];
  assign Out2[29] = IN34[4];
  assign Out2[30] = IN35[4];
  assign Out2[31] = IN36[4];
  assign Out2[32] = IN37[4];
  assign Out2[33] = IN38[4];
  assign Out2[34] = IN39[4];
  assign Out2[35] = IN40[3];
  assign Out2[36] = IN41[2];
  assign Out2[37] = IN42[1];
  assign Out2[38] = IN43[0];

endmodule
module RC_39_39(IN1, IN2, Out);
  input [38:0] IN1;
  input [38:0] IN2;
  output [39:0] Out;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w79);
  FullAdder U1 (IN1[1], IN2[1], w79, Out[1], w81);
  FullAdder U2 (IN1[2], IN2[2], w81, Out[2], w83);
  FullAdder U3 (IN1[3], IN2[3], w83, Out[3], w85);
  FullAdder U4 (IN1[4], IN2[4], w85, Out[4], w87);
  FullAdder U5 (IN1[5], IN2[5], w87, Out[5], w89);
  FullAdder U6 (IN1[6], IN2[6], w89, Out[6], w91);
  FullAdder U7 (IN1[7], IN2[7], w91, Out[7], w93);
  FullAdder U8 (IN1[8], IN2[8], w93, Out[8], w95);
  FullAdder U9 (IN1[9], IN2[9], w95, Out[9], w97);
  FullAdder U10 (IN1[10], IN2[10], w97, Out[10], w99);
  FullAdder U11 (IN1[11], IN2[11], w99, Out[11], w101);
  FullAdder U12 (IN1[12], IN2[12], w101, Out[12], w103);
  FullAdder U13 (IN1[13], IN2[13], w103, Out[13], w105);
  FullAdder U14 (IN1[14], IN2[14], w105, Out[14], w107);
  FullAdder U15 (IN1[15], IN2[15], w107, Out[15], w109);
  FullAdder U16 (IN1[16], IN2[16], w109, Out[16], w111);
  FullAdder U17 (IN1[17], IN2[17], w111, Out[17], w113);
  FullAdder U18 (IN1[18], IN2[18], w113, Out[18], w115);
  FullAdder U19 (IN1[19], IN2[19], w115, Out[19], w117);
  FullAdder U20 (IN1[20], IN2[20], w117, Out[20], w119);
  FullAdder U21 (IN1[21], IN2[21], w119, Out[21], w121);
  FullAdder U22 (IN1[22], IN2[22], w121, Out[22], w123);
  FullAdder U23 (IN1[23], IN2[23], w123, Out[23], w125);
  FullAdder U24 (IN1[24], IN2[24], w125, Out[24], w127);
  FullAdder U25 (IN1[25], IN2[25], w127, Out[25], w129);
  FullAdder U26 (IN1[26], IN2[26], w129, Out[26], w131);
  FullAdder U27 (IN1[27], IN2[27], w131, Out[27], w133);
  FullAdder U28 (IN1[28], IN2[28], w133, Out[28], w135);
  FullAdder U29 (IN1[29], IN2[29], w135, Out[29], w137);
  FullAdder U30 (IN1[30], IN2[30], w137, Out[30], w139);
  FullAdder U31 (IN1[31], IN2[31], w139, Out[31], w141);
  FullAdder U32 (IN1[32], IN2[32], w141, Out[32], w143);
  FullAdder U33 (IN1[33], IN2[33], w143, Out[33], w145);
  FullAdder U34 (IN1[34], IN2[34], w145, Out[34], w147);
  FullAdder U35 (IN1[35], IN2[35], w147, Out[35], w149);
  FullAdder U36 (IN1[36], IN2[36], w149, Out[36], w151);
  FullAdder U37 (IN1[37], IN2[37], w151, Out[37], w153);
  FullAdder U38 (IN1[38], IN2[38], w153, Out[38], Out[39]);

endmodule
module NR_5_40(IN1, IN2, Out);
  input [4:0] IN1;
  input [39:0] IN2;
  output [44:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [4:0] P5;
  wire [4:0] P6;
  wire [4:0] P7;
  wire [4:0] P8;
  wire [4:0] P9;
  wire [4:0] P10;
  wire [4:0] P11;
  wire [4:0] P12;
  wire [4:0] P13;
  wire [4:0] P14;
  wire [4:0] P15;
  wire [4:0] P16;
  wire [4:0] P17;
  wire [4:0] P18;
  wire [4:0] P19;
  wire [4:0] P20;
  wire [4:0] P21;
  wire [4:0] P22;
  wire [4:0] P23;
  wire [4:0] P24;
  wire [4:0] P25;
  wire [4:0] P26;
  wire [4:0] P27;
  wire [4:0] P28;
  wire [4:0] P29;
  wire [4:0] P30;
  wire [4:0] P31;
  wire [4:0] P32;
  wire [4:0] P33;
  wire [4:0] P34;
  wire [4:0] P35;
  wire [4:0] P36;
  wire [4:0] P37;
  wire [4:0] P38;
  wire [4:0] P39;
  wire [3:0] P40;
  wire [2:0] P41;
  wire [1:0] P42;
  wire [0:0] P43;
  wire [43:0] R1;
  wire [38:0] R2;
  wire [44:0] aOut;
  U_SP_5_40 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, R1, R2);
  RC_39_39 S2 (R1[43:5], R2, aOut[44:5]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign Out = aOut[44:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
