
module NR_36_1(
    input [35:0]IN1,
    input [0:0]IN2,
    output [35:0]Out
);
    assign Out = IN2;
endmodule
