//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 53
  second input length: 11
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_53_11(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  input [52:0] IN1;
  input [10:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [10:0] P11;
  output [10:0] P12;
  output [10:0] P13;
  output [10:0] P14;
  output [10:0] P15;
  output [10:0] P16;
  output [10:0] P17;
  output [10:0] P18;
  output [10:0] P19;
  output [10:0] P20;
  output [10:0] P21;
  output [10:0] P22;
  output [10:0] P23;
  output [10:0] P24;
  output [10:0] P25;
  output [10:0] P26;
  output [10:0] P27;
  output [10:0] P28;
  output [10:0] P29;
  output [10:0] P30;
  output [10:0] P31;
  output [10:0] P32;
  output [10:0] P33;
  output [10:0] P34;
  output [10:0] P35;
  output [10:0] P36;
  output [10:0] P37;
  output [10:0] P38;
  output [10:0] P39;
  output [10:0] P40;
  output [10:0] P41;
  output [10:0] P42;
  output [10:0] P43;
  output [10:0] P44;
  output [10:0] P45;
  output [10:0] P46;
  output [10:0] P47;
  output [10:0] P48;
  output [10:0] P49;
  output [10:0] P50;
  output [10:0] P51;
  output [10:0] P52;
  output [9:0] P53;
  output [8:0] P54;
  output [7:0] P55;
  output [6:0] P56;
  output [5:0] P57;
  output [4:0] P58;
  output [3:0] P59;
  output [2:0] P60;
  output [1:0] P61;
  output [0:0] P62;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[0] = IN1[1]&IN2[10];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[1] = IN1[2]&IN2[9];
  assign P12[0] = IN1[2]&IN2[10];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[2] = IN1[3]&IN2[8];
  assign P12[1] = IN1[3]&IN2[9];
  assign P13[0] = IN1[3]&IN2[10];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[3] = IN1[4]&IN2[7];
  assign P12[2] = IN1[4]&IN2[8];
  assign P13[1] = IN1[4]&IN2[9];
  assign P14[0] = IN1[4]&IN2[10];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[4] = IN1[5]&IN2[6];
  assign P12[3] = IN1[5]&IN2[7];
  assign P13[2] = IN1[5]&IN2[8];
  assign P14[1] = IN1[5]&IN2[9];
  assign P15[0] = IN1[5]&IN2[10];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[5] = IN1[6]&IN2[5];
  assign P12[4] = IN1[6]&IN2[6];
  assign P13[3] = IN1[6]&IN2[7];
  assign P14[2] = IN1[6]&IN2[8];
  assign P15[1] = IN1[6]&IN2[9];
  assign P16[0] = IN1[6]&IN2[10];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[6] = IN1[7]&IN2[4];
  assign P12[5] = IN1[7]&IN2[5];
  assign P13[4] = IN1[7]&IN2[6];
  assign P14[3] = IN1[7]&IN2[7];
  assign P15[2] = IN1[7]&IN2[8];
  assign P16[1] = IN1[7]&IN2[9];
  assign P17[0] = IN1[7]&IN2[10];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[7] = IN1[8]&IN2[3];
  assign P12[6] = IN1[8]&IN2[4];
  assign P13[5] = IN1[8]&IN2[5];
  assign P14[4] = IN1[8]&IN2[6];
  assign P15[3] = IN1[8]&IN2[7];
  assign P16[2] = IN1[8]&IN2[8];
  assign P17[1] = IN1[8]&IN2[9];
  assign P18[0] = IN1[8]&IN2[10];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[8] = IN1[9]&IN2[2];
  assign P12[7] = IN1[9]&IN2[3];
  assign P13[6] = IN1[9]&IN2[4];
  assign P14[5] = IN1[9]&IN2[5];
  assign P15[4] = IN1[9]&IN2[6];
  assign P16[3] = IN1[9]&IN2[7];
  assign P17[2] = IN1[9]&IN2[8];
  assign P18[1] = IN1[9]&IN2[9];
  assign P19[0] = IN1[9]&IN2[10];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[9] = IN1[10]&IN2[1];
  assign P12[8] = IN1[10]&IN2[2];
  assign P13[7] = IN1[10]&IN2[3];
  assign P14[6] = IN1[10]&IN2[4];
  assign P15[5] = IN1[10]&IN2[5];
  assign P16[4] = IN1[10]&IN2[6];
  assign P17[3] = IN1[10]&IN2[7];
  assign P18[2] = IN1[10]&IN2[8];
  assign P19[1] = IN1[10]&IN2[9];
  assign P20[0] = IN1[10]&IN2[10];
  assign P11[10] = IN1[11]&IN2[0];
  assign P12[9] = IN1[11]&IN2[1];
  assign P13[8] = IN1[11]&IN2[2];
  assign P14[7] = IN1[11]&IN2[3];
  assign P15[6] = IN1[11]&IN2[4];
  assign P16[5] = IN1[11]&IN2[5];
  assign P17[4] = IN1[11]&IN2[6];
  assign P18[3] = IN1[11]&IN2[7];
  assign P19[2] = IN1[11]&IN2[8];
  assign P20[1] = IN1[11]&IN2[9];
  assign P21[0] = IN1[11]&IN2[10];
  assign P12[10] = IN1[12]&IN2[0];
  assign P13[9] = IN1[12]&IN2[1];
  assign P14[8] = IN1[12]&IN2[2];
  assign P15[7] = IN1[12]&IN2[3];
  assign P16[6] = IN1[12]&IN2[4];
  assign P17[5] = IN1[12]&IN2[5];
  assign P18[4] = IN1[12]&IN2[6];
  assign P19[3] = IN1[12]&IN2[7];
  assign P20[2] = IN1[12]&IN2[8];
  assign P21[1] = IN1[12]&IN2[9];
  assign P22[0] = IN1[12]&IN2[10];
  assign P13[10] = IN1[13]&IN2[0];
  assign P14[9] = IN1[13]&IN2[1];
  assign P15[8] = IN1[13]&IN2[2];
  assign P16[7] = IN1[13]&IN2[3];
  assign P17[6] = IN1[13]&IN2[4];
  assign P18[5] = IN1[13]&IN2[5];
  assign P19[4] = IN1[13]&IN2[6];
  assign P20[3] = IN1[13]&IN2[7];
  assign P21[2] = IN1[13]&IN2[8];
  assign P22[1] = IN1[13]&IN2[9];
  assign P23[0] = IN1[13]&IN2[10];
  assign P14[10] = IN1[14]&IN2[0];
  assign P15[9] = IN1[14]&IN2[1];
  assign P16[8] = IN1[14]&IN2[2];
  assign P17[7] = IN1[14]&IN2[3];
  assign P18[6] = IN1[14]&IN2[4];
  assign P19[5] = IN1[14]&IN2[5];
  assign P20[4] = IN1[14]&IN2[6];
  assign P21[3] = IN1[14]&IN2[7];
  assign P22[2] = IN1[14]&IN2[8];
  assign P23[1] = IN1[14]&IN2[9];
  assign P24[0] = IN1[14]&IN2[10];
  assign P15[10] = IN1[15]&IN2[0];
  assign P16[9] = IN1[15]&IN2[1];
  assign P17[8] = IN1[15]&IN2[2];
  assign P18[7] = IN1[15]&IN2[3];
  assign P19[6] = IN1[15]&IN2[4];
  assign P20[5] = IN1[15]&IN2[5];
  assign P21[4] = IN1[15]&IN2[6];
  assign P22[3] = IN1[15]&IN2[7];
  assign P23[2] = IN1[15]&IN2[8];
  assign P24[1] = IN1[15]&IN2[9];
  assign P25[0] = IN1[15]&IN2[10];
  assign P16[10] = IN1[16]&IN2[0];
  assign P17[9] = IN1[16]&IN2[1];
  assign P18[8] = IN1[16]&IN2[2];
  assign P19[7] = IN1[16]&IN2[3];
  assign P20[6] = IN1[16]&IN2[4];
  assign P21[5] = IN1[16]&IN2[5];
  assign P22[4] = IN1[16]&IN2[6];
  assign P23[3] = IN1[16]&IN2[7];
  assign P24[2] = IN1[16]&IN2[8];
  assign P25[1] = IN1[16]&IN2[9];
  assign P26[0] = IN1[16]&IN2[10];
  assign P17[10] = IN1[17]&IN2[0];
  assign P18[9] = IN1[17]&IN2[1];
  assign P19[8] = IN1[17]&IN2[2];
  assign P20[7] = IN1[17]&IN2[3];
  assign P21[6] = IN1[17]&IN2[4];
  assign P22[5] = IN1[17]&IN2[5];
  assign P23[4] = IN1[17]&IN2[6];
  assign P24[3] = IN1[17]&IN2[7];
  assign P25[2] = IN1[17]&IN2[8];
  assign P26[1] = IN1[17]&IN2[9];
  assign P27[0] = IN1[17]&IN2[10];
  assign P18[10] = IN1[18]&IN2[0];
  assign P19[9] = IN1[18]&IN2[1];
  assign P20[8] = IN1[18]&IN2[2];
  assign P21[7] = IN1[18]&IN2[3];
  assign P22[6] = IN1[18]&IN2[4];
  assign P23[5] = IN1[18]&IN2[5];
  assign P24[4] = IN1[18]&IN2[6];
  assign P25[3] = IN1[18]&IN2[7];
  assign P26[2] = IN1[18]&IN2[8];
  assign P27[1] = IN1[18]&IN2[9];
  assign P28[0] = IN1[18]&IN2[10];
  assign P19[10] = IN1[19]&IN2[0];
  assign P20[9] = IN1[19]&IN2[1];
  assign P21[8] = IN1[19]&IN2[2];
  assign P22[7] = IN1[19]&IN2[3];
  assign P23[6] = IN1[19]&IN2[4];
  assign P24[5] = IN1[19]&IN2[5];
  assign P25[4] = IN1[19]&IN2[6];
  assign P26[3] = IN1[19]&IN2[7];
  assign P27[2] = IN1[19]&IN2[8];
  assign P28[1] = IN1[19]&IN2[9];
  assign P29[0] = IN1[19]&IN2[10];
  assign P20[10] = IN1[20]&IN2[0];
  assign P21[9] = IN1[20]&IN2[1];
  assign P22[8] = IN1[20]&IN2[2];
  assign P23[7] = IN1[20]&IN2[3];
  assign P24[6] = IN1[20]&IN2[4];
  assign P25[5] = IN1[20]&IN2[5];
  assign P26[4] = IN1[20]&IN2[6];
  assign P27[3] = IN1[20]&IN2[7];
  assign P28[2] = IN1[20]&IN2[8];
  assign P29[1] = IN1[20]&IN2[9];
  assign P30[0] = IN1[20]&IN2[10];
  assign P21[10] = IN1[21]&IN2[0];
  assign P22[9] = IN1[21]&IN2[1];
  assign P23[8] = IN1[21]&IN2[2];
  assign P24[7] = IN1[21]&IN2[3];
  assign P25[6] = IN1[21]&IN2[4];
  assign P26[5] = IN1[21]&IN2[5];
  assign P27[4] = IN1[21]&IN2[6];
  assign P28[3] = IN1[21]&IN2[7];
  assign P29[2] = IN1[21]&IN2[8];
  assign P30[1] = IN1[21]&IN2[9];
  assign P31[0] = IN1[21]&IN2[10];
  assign P22[10] = IN1[22]&IN2[0];
  assign P23[9] = IN1[22]&IN2[1];
  assign P24[8] = IN1[22]&IN2[2];
  assign P25[7] = IN1[22]&IN2[3];
  assign P26[6] = IN1[22]&IN2[4];
  assign P27[5] = IN1[22]&IN2[5];
  assign P28[4] = IN1[22]&IN2[6];
  assign P29[3] = IN1[22]&IN2[7];
  assign P30[2] = IN1[22]&IN2[8];
  assign P31[1] = IN1[22]&IN2[9];
  assign P32[0] = IN1[22]&IN2[10];
  assign P23[10] = IN1[23]&IN2[0];
  assign P24[9] = IN1[23]&IN2[1];
  assign P25[8] = IN1[23]&IN2[2];
  assign P26[7] = IN1[23]&IN2[3];
  assign P27[6] = IN1[23]&IN2[4];
  assign P28[5] = IN1[23]&IN2[5];
  assign P29[4] = IN1[23]&IN2[6];
  assign P30[3] = IN1[23]&IN2[7];
  assign P31[2] = IN1[23]&IN2[8];
  assign P32[1] = IN1[23]&IN2[9];
  assign P33[0] = IN1[23]&IN2[10];
  assign P24[10] = IN1[24]&IN2[0];
  assign P25[9] = IN1[24]&IN2[1];
  assign P26[8] = IN1[24]&IN2[2];
  assign P27[7] = IN1[24]&IN2[3];
  assign P28[6] = IN1[24]&IN2[4];
  assign P29[5] = IN1[24]&IN2[5];
  assign P30[4] = IN1[24]&IN2[6];
  assign P31[3] = IN1[24]&IN2[7];
  assign P32[2] = IN1[24]&IN2[8];
  assign P33[1] = IN1[24]&IN2[9];
  assign P34[0] = IN1[24]&IN2[10];
  assign P25[10] = IN1[25]&IN2[0];
  assign P26[9] = IN1[25]&IN2[1];
  assign P27[8] = IN1[25]&IN2[2];
  assign P28[7] = IN1[25]&IN2[3];
  assign P29[6] = IN1[25]&IN2[4];
  assign P30[5] = IN1[25]&IN2[5];
  assign P31[4] = IN1[25]&IN2[6];
  assign P32[3] = IN1[25]&IN2[7];
  assign P33[2] = IN1[25]&IN2[8];
  assign P34[1] = IN1[25]&IN2[9];
  assign P35[0] = IN1[25]&IN2[10];
  assign P26[10] = IN1[26]&IN2[0];
  assign P27[9] = IN1[26]&IN2[1];
  assign P28[8] = IN1[26]&IN2[2];
  assign P29[7] = IN1[26]&IN2[3];
  assign P30[6] = IN1[26]&IN2[4];
  assign P31[5] = IN1[26]&IN2[5];
  assign P32[4] = IN1[26]&IN2[6];
  assign P33[3] = IN1[26]&IN2[7];
  assign P34[2] = IN1[26]&IN2[8];
  assign P35[1] = IN1[26]&IN2[9];
  assign P36[0] = IN1[26]&IN2[10];
  assign P27[10] = IN1[27]&IN2[0];
  assign P28[9] = IN1[27]&IN2[1];
  assign P29[8] = IN1[27]&IN2[2];
  assign P30[7] = IN1[27]&IN2[3];
  assign P31[6] = IN1[27]&IN2[4];
  assign P32[5] = IN1[27]&IN2[5];
  assign P33[4] = IN1[27]&IN2[6];
  assign P34[3] = IN1[27]&IN2[7];
  assign P35[2] = IN1[27]&IN2[8];
  assign P36[1] = IN1[27]&IN2[9];
  assign P37[0] = IN1[27]&IN2[10];
  assign P28[10] = IN1[28]&IN2[0];
  assign P29[9] = IN1[28]&IN2[1];
  assign P30[8] = IN1[28]&IN2[2];
  assign P31[7] = IN1[28]&IN2[3];
  assign P32[6] = IN1[28]&IN2[4];
  assign P33[5] = IN1[28]&IN2[5];
  assign P34[4] = IN1[28]&IN2[6];
  assign P35[3] = IN1[28]&IN2[7];
  assign P36[2] = IN1[28]&IN2[8];
  assign P37[1] = IN1[28]&IN2[9];
  assign P38[0] = IN1[28]&IN2[10];
  assign P29[10] = IN1[29]&IN2[0];
  assign P30[9] = IN1[29]&IN2[1];
  assign P31[8] = IN1[29]&IN2[2];
  assign P32[7] = IN1[29]&IN2[3];
  assign P33[6] = IN1[29]&IN2[4];
  assign P34[5] = IN1[29]&IN2[5];
  assign P35[4] = IN1[29]&IN2[6];
  assign P36[3] = IN1[29]&IN2[7];
  assign P37[2] = IN1[29]&IN2[8];
  assign P38[1] = IN1[29]&IN2[9];
  assign P39[0] = IN1[29]&IN2[10];
  assign P30[10] = IN1[30]&IN2[0];
  assign P31[9] = IN1[30]&IN2[1];
  assign P32[8] = IN1[30]&IN2[2];
  assign P33[7] = IN1[30]&IN2[3];
  assign P34[6] = IN1[30]&IN2[4];
  assign P35[5] = IN1[30]&IN2[5];
  assign P36[4] = IN1[30]&IN2[6];
  assign P37[3] = IN1[30]&IN2[7];
  assign P38[2] = IN1[30]&IN2[8];
  assign P39[1] = IN1[30]&IN2[9];
  assign P40[0] = IN1[30]&IN2[10];
  assign P31[10] = IN1[31]&IN2[0];
  assign P32[9] = IN1[31]&IN2[1];
  assign P33[8] = IN1[31]&IN2[2];
  assign P34[7] = IN1[31]&IN2[3];
  assign P35[6] = IN1[31]&IN2[4];
  assign P36[5] = IN1[31]&IN2[5];
  assign P37[4] = IN1[31]&IN2[6];
  assign P38[3] = IN1[31]&IN2[7];
  assign P39[2] = IN1[31]&IN2[8];
  assign P40[1] = IN1[31]&IN2[9];
  assign P41[0] = IN1[31]&IN2[10];
  assign P32[10] = IN1[32]&IN2[0];
  assign P33[9] = IN1[32]&IN2[1];
  assign P34[8] = IN1[32]&IN2[2];
  assign P35[7] = IN1[32]&IN2[3];
  assign P36[6] = IN1[32]&IN2[4];
  assign P37[5] = IN1[32]&IN2[5];
  assign P38[4] = IN1[32]&IN2[6];
  assign P39[3] = IN1[32]&IN2[7];
  assign P40[2] = IN1[32]&IN2[8];
  assign P41[1] = IN1[32]&IN2[9];
  assign P42[0] = IN1[32]&IN2[10];
  assign P33[10] = IN1[33]&IN2[0];
  assign P34[9] = IN1[33]&IN2[1];
  assign P35[8] = IN1[33]&IN2[2];
  assign P36[7] = IN1[33]&IN2[3];
  assign P37[6] = IN1[33]&IN2[4];
  assign P38[5] = IN1[33]&IN2[5];
  assign P39[4] = IN1[33]&IN2[6];
  assign P40[3] = IN1[33]&IN2[7];
  assign P41[2] = IN1[33]&IN2[8];
  assign P42[1] = IN1[33]&IN2[9];
  assign P43[0] = IN1[33]&IN2[10];
  assign P34[10] = IN1[34]&IN2[0];
  assign P35[9] = IN1[34]&IN2[1];
  assign P36[8] = IN1[34]&IN2[2];
  assign P37[7] = IN1[34]&IN2[3];
  assign P38[6] = IN1[34]&IN2[4];
  assign P39[5] = IN1[34]&IN2[5];
  assign P40[4] = IN1[34]&IN2[6];
  assign P41[3] = IN1[34]&IN2[7];
  assign P42[2] = IN1[34]&IN2[8];
  assign P43[1] = IN1[34]&IN2[9];
  assign P44[0] = IN1[34]&IN2[10];
  assign P35[10] = IN1[35]&IN2[0];
  assign P36[9] = IN1[35]&IN2[1];
  assign P37[8] = IN1[35]&IN2[2];
  assign P38[7] = IN1[35]&IN2[3];
  assign P39[6] = IN1[35]&IN2[4];
  assign P40[5] = IN1[35]&IN2[5];
  assign P41[4] = IN1[35]&IN2[6];
  assign P42[3] = IN1[35]&IN2[7];
  assign P43[2] = IN1[35]&IN2[8];
  assign P44[1] = IN1[35]&IN2[9];
  assign P45[0] = IN1[35]&IN2[10];
  assign P36[10] = IN1[36]&IN2[0];
  assign P37[9] = IN1[36]&IN2[1];
  assign P38[8] = IN1[36]&IN2[2];
  assign P39[7] = IN1[36]&IN2[3];
  assign P40[6] = IN1[36]&IN2[4];
  assign P41[5] = IN1[36]&IN2[5];
  assign P42[4] = IN1[36]&IN2[6];
  assign P43[3] = IN1[36]&IN2[7];
  assign P44[2] = IN1[36]&IN2[8];
  assign P45[1] = IN1[36]&IN2[9];
  assign P46[0] = IN1[36]&IN2[10];
  assign P37[10] = IN1[37]&IN2[0];
  assign P38[9] = IN1[37]&IN2[1];
  assign P39[8] = IN1[37]&IN2[2];
  assign P40[7] = IN1[37]&IN2[3];
  assign P41[6] = IN1[37]&IN2[4];
  assign P42[5] = IN1[37]&IN2[5];
  assign P43[4] = IN1[37]&IN2[6];
  assign P44[3] = IN1[37]&IN2[7];
  assign P45[2] = IN1[37]&IN2[8];
  assign P46[1] = IN1[37]&IN2[9];
  assign P47[0] = IN1[37]&IN2[10];
  assign P38[10] = IN1[38]&IN2[0];
  assign P39[9] = IN1[38]&IN2[1];
  assign P40[8] = IN1[38]&IN2[2];
  assign P41[7] = IN1[38]&IN2[3];
  assign P42[6] = IN1[38]&IN2[4];
  assign P43[5] = IN1[38]&IN2[5];
  assign P44[4] = IN1[38]&IN2[6];
  assign P45[3] = IN1[38]&IN2[7];
  assign P46[2] = IN1[38]&IN2[8];
  assign P47[1] = IN1[38]&IN2[9];
  assign P48[0] = IN1[38]&IN2[10];
  assign P39[10] = IN1[39]&IN2[0];
  assign P40[9] = IN1[39]&IN2[1];
  assign P41[8] = IN1[39]&IN2[2];
  assign P42[7] = IN1[39]&IN2[3];
  assign P43[6] = IN1[39]&IN2[4];
  assign P44[5] = IN1[39]&IN2[5];
  assign P45[4] = IN1[39]&IN2[6];
  assign P46[3] = IN1[39]&IN2[7];
  assign P47[2] = IN1[39]&IN2[8];
  assign P48[1] = IN1[39]&IN2[9];
  assign P49[0] = IN1[39]&IN2[10];
  assign P40[10] = IN1[40]&IN2[0];
  assign P41[9] = IN1[40]&IN2[1];
  assign P42[8] = IN1[40]&IN2[2];
  assign P43[7] = IN1[40]&IN2[3];
  assign P44[6] = IN1[40]&IN2[4];
  assign P45[5] = IN1[40]&IN2[5];
  assign P46[4] = IN1[40]&IN2[6];
  assign P47[3] = IN1[40]&IN2[7];
  assign P48[2] = IN1[40]&IN2[8];
  assign P49[1] = IN1[40]&IN2[9];
  assign P50[0] = IN1[40]&IN2[10];
  assign P41[10] = IN1[41]&IN2[0];
  assign P42[9] = IN1[41]&IN2[1];
  assign P43[8] = IN1[41]&IN2[2];
  assign P44[7] = IN1[41]&IN2[3];
  assign P45[6] = IN1[41]&IN2[4];
  assign P46[5] = IN1[41]&IN2[5];
  assign P47[4] = IN1[41]&IN2[6];
  assign P48[3] = IN1[41]&IN2[7];
  assign P49[2] = IN1[41]&IN2[8];
  assign P50[1] = IN1[41]&IN2[9];
  assign P51[0] = IN1[41]&IN2[10];
  assign P42[10] = IN1[42]&IN2[0];
  assign P43[9] = IN1[42]&IN2[1];
  assign P44[8] = IN1[42]&IN2[2];
  assign P45[7] = IN1[42]&IN2[3];
  assign P46[6] = IN1[42]&IN2[4];
  assign P47[5] = IN1[42]&IN2[5];
  assign P48[4] = IN1[42]&IN2[6];
  assign P49[3] = IN1[42]&IN2[7];
  assign P50[2] = IN1[42]&IN2[8];
  assign P51[1] = IN1[42]&IN2[9];
  assign P52[0] = IN1[42]&IN2[10];
  assign P43[10] = IN1[43]&IN2[0];
  assign P44[9] = IN1[43]&IN2[1];
  assign P45[8] = IN1[43]&IN2[2];
  assign P46[7] = IN1[43]&IN2[3];
  assign P47[6] = IN1[43]&IN2[4];
  assign P48[5] = IN1[43]&IN2[5];
  assign P49[4] = IN1[43]&IN2[6];
  assign P50[3] = IN1[43]&IN2[7];
  assign P51[2] = IN1[43]&IN2[8];
  assign P52[1] = IN1[43]&IN2[9];
  assign P53[0] = IN1[43]&IN2[10];
  assign P44[10] = IN1[44]&IN2[0];
  assign P45[9] = IN1[44]&IN2[1];
  assign P46[8] = IN1[44]&IN2[2];
  assign P47[7] = IN1[44]&IN2[3];
  assign P48[6] = IN1[44]&IN2[4];
  assign P49[5] = IN1[44]&IN2[5];
  assign P50[4] = IN1[44]&IN2[6];
  assign P51[3] = IN1[44]&IN2[7];
  assign P52[2] = IN1[44]&IN2[8];
  assign P53[1] = IN1[44]&IN2[9];
  assign P54[0] = IN1[44]&IN2[10];
  assign P45[10] = IN1[45]&IN2[0];
  assign P46[9] = IN1[45]&IN2[1];
  assign P47[8] = IN1[45]&IN2[2];
  assign P48[7] = IN1[45]&IN2[3];
  assign P49[6] = IN1[45]&IN2[4];
  assign P50[5] = IN1[45]&IN2[5];
  assign P51[4] = IN1[45]&IN2[6];
  assign P52[3] = IN1[45]&IN2[7];
  assign P53[2] = IN1[45]&IN2[8];
  assign P54[1] = IN1[45]&IN2[9];
  assign P55[0] = IN1[45]&IN2[10];
  assign P46[10] = IN1[46]&IN2[0];
  assign P47[9] = IN1[46]&IN2[1];
  assign P48[8] = IN1[46]&IN2[2];
  assign P49[7] = IN1[46]&IN2[3];
  assign P50[6] = IN1[46]&IN2[4];
  assign P51[5] = IN1[46]&IN2[5];
  assign P52[4] = IN1[46]&IN2[6];
  assign P53[3] = IN1[46]&IN2[7];
  assign P54[2] = IN1[46]&IN2[8];
  assign P55[1] = IN1[46]&IN2[9];
  assign P56[0] = IN1[46]&IN2[10];
  assign P47[10] = IN1[47]&IN2[0];
  assign P48[9] = IN1[47]&IN2[1];
  assign P49[8] = IN1[47]&IN2[2];
  assign P50[7] = IN1[47]&IN2[3];
  assign P51[6] = IN1[47]&IN2[4];
  assign P52[5] = IN1[47]&IN2[5];
  assign P53[4] = IN1[47]&IN2[6];
  assign P54[3] = IN1[47]&IN2[7];
  assign P55[2] = IN1[47]&IN2[8];
  assign P56[1] = IN1[47]&IN2[9];
  assign P57[0] = IN1[47]&IN2[10];
  assign P48[10] = IN1[48]&IN2[0];
  assign P49[9] = IN1[48]&IN2[1];
  assign P50[8] = IN1[48]&IN2[2];
  assign P51[7] = IN1[48]&IN2[3];
  assign P52[6] = IN1[48]&IN2[4];
  assign P53[5] = IN1[48]&IN2[5];
  assign P54[4] = IN1[48]&IN2[6];
  assign P55[3] = IN1[48]&IN2[7];
  assign P56[2] = IN1[48]&IN2[8];
  assign P57[1] = IN1[48]&IN2[9];
  assign P58[0] = IN1[48]&IN2[10];
  assign P49[10] = IN1[49]&IN2[0];
  assign P50[9] = IN1[49]&IN2[1];
  assign P51[8] = IN1[49]&IN2[2];
  assign P52[7] = IN1[49]&IN2[3];
  assign P53[6] = IN1[49]&IN2[4];
  assign P54[5] = IN1[49]&IN2[5];
  assign P55[4] = IN1[49]&IN2[6];
  assign P56[3] = IN1[49]&IN2[7];
  assign P57[2] = IN1[49]&IN2[8];
  assign P58[1] = IN1[49]&IN2[9];
  assign P59[0] = IN1[49]&IN2[10];
  assign P50[10] = IN1[50]&IN2[0];
  assign P51[9] = IN1[50]&IN2[1];
  assign P52[8] = IN1[50]&IN2[2];
  assign P53[7] = IN1[50]&IN2[3];
  assign P54[6] = IN1[50]&IN2[4];
  assign P55[5] = IN1[50]&IN2[5];
  assign P56[4] = IN1[50]&IN2[6];
  assign P57[3] = IN1[50]&IN2[7];
  assign P58[2] = IN1[50]&IN2[8];
  assign P59[1] = IN1[50]&IN2[9];
  assign P60[0] = IN1[50]&IN2[10];
  assign P51[10] = IN1[51]&IN2[0];
  assign P52[9] = IN1[51]&IN2[1];
  assign P53[8] = IN1[51]&IN2[2];
  assign P54[7] = IN1[51]&IN2[3];
  assign P55[6] = IN1[51]&IN2[4];
  assign P56[5] = IN1[51]&IN2[5];
  assign P57[4] = IN1[51]&IN2[6];
  assign P58[3] = IN1[51]&IN2[7];
  assign P59[2] = IN1[51]&IN2[8];
  assign P60[1] = IN1[51]&IN2[9];
  assign P61[0] = IN1[51]&IN2[10];
  assign P52[10] = IN1[52]&IN2[0];
  assign P53[9] = IN1[52]&IN2[1];
  assign P54[8] = IN1[52]&IN2[2];
  assign P55[7] = IN1[52]&IN2[3];
  assign P56[6] = IN1[52]&IN2[4];
  assign P57[5] = IN1[52]&IN2[5];
  assign P58[4] = IN1[52]&IN2[6];
  assign P59[3] = IN1[52]&IN2[7];
  assign P60[2] = IN1[52]&IN2[8];
  assign P61[1] = IN1[52]&IN2[9];
  assign P62[0] = IN1[52]&IN2[10];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [10:0] IN11;
  input [10:0] IN12;
  input [10:0] IN13;
  input [10:0] IN14;
  input [10:0] IN15;
  input [10:0] IN16;
  input [10:0] IN17;
  input [10:0] IN18;
  input [10:0] IN19;
  input [10:0] IN20;
  input [10:0] IN21;
  input [10:0] IN22;
  input [10:0] IN23;
  input [10:0] IN24;
  input [10:0] IN25;
  input [10:0] IN26;
  input [10:0] IN27;
  input [10:0] IN28;
  input [10:0] IN29;
  input [10:0] IN30;
  input [10:0] IN31;
  input [10:0] IN32;
  input [10:0] IN33;
  input [10:0] IN34;
  input [10:0] IN35;
  input [10:0] IN36;
  input [10:0] IN37;
  input [10:0] IN38;
  input [10:0] IN39;
  input [10:0] IN40;
  input [10:0] IN41;
  input [10:0] IN42;
  input [10:0] IN43;
  input [10:0] IN44;
  input [10:0] IN45;
  input [10:0] IN46;
  input [10:0] IN47;
  input [10:0] IN48;
  input [10:0] IN49;
  input [10:0] IN50;
  input [10:0] IN51;
  input [10:0] IN52;
  input [9:0] IN53;
  input [8:0] IN54;
  input [7:0] IN55;
  input [6:0] IN56;
  input [5:0] IN57;
  input [4:0] IN58;
  input [3:0] IN59;
  input [2:0] IN60;
  input [1:0] IN61;
  input [0:0] IN62;
  output [62:0] Out1;
  output [9:0] Out2;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1520;
  wire w1522;
  wire w1524;
  wire w1526;
  wire w1528;
  wire w1530;
  wire w1532;
  wire w1534;
  wire w1536;
  wire w1538;
  wire w1540;
  wire w1542;
  wire w1544;
  wire w1546;
  wire w1548;
  wire w1550;
  wire w1552;
  wire w1554;
  wire w1556;
  wire w1558;
  wire w1560;
  wire w1562;
  wire w1564;
  wire w1566;
  wire w1568;
  wire w1570;
  wire w1572;
  wire w1574;
  wire w1576;
  wire w1578;
  wire w1580;
  wire w1582;
  wire w1584;
  wire w1586;
  wire w1588;
  wire w1590;
  wire w1592;
  wire w1594;
  wire w1596;
  wire w1598;
  wire w1600;
  wire w1602;
  wire w1604;
  wire w1606;
  wire w1608;
  wire w1610;
  wire w1612;
  wire w1614;
  wire w1616;
  wire w1618;
  wire w1620;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w584);
  FullAdder U1 (w584, IN2[0], IN2[1], w585, w586);
  FullAdder U2 (w586, IN3[0], IN3[1], w587, w588);
  FullAdder U3 (w588, IN4[0], IN4[1], w589, w590);
  FullAdder U4 (w590, IN5[0], IN5[1], w591, w592);
  FullAdder U5 (w592, IN6[0], IN6[1], w593, w594);
  FullAdder U6 (w594, IN7[0], IN7[1], w595, w596);
  FullAdder U7 (w596, IN8[0], IN8[1], w597, w598);
  FullAdder U8 (w598, IN9[0], IN9[1], w599, w600);
  FullAdder U9 (w600, IN10[0], IN10[1], w601, w602);
  FullAdder U10 (w602, IN11[0], IN11[1], w603, w604);
  FullAdder U11 (w604, IN12[0], IN12[1], w605, w606);
  FullAdder U12 (w606, IN13[0], IN13[1], w607, w608);
  FullAdder U13 (w608, IN14[0], IN14[1], w609, w610);
  FullAdder U14 (w610, IN15[0], IN15[1], w611, w612);
  FullAdder U15 (w612, IN16[0], IN16[1], w613, w614);
  FullAdder U16 (w614, IN17[0], IN17[1], w615, w616);
  FullAdder U17 (w616, IN18[0], IN18[1], w617, w618);
  FullAdder U18 (w618, IN19[0], IN19[1], w619, w620);
  FullAdder U19 (w620, IN20[0], IN20[1], w621, w622);
  FullAdder U20 (w622, IN21[0], IN21[1], w623, w624);
  FullAdder U21 (w624, IN22[0], IN22[1], w625, w626);
  FullAdder U22 (w626, IN23[0], IN23[1], w627, w628);
  FullAdder U23 (w628, IN24[0], IN24[1], w629, w630);
  FullAdder U24 (w630, IN25[0], IN25[1], w631, w632);
  FullAdder U25 (w632, IN26[0], IN26[1], w633, w634);
  FullAdder U26 (w634, IN27[0], IN27[1], w635, w636);
  FullAdder U27 (w636, IN28[0], IN28[1], w637, w638);
  FullAdder U28 (w638, IN29[0], IN29[1], w639, w640);
  FullAdder U29 (w640, IN30[0], IN30[1], w641, w642);
  FullAdder U30 (w642, IN31[0], IN31[1], w643, w644);
  FullAdder U31 (w644, IN32[0], IN32[1], w645, w646);
  FullAdder U32 (w646, IN33[0], IN33[1], w647, w648);
  FullAdder U33 (w648, IN34[0], IN34[1], w649, w650);
  FullAdder U34 (w650, IN35[0], IN35[1], w651, w652);
  FullAdder U35 (w652, IN36[0], IN36[1], w653, w654);
  FullAdder U36 (w654, IN37[0], IN37[1], w655, w656);
  FullAdder U37 (w656, IN38[0], IN38[1], w657, w658);
  FullAdder U38 (w658, IN39[0], IN39[1], w659, w660);
  FullAdder U39 (w660, IN40[0], IN40[1], w661, w662);
  FullAdder U40 (w662, IN41[0], IN41[1], w663, w664);
  FullAdder U41 (w664, IN42[0], IN42[1], w665, w666);
  FullAdder U42 (w666, IN43[0], IN43[1], w667, w668);
  FullAdder U43 (w668, IN44[0], IN44[1], w669, w670);
  FullAdder U44 (w670, IN45[0], IN45[1], w671, w672);
  FullAdder U45 (w672, IN46[0], IN46[1], w673, w674);
  FullAdder U46 (w674, IN47[0], IN47[1], w675, w676);
  FullAdder U47 (w676, IN48[0], IN48[1], w677, w678);
  FullAdder U48 (w678, IN49[0], IN49[1], w679, w680);
  FullAdder U49 (w680, IN50[0], IN50[1], w681, w682);
  FullAdder U50 (w682, IN51[0], IN51[1], w683, w684);
  FullAdder U51 (w684, IN52[0], IN52[1], w685, w686);
  HalfAdder U52 (w585, IN2[2], Out1[2], w688);
  FullAdder U53 (w688, w587, IN3[2], w689, w690);
  FullAdder U54 (w690, w589, IN4[2], w691, w692);
  FullAdder U55 (w692, w591, IN5[2], w693, w694);
  FullAdder U56 (w694, w593, IN6[2], w695, w696);
  FullAdder U57 (w696, w595, IN7[2], w697, w698);
  FullAdder U58 (w698, w597, IN8[2], w699, w700);
  FullAdder U59 (w700, w599, IN9[2], w701, w702);
  FullAdder U60 (w702, w601, IN10[2], w703, w704);
  FullAdder U61 (w704, w603, IN11[2], w705, w706);
  FullAdder U62 (w706, w605, IN12[2], w707, w708);
  FullAdder U63 (w708, w607, IN13[2], w709, w710);
  FullAdder U64 (w710, w609, IN14[2], w711, w712);
  FullAdder U65 (w712, w611, IN15[2], w713, w714);
  FullAdder U66 (w714, w613, IN16[2], w715, w716);
  FullAdder U67 (w716, w615, IN17[2], w717, w718);
  FullAdder U68 (w718, w617, IN18[2], w719, w720);
  FullAdder U69 (w720, w619, IN19[2], w721, w722);
  FullAdder U70 (w722, w621, IN20[2], w723, w724);
  FullAdder U71 (w724, w623, IN21[2], w725, w726);
  FullAdder U72 (w726, w625, IN22[2], w727, w728);
  FullAdder U73 (w728, w627, IN23[2], w729, w730);
  FullAdder U74 (w730, w629, IN24[2], w731, w732);
  FullAdder U75 (w732, w631, IN25[2], w733, w734);
  FullAdder U76 (w734, w633, IN26[2], w735, w736);
  FullAdder U77 (w736, w635, IN27[2], w737, w738);
  FullAdder U78 (w738, w637, IN28[2], w739, w740);
  FullAdder U79 (w740, w639, IN29[2], w741, w742);
  FullAdder U80 (w742, w641, IN30[2], w743, w744);
  FullAdder U81 (w744, w643, IN31[2], w745, w746);
  FullAdder U82 (w746, w645, IN32[2], w747, w748);
  FullAdder U83 (w748, w647, IN33[2], w749, w750);
  FullAdder U84 (w750, w649, IN34[2], w751, w752);
  FullAdder U85 (w752, w651, IN35[2], w753, w754);
  FullAdder U86 (w754, w653, IN36[2], w755, w756);
  FullAdder U87 (w756, w655, IN37[2], w757, w758);
  FullAdder U88 (w758, w657, IN38[2], w759, w760);
  FullAdder U89 (w760, w659, IN39[2], w761, w762);
  FullAdder U90 (w762, w661, IN40[2], w763, w764);
  FullAdder U91 (w764, w663, IN41[2], w765, w766);
  FullAdder U92 (w766, w665, IN42[2], w767, w768);
  FullAdder U93 (w768, w667, IN43[2], w769, w770);
  FullAdder U94 (w770, w669, IN44[2], w771, w772);
  FullAdder U95 (w772, w671, IN45[2], w773, w774);
  FullAdder U96 (w774, w673, IN46[2], w775, w776);
  FullAdder U97 (w776, w675, IN47[2], w777, w778);
  FullAdder U98 (w778, w677, IN48[2], w779, w780);
  FullAdder U99 (w780, w679, IN49[2], w781, w782);
  FullAdder U100 (w782, w681, IN50[2], w783, w784);
  FullAdder U101 (w784, w683, IN51[2], w785, w786);
  FullAdder U102 (w786, w685, IN52[2], w787, w788);
  FullAdder U103 (w788, w686, IN53[0], w789, w790);
  HalfAdder U104 (w689, IN3[3], Out1[3], w792);
  FullAdder U105 (w792, w691, IN4[3], w793, w794);
  FullAdder U106 (w794, w693, IN5[3], w795, w796);
  FullAdder U107 (w796, w695, IN6[3], w797, w798);
  FullAdder U108 (w798, w697, IN7[3], w799, w800);
  FullAdder U109 (w800, w699, IN8[3], w801, w802);
  FullAdder U110 (w802, w701, IN9[3], w803, w804);
  FullAdder U111 (w804, w703, IN10[3], w805, w806);
  FullAdder U112 (w806, w705, IN11[3], w807, w808);
  FullAdder U113 (w808, w707, IN12[3], w809, w810);
  FullAdder U114 (w810, w709, IN13[3], w811, w812);
  FullAdder U115 (w812, w711, IN14[3], w813, w814);
  FullAdder U116 (w814, w713, IN15[3], w815, w816);
  FullAdder U117 (w816, w715, IN16[3], w817, w818);
  FullAdder U118 (w818, w717, IN17[3], w819, w820);
  FullAdder U119 (w820, w719, IN18[3], w821, w822);
  FullAdder U120 (w822, w721, IN19[3], w823, w824);
  FullAdder U121 (w824, w723, IN20[3], w825, w826);
  FullAdder U122 (w826, w725, IN21[3], w827, w828);
  FullAdder U123 (w828, w727, IN22[3], w829, w830);
  FullAdder U124 (w830, w729, IN23[3], w831, w832);
  FullAdder U125 (w832, w731, IN24[3], w833, w834);
  FullAdder U126 (w834, w733, IN25[3], w835, w836);
  FullAdder U127 (w836, w735, IN26[3], w837, w838);
  FullAdder U128 (w838, w737, IN27[3], w839, w840);
  FullAdder U129 (w840, w739, IN28[3], w841, w842);
  FullAdder U130 (w842, w741, IN29[3], w843, w844);
  FullAdder U131 (w844, w743, IN30[3], w845, w846);
  FullAdder U132 (w846, w745, IN31[3], w847, w848);
  FullAdder U133 (w848, w747, IN32[3], w849, w850);
  FullAdder U134 (w850, w749, IN33[3], w851, w852);
  FullAdder U135 (w852, w751, IN34[3], w853, w854);
  FullAdder U136 (w854, w753, IN35[3], w855, w856);
  FullAdder U137 (w856, w755, IN36[3], w857, w858);
  FullAdder U138 (w858, w757, IN37[3], w859, w860);
  FullAdder U139 (w860, w759, IN38[3], w861, w862);
  FullAdder U140 (w862, w761, IN39[3], w863, w864);
  FullAdder U141 (w864, w763, IN40[3], w865, w866);
  FullAdder U142 (w866, w765, IN41[3], w867, w868);
  FullAdder U143 (w868, w767, IN42[3], w869, w870);
  FullAdder U144 (w870, w769, IN43[3], w871, w872);
  FullAdder U145 (w872, w771, IN44[3], w873, w874);
  FullAdder U146 (w874, w773, IN45[3], w875, w876);
  FullAdder U147 (w876, w775, IN46[3], w877, w878);
  FullAdder U148 (w878, w777, IN47[3], w879, w880);
  FullAdder U149 (w880, w779, IN48[3], w881, w882);
  FullAdder U150 (w882, w781, IN49[3], w883, w884);
  FullAdder U151 (w884, w783, IN50[3], w885, w886);
  FullAdder U152 (w886, w785, IN51[3], w887, w888);
  FullAdder U153 (w888, w787, IN52[3], w889, w890);
  FullAdder U154 (w890, w789, IN53[1], w891, w892);
  FullAdder U155 (w892, w790, IN54[0], w893, w894);
  HalfAdder U156 (w793, IN4[4], Out1[4], w896);
  FullAdder U157 (w896, w795, IN5[4], w897, w898);
  FullAdder U158 (w898, w797, IN6[4], w899, w900);
  FullAdder U159 (w900, w799, IN7[4], w901, w902);
  FullAdder U160 (w902, w801, IN8[4], w903, w904);
  FullAdder U161 (w904, w803, IN9[4], w905, w906);
  FullAdder U162 (w906, w805, IN10[4], w907, w908);
  FullAdder U163 (w908, w807, IN11[4], w909, w910);
  FullAdder U164 (w910, w809, IN12[4], w911, w912);
  FullAdder U165 (w912, w811, IN13[4], w913, w914);
  FullAdder U166 (w914, w813, IN14[4], w915, w916);
  FullAdder U167 (w916, w815, IN15[4], w917, w918);
  FullAdder U168 (w918, w817, IN16[4], w919, w920);
  FullAdder U169 (w920, w819, IN17[4], w921, w922);
  FullAdder U170 (w922, w821, IN18[4], w923, w924);
  FullAdder U171 (w924, w823, IN19[4], w925, w926);
  FullAdder U172 (w926, w825, IN20[4], w927, w928);
  FullAdder U173 (w928, w827, IN21[4], w929, w930);
  FullAdder U174 (w930, w829, IN22[4], w931, w932);
  FullAdder U175 (w932, w831, IN23[4], w933, w934);
  FullAdder U176 (w934, w833, IN24[4], w935, w936);
  FullAdder U177 (w936, w835, IN25[4], w937, w938);
  FullAdder U178 (w938, w837, IN26[4], w939, w940);
  FullAdder U179 (w940, w839, IN27[4], w941, w942);
  FullAdder U180 (w942, w841, IN28[4], w943, w944);
  FullAdder U181 (w944, w843, IN29[4], w945, w946);
  FullAdder U182 (w946, w845, IN30[4], w947, w948);
  FullAdder U183 (w948, w847, IN31[4], w949, w950);
  FullAdder U184 (w950, w849, IN32[4], w951, w952);
  FullAdder U185 (w952, w851, IN33[4], w953, w954);
  FullAdder U186 (w954, w853, IN34[4], w955, w956);
  FullAdder U187 (w956, w855, IN35[4], w957, w958);
  FullAdder U188 (w958, w857, IN36[4], w959, w960);
  FullAdder U189 (w960, w859, IN37[4], w961, w962);
  FullAdder U190 (w962, w861, IN38[4], w963, w964);
  FullAdder U191 (w964, w863, IN39[4], w965, w966);
  FullAdder U192 (w966, w865, IN40[4], w967, w968);
  FullAdder U193 (w968, w867, IN41[4], w969, w970);
  FullAdder U194 (w970, w869, IN42[4], w971, w972);
  FullAdder U195 (w972, w871, IN43[4], w973, w974);
  FullAdder U196 (w974, w873, IN44[4], w975, w976);
  FullAdder U197 (w976, w875, IN45[4], w977, w978);
  FullAdder U198 (w978, w877, IN46[4], w979, w980);
  FullAdder U199 (w980, w879, IN47[4], w981, w982);
  FullAdder U200 (w982, w881, IN48[4], w983, w984);
  FullAdder U201 (w984, w883, IN49[4], w985, w986);
  FullAdder U202 (w986, w885, IN50[4], w987, w988);
  FullAdder U203 (w988, w887, IN51[4], w989, w990);
  FullAdder U204 (w990, w889, IN52[4], w991, w992);
  FullAdder U205 (w992, w891, IN53[2], w993, w994);
  FullAdder U206 (w994, w893, IN54[1], w995, w996);
  FullAdder U207 (w996, w894, IN55[0], w997, w998);
  HalfAdder U208 (w897, IN5[5], Out1[5], w1000);
  FullAdder U209 (w1000, w899, IN6[5], w1001, w1002);
  FullAdder U210 (w1002, w901, IN7[5], w1003, w1004);
  FullAdder U211 (w1004, w903, IN8[5], w1005, w1006);
  FullAdder U212 (w1006, w905, IN9[5], w1007, w1008);
  FullAdder U213 (w1008, w907, IN10[5], w1009, w1010);
  FullAdder U214 (w1010, w909, IN11[5], w1011, w1012);
  FullAdder U215 (w1012, w911, IN12[5], w1013, w1014);
  FullAdder U216 (w1014, w913, IN13[5], w1015, w1016);
  FullAdder U217 (w1016, w915, IN14[5], w1017, w1018);
  FullAdder U218 (w1018, w917, IN15[5], w1019, w1020);
  FullAdder U219 (w1020, w919, IN16[5], w1021, w1022);
  FullAdder U220 (w1022, w921, IN17[5], w1023, w1024);
  FullAdder U221 (w1024, w923, IN18[5], w1025, w1026);
  FullAdder U222 (w1026, w925, IN19[5], w1027, w1028);
  FullAdder U223 (w1028, w927, IN20[5], w1029, w1030);
  FullAdder U224 (w1030, w929, IN21[5], w1031, w1032);
  FullAdder U225 (w1032, w931, IN22[5], w1033, w1034);
  FullAdder U226 (w1034, w933, IN23[5], w1035, w1036);
  FullAdder U227 (w1036, w935, IN24[5], w1037, w1038);
  FullAdder U228 (w1038, w937, IN25[5], w1039, w1040);
  FullAdder U229 (w1040, w939, IN26[5], w1041, w1042);
  FullAdder U230 (w1042, w941, IN27[5], w1043, w1044);
  FullAdder U231 (w1044, w943, IN28[5], w1045, w1046);
  FullAdder U232 (w1046, w945, IN29[5], w1047, w1048);
  FullAdder U233 (w1048, w947, IN30[5], w1049, w1050);
  FullAdder U234 (w1050, w949, IN31[5], w1051, w1052);
  FullAdder U235 (w1052, w951, IN32[5], w1053, w1054);
  FullAdder U236 (w1054, w953, IN33[5], w1055, w1056);
  FullAdder U237 (w1056, w955, IN34[5], w1057, w1058);
  FullAdder U238 (w1058, w957, IN35[5], w1059, w1060);
  FullAdder U239 (w1060, w959, IN36[5], w1061, w1062);
  FullAdder U240 (w1062, w961, IN37[5], w1063, w1064);
  FullAdder U241 (w1064, w963, IN38[5], w1065, w1066);
  FullAdder U242 (w1066, w965, IN39[5], w1067, w1068);
  FullAdder U243 (w1068, w967, IN40[5], w1069, w1070);
  FullAdder U244 (w1070, w969, IN41[5], w1071, w1072);
  FullAdder U245 (w1072, w971, IN42[5], w1073, w1074);
  FullAdder U246 (w1074, w973, IN43[5], w1075, w1076);
  FullAdder U247 (w1076, w975, IN44[5], w1077, w1078);
  FullAdder U248 (w1078, w977, IN45[5], w1079, w1080);
  FullAdder U249 (w1080, w979, IN46[5], w1081, w1082);
  FullAdder U250 (w1082, w981, IN47[5], w1083, w1084);
  FullAdder U251 (w1084, w983, IN48[5], w1085, w1086);
  FullAdder U252 (w1086, w985, IN49[5], w1087, w1088);
  FullAdder U253 (w1088, w987, IN50[5], w1089, w1090);
  FullAdder U254 (w1090, w989, IN51[5], w1091, w1092);
  FullAdder U255 (w1092, w991, IN52[5], w1093, w1094);
  FullAdder U256 (w1094, w993, IN53[3], w1095, w1096);
  FullAdder U257 (w1096, w995, IN54[2], w1097, w1098);
  FullAdder U258 (w1098, w997, IN55[1], w1099, w1100);
  FullAdder U259 (w1100, w998, IN56[0], w1101, w1102);
  HalfAdder U260 (w1001, IN6[6], Out1[6], w1104);
  FullAdder U261 (w1104, w1003, IN7[6], w1105, w1106);
  FullAdder U262 (w1106, w1005, IN8[6], w1107, w1108);
  FullAdder U263 (w1108, w1007, IN9[6], w1109, w1110);
  FullAdder U264 (w1110, w1009, IN10[6], w1111, w1112);
  FullAdder U265 (w1112, w1011, IN11[6], w1113, w1114);
  FullAdder U266 (w1114, w1013, IN12[6], w1115, w1116);
  FullAdder U267 (w1116, w1015, IN13[6], w1117, w1118);
  FullAdder U268 (w1118, w1017, IN14[6], w1119, w1120);
  FullAdder U269 (w1120, w1019, IN15[6], w1121, w1122);
  FullAdder U270 (w1122, w1021, IN16[6], w1123, w1124);
  FullAdder U271 (w1124, w1023, IN17[6], w1125, w1126);
  FullAdder U272 (w1126, w1025, IN18[6], w1127, w1128);
  FullAdder U273 (w1128, w1027, IN19[6], w1129, w1130);
  FullAdder U274 (w1130, w1029, IN20[6], w1131, w1132);
  FullAdder U275 (w1132, w1031, IN21[6], w1133, w1134);
  FullAdder U276 (w1134, w1033, IN22[6], w1135, w1136);
  FullAdder U277 (w1136, w1035, IN23[6], w1137, w1138);
  FullAdder U278 (w1138, w1037, IN24[6], w1139, w1140);
  FullAdder U279 (w1140, w1039, IN25[6], w1141, w1142);
  FullAdder U280 (w1142, w1041, IN26[6], w1143, w1144);
  FullAdder U281 (w1144, w1043, IN27[6], w1145, w1146);
  FullAdder U282 (w1146, w1045, IN28[6], w1147, w1148);
  FullAdder U283 (w1148, w1047, IN29[6], w1149, w1150);
  FullAdder U284 (w1150, w1049, IN30[6], w1151, w1152);
  FullAdder U285 (w1152, w1051, IN31[6], w1153, w1154);
  FullAdder U286 (w1154, w1053, IN32[6], w1155, w1156);
  FullAdder U287 (w1156, w1055, IN33[6], w1157, w1158);
  FullAdder U288 (w1158, w1057, IN34[6], w1159, w1160);
  FullAdder U289 (w1160, w1059, IN35[6], w1161, w1162);
  FullAdder U290 (w1162, w1061, IN36[6], w1163, w1164);
  FullAdder U291 (w1164, w1063, IN37[6], w1165, w1166);
  FullAdder U292 (w1166, w1065, IN38[6], w1167, w1168);
  FullAdder U293 (w1168, w1067, IN39[6], w1169, w1170);
  FullAdder U294 (w1170, w1069, IN40[6], w1171, w1172);
  FullAdder U295 (w1172, w1071, IN41[6], w1173, w1174);
  FullAdder U296 (w1174, w1073, IN42[6], w1175, w1176);
  FullAdder U297 (w1176, w1075, IN43[6], w1177, w1178);
  FullAdder U298 (w1178, w1077, IN44[6], w1179, w1180);
  FullAdder U299 (w1180, w1079, IN45[6], w1181, w1182);
  FullAdder U300 (w1182, w1081, IN46[6], w1183, w1184);
  FullAdder U301 (w1184, w1083, IN47[6], w1185, w1186);
  FullAdder U302 (w1186, w1085, IN48[6], w1187, w1188);
  FullAdder U303 (w1188, w1087, IN49[6], w1189, w1190);
  FullAdder U304 (w1190, w1089, IN50[6], w1191, w1192);
  FullAdder U305 (w1192, w1091, IN51[6], w1193, w1194);
  FullAdder U306 (w1194, w1093, IN52[6], w1195, w1196);
  FullAdder U307 (w1196, w1095, IN53[4], w1197, w1198);
  FullAdder U308 (w1198, w1097, IN54[3], w1199, w1200);
  FullAdder U309 (w1200, w1099, IN55[2], w1201, w1202);
  FullAdder U310 (w1202, w1101, IN56[1], w1203, w1204);
  FullAdder U311 (w1204, w1102, IN57[0], w1205, w1206);
  HalfAdder U312 (w1105, IN7[7], Out1[7], w1208);
  FullAdder U313 (w1208, w1107, IN8[7], w1209, w1210);
  FullAdder U314 (w1210, w1109, IN9[7], w1211, w1212);
  FullAdder U315 (w1212, w1111, IN10[7], w1213, w1214);
  FullAdder U316 (w1214, w1113, IN11[7], w1215, w1216);
  FullAdder U317 (w1216, w1115, IN12[7], w1217, w1218);
  FullAdder U318 (w1218, w1117, IN13[7], w1219, w1220);
  FullAdder U319 (w1220, w1119, IN14[7], w1221, w1222);
  FullAdder U320 (w1222, w1121, IN15[7], w1223, w1224);
  FullAdder U321 (w1224, w1123, IN16[7], w1225, w1226);
  FullAdder U322 (w1226, w1125, IN17[7], w1227, w1228);
  FullAdder U323 (w1228, w1127, IN18[7], w1229, w1230);
  FullAdder U324 (w1230, w1129, IN19[7], w1231, w1232);
  FullAdder U325 (w1232, w1131, IN20[7], w1233, w1234);
  FullAdder U326 (w1234, w1133, IN21[7], w1235, w1236);
  FullAdder U327 (w1236, w1135, IN22[7], w1237, w1238);
  FullAdder U328 (w1238, w1137, IN23[7], w1239, w1240);
  FullAdder U329 (w1240, w1139, IN24[7], w1241, w1242);
  FullAdder U330 (w1242, w1141, IN25[7], w1243, w1244);
  FullAdder U331 (w1244, w1143, IN26[7], w1245, w1246);
  FullAdder U332 (w1246, w1145, IN27[7], w1247, w1248);
  FullAdder U333 (w1248, w1147, IN28[7], w1249, w1250);
  FullAdder U334 (w1250, w1149, IN29[7], w1251, w1252);
  FullAdder U335 (w1252, w1151, IN30[7], w1253, w1254);
  FullAdder U336 (w1254, w1153, IN31[7], w1255, w1256);
  FullAdder U337 (w1256, w1155, IN32[7], w1257, w1258);
  FullAdder U338 (w1258, w1157, IN33[7], w1259, w1260);
  FullAdder U339 (w1260, w1159, IN34[7], w1261, w1262);
  FullAdder U340 (w1262, w1161, IN35[7], w1263, w1264);
  FullAdder U341 (w1264, w1163, IN36[7], w1265, w1266);
  FullAdder U342 (w1266, w1165, IN37[7], w1267, w1268);
  FullAdder U343 (w1268, w1167, IN38[7], w1269, w1270);
  FullAdder U344 (w1270, w1169, IN39[7], w1271, w1272);
  FullAdder U345 (w1272, w1171, IN40[7], w1273, w1274);
  FullAdder U346 (w1274, w1173, IN41[7], w1275, w1276);
  FullAdder U347 (w1276, w1175, IN42[7], w1277, w1278);
  FullAdder U348 (w1278, w1177, IN43[7], w1279, w1280);
  FullAdder U349 (w1280, w1179, IN44[7], w1281, w1282);
  FullAdder U350 (w1282, w1181, IN45[7], w1283, w1284);
  FullAdder U351 (w1284, w1183, IN46[7], w1285, w1286);
  FullAdder U352 (w1286, w1185, IN47[7], w1287, w1288);
  FullAdder U353 (w1288, w1187, IN48[7], w1289, w1290);
  FullAdder U354 (w1290, w1189, IN49[7], w1291, w1292);
  FullAdder U355 (w1292, w1191, IN50[7], w1293, w1294);
  FullAdder U356 (w1294, w1193, IN51[7], w1295, w1296);
  FullAdder U357 (w1296, w1195, IN52[7], w1297, w1298);
  FullAdder U358 (w1298, w1197, IN53[5], w1299, w1300);
  FullAdder U359 (w1300, w1199, IN54[4], w1301, w1302);
  FullAdder U360 (w1302, w1201, IN55[3], w1303, w1304);
  FullAdder U361 (w1304, w1203, IN56[2], w1305, w1306);
  FullAdder U362 (w1306, w1205, IN57[1], w1307, w1308);
  FullAdder U363 (w1308, w1206, IN58[0], w1309, w1310);
  HalfAdder U364 (w1209, IN8[8], Out1[8], w1312);
  FullAdder U365 (w1312, w1211, IN9[8], w1313, w1314);
  FullAdder U366 (w1314, w1213, IN10[8], w1315, w1316);
  FullAdder U367 (w1316, w1215, IN11[8], w1317, w1318);
  FullAdder U368 (w1318, w1217, IN12[8], w1319, w1320);
  FullAdder U369 (w1320, w1219, IN13[8], w1321, w1322);
  FullAdder U370 (w1322, w1221, IN14[8], w1323, w1324);
  FullAdder U371 (w1324, w1223, IN15[8], w1325, w1326);
  FullAdder U372 (w1326, w1225, IN16[8], w1327, w1328);
  FullAdder U373 (w1328, w1227, IN17[8], w1329, w1330);
  FullAdder U374 (w1330, w1229, IN18[8], w1331, w1332);
  FullAdder U375 (w1332, w1231, IN19[8], w1333, w1334);
  FullAdder U376 (w1334, w1233, IN20[8], w1335, w1336);
  FullAdder U377 (w1336, w1235, IN21[8], w1337, w1338);
  FullAdder U378 (w1338, w1237, IN22[8], w1339, w1340);
  FullAdder U379 (w1340, w1239, IN23[8], w1341, w1342);
  FullAdder U380 (w1342, w1241, IN24[8], w1343, w1344);
  FullAdder U381 (w1344, w1243, IN25[8], w1345, w1346);
  FullAdder U382 (w1346, w1245, IN26[8], w1347, w1348);
  FullAdder U383 (w1348, w1247, IN27[8], w1349, w1350);
  FullAdder U384 (w1350, w1249, IN28[8], w1351, w1352);
  FullAdder U385 (w1352, w1251, IN29[8], w1353, w1354);
  FullAdder U386 (w1354, w1253, IN30[8], w1355, w1356);
  FullAdder U387 (w1356, w1255, IN31[8], w1357, w1358);
  FullAdder U388 (w1358, w1257, IN32[8], w1359, w1360);
  FullAdder U389 (w1360, w1259, IN33[8], w1361, w1362);
  FullAdder U390 (w1362, w1261, IN34[8], w1363, w1364);
  FullAdder U391 (w1364, w1263, IN35[8], w1365, w1366);
  FullAdder U392 (w1366, w1265, IN36[8], w1367, w1368);
  FullAdder U393 (w1368, w1267, IN37[8], w1369, w1370);
  FullAdder U394 (w1370, w1269, IN38[8], w1371, w1372);
  FullAdder U395 (w1372, w1271, IN39[8], w1373, w1374);
  FullAdder U396 (w1374, w1273, IN40[8], w1375, w1376);
  FullAdder U397 (w1376, w1275, IN41[8], w1377, w1378);
  FullAdder U398 (w1378, w1277, IN42[8], w1379, w1380);
  FullAdder U399 (w1380, w1279, IN43[8], w1381, w1382);
  FullAdder U400 (w1382, w1281, IN44[8], w1383, w1384);
  FullAdder U401 (w1384, w1283, IN45[8], w1385, w1386);
  FullAdder U402 (w1386, w1285, IN46[8], w1387, w1388);
  FullAdder U403 (w1388, w1287, IN47[8], w1389, w1390);
  FullAdder U404 (w1390, w1289, IN48[8], w1391, w1392);
  FullAdder U405 (w1392, w1291, IN49[8], w1393, w1394);
  FullAdder U406 (w1394, w1293, IN50[8], w1395, w1396);
  FullAdder U407 (w1396, w1295, IN51[8], w1397, w1398);
  FullAdder U408 (w1398, w1297, IN52[8], w1399, w1400);
  FullAdder U409 (w1400, w1299, IN53[6], w1401, w1402);
  FullAdder U410 (w1402, w1301, IN54[5], w1403, w1404);
  FullAdder U411 (w1404, w1303, IN55[4], w1405, w1406);
  FullAdder U412 (w1406, w1305, IN56[3], w1407, w1408);
  FullAdder U413 (w1408, w1307, IN57[2], w1409, w1410);
  FullAdder U414 (w1410, w1309, IN58[1], w1411, w1412);
  FullAdder U415 (w1412, w1310, IN59[0], w1413, w1414);
  HalfAdder U416 (w1313, IN9[9], Out1[9], w1416);
  FullAdder U417 (w1416, w1315, IN10[9], w1417, w1418);
  FullAdder U418 (w1418, w1317, IN11[9], w1419, w1420);
  FullAdder U419 (w1420, w1319, IN12[9], w1421, w1422);
  FullAdder U420 (w1422, w1321, IN13[9], w1423, w1424);
  FullAdder U421 (w1424, w1323, IN14[9], w1425, w1426);
  FullAdder U422 (w1426, w1325, IN15[9], w1427, w1428);
  FullAdder U423 (w1428, w1327, IN16[9], w1429, w1430);
  FullAdder U424 (w1430, w1329, IN17[9], w1431, w1432);
  FullAdder U425 (w1432, w1331, IN18[9], w1433, w1434);
  FullAdder U426 (w1434, w1333, IN19[9], w1435, w1436);
  FullAdder U427 (w1436, w1335, IN20[9], w1437, w1438);
  FullAdder U428 (w1438, w1337, IN21[9], w1439, w1440);
  FullAdder U429 (w1440, w1339, IN22[9], w1441, w1442);
  FullAdder U430 (w1442, w1341, IN23[9], w1443, w1444);
  FullAdder U431 (w1444, w1343, IN24[9], w1445, w1446);
  FullAdder U432 (w1446, w1345, IN25[9], w1447, w1448);
  FullAdder U433 (w1448, w1347, IN26[9], w1449, w1450);
  FullAdder U434 (w1450, w1349, IN27[9], w1451, w1452);
  FullAdder U435 (w1452, w1351, IN28[9], w1453, w1454);
  FullAdder U436 (w1454, w1353, IN29[9], w1455, w1456);
  FullAdder U437 (w1456, w1355, IN30[9], w1457, w1458);
  FullAdder U438 (w1458, w1357, IN31[9], w1459, w1460);
  FullAdder U439 (w1460, w1359, IN32[9], w1461, w1462);
  FullAdder U440 (w1462, w1361, IN33[9], w1463, w1464);
  FullAdder U441 (w1464, w1363, IN34[9], w1465, w1466);
  FullAdder U442 (w1466, w1365, IN35[9], w1467, w1468);
  FullAdder U443 (w1468, w1367, IN36[9], w1469, w1470);
  FullAdder U444 (w1470, w1369, IN37[9], w1471, w1472);
  FullAdder U445 (w1472, w1371, IN38[9], w1473, w1474);
  FullAdder U446 (w1474, w1373, IN39[9], w1475, w1476);
  FullAdder U447 (w1476, w1375, IN40[9], w1477, w1478);
  FullAdder U448 (w1478, w1377, IN41[9], w1479, w1480);
  FullAdder U449 (w1480, w1379, IN42[9], w1481, w1482);
  FullAdder U450 (w1482, w1381, IN43[9], w1483, w1484);
  FullAdder U451 (w1484, w1383, IN44[9], w1485, w1486);
  FullAdder U452 (w1486, w1385, IN45[9], w1487, w1488);
  FullAdder U453 (w1488, w1387, IN46[9], w1489, w1490);
  FullAdder U454 (w1490, w1389, IN47[9], w1491, w1492);
  FullAdder U455 (w1492, w1391, IN48[9], w1493, w1494);
  FullAdder U456 (w1494, w1393, IN49[9], w1495, w1496);
  FullAdder U457 (w1496, w1395, IN50[9], w1497, w1498);
  FullAdder U458 (w1498, w1397, IN51[9], w1499, w1500);
  FullAdder U459 (w1500, w1399, IN52[9], w1501, w1502);
  FullAdder U460 (w1502, w1401, IN53[7], w1503, w1504);
  FullAdder U461 (w1504, w1403, IN54[6], w1505, w1506);
  FullAdder U462 (w1506, w1405, IN55[5], w1507, w1508);
  FullAdder U463 (w1508, w1407, IN56[4], w1509, w1510);
  FullAdder U464 (w1510, w1409, IN57[3], w1511, w1512);
  FullAdder U465 (w1512, w1411, IN58[2], w1513, w1514);
  FullAdder U466 (w1514, w1413, IN59[1], w1515, w1516);
  FullAdder U467 (w1516, w1414, IN60[0], w1517, w1518);
  HalfAdder U468 (w1417, IN10[10], Out1[10], w1520);
  FullAdder U469 (w1520, w1419, IN11[10], Out1[11], w1522);
  FullAdder U470 (w1522, w1421, IN12[10], Out1[12], w1524);
  FullAdder U471 (w1524, w1423, IN13[10], Out1[13], w1526);
  FullAdder U472 (w1526, w1425, IN14[10], Out1[14], w1528);
  FullAdder U473 (w1528, w1427, IN15[10], Out1[15], w1530);
  FullAdder U474 (w1530, w1429, IN16[10], Out1[16], w1532);
  FullAdder U475 (w1532, w1431, IN17[10], Out1[17], w1534);
  FullAdder U476 (w1534, w1433, IN18[10], Out1[18], w1536);
  FullAdder U477 (w1536, w1435, IN19[10], Out1[19], w1538);
  FullAdder U478 (w1538, w1437, IN20[10], Out1[20], w1540);
  FullAdder U479 (w1540, w1439, IN21[10], Out1[21], w1542);
  FullAdder U480 (w1542, w1441, IN22[10], Out1[22], w1544);
  FullAdder U481 (w1544, w1443, IN23[10], Out1[23], w1546);
  FullAdder U482 (w1546, w1445, IN24[10], Out1[24], w1548);
  FullAdder U483 (w1548, w1447, IN25[10], Out1[25], w1550);
  FullAdder U484 (w1550, w1449, IN26[10], Out1[26], w1552);
  FullAdder U485 (w1552, w1451, IN27[10], Out1[27], w1554);
  FullAdder U486 (w1554, w1453, IN28[10], Out1[28], w1556);
  FullAdder U487 (w1556, w1455, IN29[10], Out1[29], w1558);
  FullAdder U488 (w1558, w1457, IN30[10], Out1[30], w1560);
  FullAdder U489 (w1560, w1459, IN31[10], Out1[31], w1562);
  FullAdder U490 (w1562, w1461, IN32[10], Out1[32], w1564);
  FullAdder U491 (w1564, w1463, IN33[10], Out1[33], w1566);
  FullAdder U492 (w1566, w1465, IN34[10], Out1[34], w1568);
  FullAdder U493 (w1568, w1467, IN35[10], Out1[35], w1570);
  FullAdder U494 (w1570, w1469, IN36[10], Out1[36], w1572);
  FullAdder U495 (w1572, w1471, IN37[10], Out1[37], w1574);
  FullAdder U496 (w1574, w1473, IN38[10], Out1[38], w1576);
  FullAdder U497 (w1576, w1475, IN39[10], Out1[39], w1578);
  FullAdder U498 (w1578, w1477, IN40[10], Out1[40], w1580);
  FullAdder U499 (w1580, w1479, IN41[10], Out1[41], w1582);
  FullAdder U500 (w1582, w1481, IN42[10], Out1[42], w1584);
  FullAdder U501 (w1584, w1483, IN43[10], Out1[43], w1586);
  FullAdder U502 (w1586, w1485, IN44[10], Out1[44], w1588);
  FullAdder U503 (w1588, w1487, IN45[10], Out1[45], w1590);
  FullAdder U504 (w1590, w1489, IN46[10], Out1[46], w1592);
  FullAdder U505 (w1592, w1491, IN47[10], Out1[47], w1594);
  FullAdder U506 (w1594, w1493, IN48[10], Out1[48], w1596);
  FullAdder U507 (w1596, w1495, IN49[10], Out1[49], w1598);
  FullAdder U508 (w1598, w1497, IN50[10], Out1[50], w1600);
  FullAdder U509 (w1600, w1499, IN51[10], Out1[51], w1602);
  FullAdder U510 (w1602, w1501, IN52[10], Out1[52], w1604);
  FullAdder U511 (w1604, w1503, IN53[8], Out1[53], w1606);
  FullAdder U512 (w1606, w1505, IN54[7], Out1[54], w1608);
  FullAdder U513 (w1608, w1507, IN55[6], Out1[55], w1610);
  FullAdder U514 (w1610, w1509, IN56[5], Out1[56], w1612);
  FullAdder U515 (w1612, w1511, IN57[4], Out1[57], w1614);
  FullAdder U516 (w1614, w1513, IN58[3], Out1[58], w1616);
  FullAdder U517 (w1616, w1515, IN59[2], Out1[59], w1618);
  FullAdder U518 (w1618, w1517, IN60[1], Out1[60], w1620);
  FullAdder U519 (w1620, w1518, IN61[0], Out1[61], Out1[62]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN53[9];
  assign Out2[1] = IN54[8];
  assign Out2[2] = IN55[7];
  assign Out2[3] = IN56[6];
  assign Out2[4] = IN57[5];
  assign Out2[5] = IN58[4];
  assign Out2[6] = IN59[3];
  assign Out2[7] = IN60[2];
  assign Out2[8] = IN61[1];
  assign Out2[9] = IN62[0];

endmodule
module RC_10_10(IN1, IN2, Out);
  input [9:0] IN1;
  input [9:0] IN2;
  output [10:0] Out;
  wire w21;
  wire w23;
  wire w25;
  wire w27;
  wire w29;
  wire w31;
  wire w33;
  wire w35;
  wire w37;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w21);
  FullAdder U1 (IN1[1], IN2[1], w21, Out[1], w23);
  FullAdder U2 (IN1[2], IN2[2], w23, Out[2], w25);
  FullAdder U3 (IN1[3], IN2[3], w25, Out[3], w27);
  FullAdder U4 (IN1[4], IN2[4], w27, Out[4], w29);
  FullAdder U5 (IN1[5], IN2[5], w29, Out[5], w31);
  FullAdder U6 (IN1[6], IN2[6], w31, Out[6], w33);
  FullAdder U7 (IN1[7], IN2[7], w33, Out[7], w35);
  FullAdder U8 (IN1[8], IN2[8], w35, Out[8], w37);
  FullAdder U9 (IN1[9], IN2[9], w37, Out[9], Out[10]);

endmodule
module NR_53_11(IN1, IN2, Out);
  input [52:0] IN1;
  input [10:0] IN2;
  output [63:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [10:0] P11;
  wire [10:0] P12;
  wire [10:0] P13;
  wire [10:0] P14;
  wire [10:0] P15;
  wire [10:0] P16;
  wire [10:0] P17;
  wire [10:0] P18;
  wire [10:0] P19;
  wire [10:0] P20;
  wire [10:0] P21;
  wire [10:0] P22;
  wire [10:0] P23;
  wire [10:0] P24;
  wire [10:0] P25;
  wire [10:0] P26;
  wire [10:0] P27;
  wire [10:0] P28;
  wire [10:0] P29;
  wire [10:0] P30;
  wire [10:0] P31;
  wire [10:0] P32;
  wire [10:0] P33;
  wire [10:0] P34;
  wire [10:0] P35;
  wire [10:0] P36;
  wire [10:0] P37;
  wire [10:0] P38;
  wire [10:0] P39;
  wire [10:0] P40;
  wire [10:0] P41;
  wire [10:0] P42;
  wire [10:0] P43;
  wire [10:0] P44;
  wire [10:0] P45;
  wire [10:0] P46;
  wire [10:0] P47;
  wire [10:0] P48;
  wire [10:0] P49;
  wire [10:0] P50;
  wire [10:0] P51;
  wire [10:0] P52;
  wire [9:0] P53;
  wire [8:0] P54;
  wire [7:0] P55;
  wire [6:0] P56;
  wire [5:0] P57;
  wire [4:0] P58;
  wire [3:0] P59;
  wire [2:0] P60;
  wire [1:0] P61;
  wire [0:0] P62;
  wire [62:0] R1;
  wire [9:0] R2;
  wire [63:0] aOut;
  U_SP_53_11 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, R1, R2);
  RC_10_10 S2 (R1[62:53], R2, aOut[63:53]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign Out = aOut[63:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
