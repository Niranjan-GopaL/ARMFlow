
module NR_35_1(
    input [34:0]IN1,
    input [0:0]IN2,
    output [34:0]Out
);
    assign Out = IN2;
endmodule
