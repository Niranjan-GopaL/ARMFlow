//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 9
  second input length: 44
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_9_44(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51);
  input [8:0] IN1;
  input [43:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [8:0] P9;
  output [8:0] P10;
  output [8:0] P11;
  output [8:0] P12;
  output [8:0] P13;
  output [8:0] P14;
  output [8:0] P15;
  output [8:0] P16;
  output [8:0] P17;
  output [8:0] P18;
  output [8:0] P19;
  output [8:0] P20;
  output [8:0] P21;
  output [8:0] P22;
  output [8:0] P23;
  output [8:0] P24;
  output [8:0] P25;
  output [8:0] P26;
  output [8:0] P27;
  output [8:0] P28;
  output [8:0] P29;
  output [8:0] P30;
  output [8:0] P31;
  output [8:0] P32;
  output [8:0] P33;
  output [8:0] P34;
  output [8:0] P35;
  output [8:0] P36;
  output [8:0] P37;
  output [8:0] P38;
  output [8:0] P39;
  output [8:0] P40;
  output [8:0] P41;
  output [8:0] P42;
  output [8:0] P43;
  output [7:0] P44;
  output [6:0] P45;
  output [5:0] P46;
  output [4:0] P47;
  output [3:0] P48;
  output [2:0] P49;
  output [1:0] P50;
  output [0:0] P51;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[0] = IN1[1]&IN2[43];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[1] = IN1[2]&IN2[42];
  assign P45[0] = IN1[2]&IN2[43];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[2] = IN1[3]&IN2[41];
  assign P45[1] = IN1[3]&IN2[42];
  assign P46[0] = IN1[3]&IN2[43];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[3] = IN1[4]&IN2[40];
  assign P45[2] = IN1[4]&IN2[41];
  assign P46[1] = IN1[4]&IN2[42];
  assign P47[0] = IN1[4]&IN2[43];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[4] = IN1[5]&IN2[39];
  assign P45[3] = IN1[5]&IN2[40];
  assign P46[2] = IN1[5]&IN2[41];
  assign P47[1] = IN1[5]&IN2[42];
  assign P48[0] = IN1[5]&IN2[43];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[5] = IN1[6]&IN2[38];
  assign P45[4] = IN1[6]&IN2[39];
  assign P46[3] = IN1[6]&IN2[40];
  assign P47[2] = IN1[6]&IN2[41];
  assign P48[1] = IN1[6]&IN2[42];
  assign P49[0] = IN1[6]&IN2[43];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[6] = IN1[7]&IN2[37];
  assign P45[5] = IN1[7]&IN2[38];
  assign P46[4] = IN1[7]&IN2[39];
  assign P47[3] = IN1[7]&IN2[40];
  assign P48[2] = IN1[7]&IN2[41];
  assign P49[1] = IN1[7]&IN2[42];
  assign P50[0] = IN1[7]&IN2[43];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[7] = IN1[8]&IN2[36];
  assign P45[6] = IN1[8]&IN2[37];
  assign P46[5] = IN1[8]&IN2[38];
  assign P47[4] = IN1[8]&IN2[39];
  assign P48[3] = IN1[8]&IN2[40];
  assign P49[2] = IN1[8]&IN2[41];
  assign P50[1] = IN1[8]&IN2[42];
  assign P51[0] = IN1[8]&IN2[43];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [8:0] IN9;
  input [8:0] IN10;
  input [8:0] IN11;
  input [8:0] IN12;
  input [8:0] IN13;
  input [8:0] IN14;
  input [8:0] IN15;
  input [8:0] IN16;
  input [8:0] IN17;
  input [8:0] IN18;
  input [8:0] IN19;
  input [8:0] IN20;
  input [8:0] IN21;
  input [8:0] IN22;
  input [8:0] IN23;
  input [8:0] IN24;
  input [8:0] IN25;
  input [8:0] IN26;
  input [8:0] IN27;
  input [8:0] IN28;
  input [8:0] IN29;
  input [8:0] IN30;
  input [8:0] IN31;
  input [8:0] IN32;
  input [8:0] IN33;
  input [8:0] IN34;
  input [8:0] IN35;
  input [8:0] IN36;
  input [8:0] IN37;
  input [8:0] IN38;
  input [8:0] IN39;
  input [8:0] IN40;
  input [8:0] IN41;
  input [8:0] IN42;
  input [8:0] IN43;
  input [7:0] IN44;
  input [6:0] IN45;
  input [5:0] IN46;
  input [4:0] IN47;
  input [3:0] IN48;
  input [2:0] IN49;
  input [1:0] IN50;
  input [0:0] IN51;
  output [51:0] Out1;
  output [42:0] Out2;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1069;
  wire w1071;
  wire w1073;
  wire w1075;
  wire w1077;
  wire w1079;
  wire w1081;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w397);
  FullAdder U1 (w397, IN2[0], IN2[1], w398, w399);
  FullAdder U2 (w399, IN3[0], IN3[1], w400, w401);
  FullAdder U3 (w401, IN4[0], IN4[1], w402, w403);
  FullAdder U4 (w403, IN5[0], IN5[1], w404, w405);
  FullAdder U5 (w405, IN6[0], IN6[1], w406, w407);
  FullAdder U6 (w407, IN7[0], IN7[1], w408, w409);
  FullAdder U7 (w409, IN8[0], IN8[1], w410, w411);
  HalfAdder U8 (w398, IN2[2], Out1[2], w413);
  FullAdder U9 (w413, w400, IN3[2], w414, w415);
  FullAdder U10 (w415, w402, IN4[2], w416, w417);
  FullAdder U11 (w417, w404, IN5[2], w418, w419);
  FullAdder U12 (w419, w406, IN6[2], w420, w421);
  FullAdder U13 (w421, w408, IN7[2], w422, w423);
  FullAdder U14 (w423, w410, IN8[2], w424, w425);
  FullAdder U15 (w425, w411, IN9[0], w426, w427);
  HalfAdder U16 (w414, IN3[3], Out1[3], w429);
  FullAdder U17 (w429, w416, IN4[3], w430, w431);
  FullAdder U18 (w431, w418, IN5[3], w432, w433);
  FullAdder U19 (w433, w420, IN6[3], w434, w435);
  FullAdder U20 (w435, w422, IN7[3], w436, w437);
  FullAdder U21 (w437, w424, IN8[3], w438, w439);
  FullAdder U22 (w439, w426, IN9[1], w440, w441);
  FullAdder U23 (w441, w427, IN10[0], w442, w443);
  HalfAdder U24 (w430, IN4[4], Out1[4], w445);
  FullAdder U25 (w445, w432, IN5[4], w446, w447);
  FullAdder U26 (w447, w434, IN6[4], w448, w449);
  FullAdder U27 (w449, w436, IN7[4], w450, w451);
  FullAdder U28 (w451, w438, IN8[4], w452, w453);
  FullAdder U29 (w453, w440, IN9[2], w454, w455);
  FullAdder U30 (w455, w442, IN10[1], w456, w457);
  FullAdder U31 (w457, w443, IN11[0], w458, w459);
  HalfAdder U32 (w446, IN5[5], Out1[5], w461);
  FullAdder U33 (w461, w448, IN6[5], w462, w463);
  FullAdder U34 (w463, w450, IN7[5], w464, w465);
  FullAdder U35 (w465, w452, IN8[5], w466, w467);
  FullAdder U36 (w467, w454, IN9[3], w468, w469);
  FullAdder U37 (w469, w456, IN10[2], w470, w471);
  FullAdder U38 (w471, w458, IN11[1], w472, w473);
  FullAdder U39 (w473, w459, IN12[0], w474, w475);
  HalfAdder U40 (w462, IN6[6], Out1[6], w477);
  FullAdder U41 (w477, w464, IN7[6], w478, w479);
  FullAdder U42 (w479, w466, IN8[6], w480, w481);
  FullAdder U43 (w481, w468, IN9[4], w482, w483);
  FullAdder U44 (w483, w470, IN10[3], w484, w485);
  FullAdder U45 (w485, w472, IN11[2], w486, w487);
  FullAdder U46 (w487, w474, IN12[1], w488, w489);
  FullAdder U47 (w489, w475, IN13[0], w490, w491);
  HalfAdder U48 (w478, IN7[7], Out1[7], w493);
  FullAdder U49 (w493, w480, IN8[7], w494, w495);
  FullAdder U50 (w495, w482, IN9[5], w496, w497);
  FullAdder U51 (w497, w484, IN10[4], w498, w499);
  FullAdder U52 (w499, w486, IN11[3], w500, w501);
  FullAdder U53 (w501, w488, IN12[2], w502, w503);
  FullAdder U54 (w503, w490, IN13[1], w504, w505);
  FullAdder U55 (w505, w491, IN14[0], w506, w507);
  HalfAdder U56 (w494, IN8[8], Out1[8], w509);
  FullAdder U57 (w509, w496, IN9[6], w510, w511);
  FullAdder U58 (w511, w498, IN10[5], w512, w513);
  FullAdder U59 (w513, w500, IN11[4], w514, w515);
  FullAdder U60 (w515, w502, IN12[3], w516, w517);
  FullAdder U61 (w517, w504, IN13[2], w518, w519);
  FullAdder U62 (w519, w506, IN14[1], w520, w521);
  FullAdder U63 (w521, w507, IN15[0], w522, w523);
  HalfAdder U64 (w510, IN9[7], Out1[9], w525);
  FullAdder U65 (w525, w512, IN10[6], w526, w527);
  FullAdder U66 (w527, w514, IN11[5], w528, w529);
  FullAdder U67 (w529, w516, IN12[4], w530, w531);
  FullAdder U68 (w531, w518, IN13[3], w532, w533);
  FullAdder U69 (w533, w520, IN14[2], w534, w535);
  FullAdder U70 (w535, w522, IN15[1], w536, w537);
  FullAdder U71 (w537, w523, IN16[0], w538, w539);
  HalfAdder U72 (w526, IN10[7], Out1[10], w541);
  FullAdder U73 (w541, w528, IN11[6], w542, w543);
  FullAdder U74 (w543, w530, IN12[5], w544, w545);
  FullAdder U75 (w545, w532, IN13[4], w546, w547);
  FullAdder U76 (w547, w534, IN14[3], w548, w549);
  FullAdder U77 (w549, w536, IN15[2], w550, w551);
  FullAdder U78 (w551, w538, IN16[1], w552, w553);
  FullAdder U79 (w553, w539, IN17[0], w554, w555);
  HalfAdder U80 (w542, IN11[7], Out1[11], w557);
  FullAdder U81 (w557, w544, IN12[6], w558, w559);
  FullAdder U82 (w559, w546, IN13[5], w560, w561);
  FullAdder U83 (w561, w548, IN14[4], w562, w563);
  FullAdder U84 (w563, w550, IN15[3], w564, w565);
  FullAdder U85 (w565, w552, IN16[2], w566, w567);
  FullAdder U86 (w567, w554, IN17[1], w568, w569);
  FullAdder U87 (w569, w555, IN18[0], w570, w571);
  HalfAdder U88 (w558, IN12[7], Out1[12], w573);
  FullAdder U89 (w573, w560, IN13[6], w574, w575);
  FullAdder U90 (w575, w562, IN14[5], w576, w577);
  FullAdder U91 (w577, w564, IN15[4], w578, w579);
  FullAdder U92 (w579, w566, IN16[3], w580, w581);
  FullAdder U93 (w581, w568, IN17[2], w582, w583);
  FullAdder U94 (w583, w570, IN18[1], w584, w585);
  FullAdder U95 (w585, w571, IN19[0], w586, w587);
  HalfAdder U96 (w574, IN13[7], Out1[13], w589);
  FullAdder U97 (w589, w576, IN14[6], w590, w591);
  FullAdder U98 (w591, w578, IN15[5], w592, w593);
  FullAdder U99 (w593, w580, IN16[4], w594, w595);
  FullAdder U100 (w595, w582, IN17[3], w596, w597);
  FullAdder U101 (w597, w584, IN18[2], w598, w599);
  FullAdder U102 (w599, w586, IN19[1], w600, w601);
  FullAdder U103 (w601, w587, IN20[0], w602, w603);
  HalfAdder U104 (w590, IN14[7], Out1[14], w605);
  FullAdder U105 (w605, w592, IN15[6], w606, w607);
  FullAdder U106 (w607, w594, IN16[5], w608, w609);
  FullAdder U107 (w609, w596, IN17[4], w610, w611);
  FullAdder U108 (w611, w598, IN18[3], w612, w613);
  FullAdder U109 (w613, w600, IN19[2], w614, w615);
  FullAdder U110 (w615, w602, IN20[1], w616, w617);
  FullAdder U111 (w617, w603, IN21[0], w618, w619);
  HalfAdder U112 (w606, IN15[7], Out1[15], w621);
  FullAdder U113 (w621, w608, IN16[6], w622, w623);
  FullAdder U114 (w623, w610, IN17[5], w624, w625);
  FullAdder U115 (w625, w612, IN18[4], w626, w627);
  FullAdder U116 (w627, w614, IN19[3], w628, w629);
  FullAdder U117 (w629, w616, IN20[2], w630, w631);
  FullAdder U118 (w631, w618, IN21[1], w632, w633);
  FullAdder U119 (w633, w619, IN22[0], w634, w635);
  HalfAdder U120 (w622, IN16[7], Out1[16], w637);
  FullAdder U121 (w637, w624, IN17[6], w638, w639);
  FullAdder U122 (w639, w626, IN18[5], w640, w641);
  FullAdder U123 (w641, w628, IN19[4], w642, w643);
  FullAdder U124 (w643, w630, IN20[3], w644, w645);
  FullAdder U125 (w645, w632, IN21[2], w646, w647);
  FullAdder U126 (w647, w634, IN22[1], w648, w649);
  FullAdder U127 (w649, w635, IN23[0], w650, w651);
  HalfAdder U128 (w638, IN17[7], Out1[17], w653);
  FullAdder U129 (w653, w640, IN18[6], w654, w655);
  FullAdder U130 (w655, w642, IN19[5], w656, w657);
  FullAdder U131 (w657, w644, IN20[4], w658, w659);
  FullAdder U132 (w659, w646, IN21[3], w660, w661);
  FullAdder U133 (w661, w648, IN22[2], w662, w663);
  FullAdder U134 (w663, w650, IN23[1], w664, w665);
  FullAdder U135 (w665, w651, IN24[0], w666, w667);
  HalfAdder U136 (w654, IN18[7], Out1[18], w669);
  FullAdder U137 (w669, w656, IN19[6], w670, w671);
  FullAdder U138 (w671, w658, IN20[5], w672, w673);
  FullAdder U139 (w673, w660, IN21[4], w674, w675);
  FullAdder U140 (w675, w662, IN22[3], w676, w677);
  FullAdder U141 (w677, w664, IN23[2], w678, w679);
  FullAdder U142 (w679, w666, IN24[1], w680, w681);
  FullAdder U143 (w681, w667, IN25[0], w682, w683);
  HalfAdder U144 (w670, IN19[7], Out1[19], w685);
  FullAdder U145 (w685, w672, IN20[6], w686, w687);
  FullAdder U146 (w687, w674, IN21[5], w688, w689);
  FullAdder U147 (w689, w676, IN22[4], w690, w691);
  FullAdder U148 (w691, w678, IN23[3], w692, w693);
  FullAdder U149 (w693, w680, IN24[2], w694, w695);
  FullAdder U150 (w695, w682, IN25[1], w696, w697);
  FullAdder U151 (w697, w683, IN26[0], w698, w699);
  HalfAdder U152 (w686, IN20[7], Out1[20], w701);
  FullAdder U153 (w701, w688, IN21[6], w702, w703);
  FullAdder U154 (w703, w690, IN22[5], w704, w705);
  FullAdder U155 (w705, w692, IN23[4], w706, w707);
  FullAdder U156 (w707, w694, IN24[3], w708, w709);
  FullAdder U157 (w709, w696, IN25[2], w710, w711);
  FullAdder U158 (w711, w698, IN26[1], w712, w713);
  FullAdder U159 (w713, w699, IN27[0], w714, w715);
  HalfAdder U160 (w702, IN21[7], Out1[21], w717);
  FullAdder U161 (w717, w704, IN22[6], w718, w719);
  FullAdder U162 (w719, w706, IN23[5], w720, w721);
  FullAdder U163 (w721, w708, IN24[4], w722, w723);
  FullAdder U164 (w723, w710, IN25[3], w724, w725);
  FullAdder U165 (w725, w712, IN26[2], w726, w727);
  FullAdder U166 (w727, w714, IN27[1], w728, w729);
  FullAdder U167 (w729, w715, IN28[0], w730, w731);
  HalfAdder U168 (w718, IN22[7], Out1[22], w733);
  FullAdder U169 (w733, w720, IN23[6], w734, w735);
  FullAdder U170 (w735, w722, IN24[5], w736, w737);
  FullAdder U171 (w737, w724, IN25[4], w738, w739);
  FullAdder U172 (w739, w726, IN26[3], w740, w741);
  FullAdder U173 (w741, w728, IN27[2], w742, w743);
  FullAdder U174 (w743, w730, IN28[1], w744, w745);
  FullAdder U175 (w745, w731, IN29[0], w746, w747);
  HalfAdder U176 (w734, IN23[7], Out1[23], w749);
  FullAdder U177 (w749, w736, IN24[6], w750, w751);
  FullAdder U178 (w751, w738, IN25[5], w752, w753);
  FullAdder U179 (w753, w740, IN26[4], w754, w755);
  FullAdder U180 (w755, w742, IN27[3], w756, w757);
  FullAdder U181 (w757, w744, IN28[2], w758, w759);
  FullAdder U182 (w759, w746, IN29[1], w760, w761);
  FullAdder U183 (w761, w747, IN30[0], w762, w763);
  HalfAdder U184 (w750, IN24[7], Out1[24], w765);
  FullAdder U185 (w765, w752, IN25[6], w766, w767);
  FullAdder U186 (w767, w754, IN26[5], w768, w769);
  FullAdder U187 (w769, w756, IN27[4], w770, w771);
  FullAdder U188 (w771, w758, IN28[3], w772, w773);
  FullAdder U189 (w773, w760, IN29[2], w774, w775);
  FullAdder U190 (w775, w762, IN30[1], w776, w777);
  FullAdder U191 (w777, w763, IN31[0], w778, w779);
  HalfAdder U192 (w766, IN25[7], Out1[25], w781);
  FullAdder U193 (w781, w768, IN26[6], w782, w783);
  FullAdder U194 (w783, w770, IN27[5], w784, w785);
  FullAdder U195 (w785, w772, IN28[4], w786, w787);
  FullAdder U196 (w787, w774, IN29[3], w788, w789);
  FullAdder U197 (w789, w776, IN30[2], w790, w791);
  FullAdder U198 (w791, w778, IN31[1], w792, w793);
  FullAdder U199 (w793, w779, IN32[0], w794, w795);
  HalfAdder U200 (w782, IN26[7], Out1[26], w797);
  FullAdder U201 (w797, w784, IN27[6], w798, w799);
  FullAdder U202 (w799, w786, IN28[5], w800, w801);
  FullAdder U203 (w801, w788, IN29[4], w802, w803);
  FullAdder U204 (w803, w790, IN30[3], w804, w805);
  FullAdder U205 (w805, w792, IN31[2], w806, w807);
  FullAdder U206 (w807, w794, IN32[1], w808, w809);
  FullAdder U207 (w809, w795, IN33[0], w810, w811);
  HalfAdder U208 (w798, IN27[7], Out1[27], w813);
  FullAdder U209 (w813, w800, IN28[6], w814, w815);
  FullAdder U210 (w815, w802, IN29[5], w816, w817);
  FullAdder U211 (w817, w804, IN30[4], w818, w819);
  FullAdder U212 (w819, w806, IN31[3], w820, w821);
  FullAdder U213 (w821, w808, IN32[2], w822, w823);
  FullAdder U214 (w823, w810, IN33[1], w824, w825);
  FullAdder U215 (w825, w811, IN34[0], w826, w827);
  HalfAdder U216 (w814, IN28[7], Out1[28], w829);
  FullAdder U217 (w829, w816, IN29[6], w830, w831);
  FullAdder U218 (w831, w818, IN30[5], w832, w833);
  FullAdder U219 (w833, w820, IN31[4], w834, w835);
  FullAdder U220 (w835, w822, IN32[3], w836, w837);
  FullAdder U221 (w837, w824, IN33[2], w838, w839);
  FullAdder U222 (w839, w826, IN34[1], w840, w841);
  FullAdder U223 (w841, w827, IN35[0], w842, w843);
  HalfAdder U224 (w830, IN29[7], Out1[29], w845);
  FullAdder U225 (w845, w832, IN30[6], w846, w847);
  FullAdder U226 (w847, w834, IN31[5], w848, w849);
  FullAdder U227 (w849, w836, IN32[4], w850, w851);
  FullAdder U228 (w851, w838, IN33[3], w852, w853);
  FullAdder U229 (w853, w840, IN34[2], w854, w855);
  FullAdder U230 (w855, w842, IN35[1], w856, w857);
  FullAdder U231 (w857, w843, IN36[0], w858, w859);
  HalfAdder U232 (w846, IN30[7], Out1[30], w861);
  FullAdder U233 (w861, w848, IN31[6], w862, w863);
  FullAdder U234 (w863, w850, IN32[5], w864, w865);
  FullAdder U235 (w865, w852, IN33[4], w866, w867);
  FullAdder U236 (w867, w854, IN34[3], w868, w869);
  FullAdder U237 (w869, w856, IN35[2], w870, w871);
  FullAdder U238 (w871, w858, IN36[1], w872, w873);
  FullAdder U239 (w873, w859, IN37[0], w874, w875);
  HalfAdder U240 (w862, IN31[7], Out1[31], w877);
  FullAdder U241 (w877, w864, IN32[6], w878, w879);
  FullAdder U242 (w879, w866, IN33[5], w880, w881);
  FullAdder U243 (w881, w868, IN34[4], w882, w883);
  FullAdder U244 (w883, w870, IN35[3], w884, w885);
  FullAdder U245 (w885, w872, IN36[2], w886, w887);
  FullAdder U246 (w887, w874, IN37[1], w888, w889);
  FullAdder U247 (w889, w875, IN38[0], w890, w891);
  HalfAdder U248 (w878, IN32[7], Out1[32], w893);
  FullAdder U249 (w893, w880, IN33[6], w894, w895);
  FullAdder U250 (w895, w882, IN34[5], w896, w897);
  FullAdder U251 (w897, w884, IN35[4], w898, w899);
  FullAdder U252 (w899, w886, IN36[3], w900, w901);
  FullAdder U253 (w901, w888, IN37[2], w902, w903);
  FullAdder U254 (w903, w890, IN38[1], w904, w905);
  FullAdder U255 (w905, w891, IN39[0], w906, w907);
  HalfAdder U256 (w894, IN33[7], Out1[33], w909);
  FullAdder U257 (w909, w896, IN34[6], w910, w911);
  FullAdder U258 (w911, w898, IN35[5], w912, w913);
  FullAdder U259 (w913, w900, IN36[4], w914, w915);
  FullAdder U260 (w915, w902, IN37[3], w916, w917);
  FullAdder U261 (w917, w904, IN38[2], w918, w919);
  FullAdder U262 (w919, w906, IN39[1], w920, w921);
  FullAdder U263 (w921, w907, IN40[0], w922, w923);
  HalfAdder U264 (w910, IN34[7], Out1[34], w925);
  FullAdder U265 (w925, w912, IN35[6], w926, w927);
  FullAdder U266 (w927, w914, IN36[5], w928, w929);
  FullAdder U267 (w929, w916, IN37[4], w930, w931);
  FullAdder U268 (w931, w918, IN38[3], w932, w933);
  FullAdder U269 (w933, w920, IN39[2], w934, w935);
  FullAdder U270 (w935, w922, IN40[1], w936, w937);
  FullAdder U271 (w937, w923, IN41[0], w938, w939);
  HalfAdder U272 (w926, IN35[7], Out1[35], w941);
  FullAdder U273 (w941, w928, IN36[6], w942, w943);
  FullAdder U274 (w943, w930, IN37[5], w944, w945);
  FullAdder U275 (w945, w932, IN38[4], w946, w947);
  FullAdder U276 (w947, w934, IN39[3], w948, w949);
  FullAdder U277 (w949, w936, IN40[2], w950, w951);
  FullAdder U278 (w951, w938, IN41[1], w952, w953);
  FullAdder U279 (w953, w939, IN42[0], w954, w955);
  HalfAdder U280 (w942, IN36[7], Out1[36], w957);
  FullAdder U281 (w957, w944, IN37[6], w958, w959);
  FullAdder U282 (w959, w946, IN38[5], w960, w961);
  FullAdder U283 (w961, w948, IN39[4], w962, w963);
  FullAdder U284 (w963, w950, IN40[3], w964, w965);
  FullAdder U285 (w965, w952, IN41[2], w966, w967);
  FullAdder U286 (w967, w954, IN42[1], w968, w969);
  FullAdder U287 (w969, w955, IN43[0], w970, w971);
  HalfAdder U288 (w958, IN37[7], Out1[37], w973);
  FullAdder U289 (w973, w960, IN38[6], w974, w975);
  FullAdder U290 (w975, w962, IN39[5], w976, w977);
  FullAdder U291 (w977, w964, IN40[4], w978, w979);
  FullAdder U292 (w979, w966, IN41[3], w980, w981);
  FullAdder U293 (w981, w968, IN42[2], w982, w983);
  FullAdder U294 (w983, w970, IN43[1], w984, w985);
  FullAdder U295 (w985, w971, IN44[0], w986, w987);
  HalfAdder U296 (w974, IN38[7], Out1[38], w989);
  FullAdder U297 (w989, w976, IN39[6], w990, w991);
  FullAdder U298 (w991, w978, IN40[5], w992, w993);
  FullAdder U299 (w993, w980, IN41[4], w994, w995);
  FullAdder U300 (w995, w982, IN42[3], w996, w997);
  FullAdder U301 (w997, w984, IN43[2], w998, w999);
  FullAdder U302 (w999, w986, IN44[1], w1000, w1001);
  FullAdder U303 (w1001, w987, IN45[0], w1002, w1003);
  HalfAdder U304 (w990, IN39[7], Out1[39], w1005);
  FullAdder U305 (w1005, w992, IN40[6], w1006, w1007);
  FullAdder U306 (w1007, w994, IN41[5], w1008, w1009);
  FullAdder U307 (w1009, w996, IN42[4], w1010, w1011);
  FullAdder U308 (w1011, w998, IN43[3], w1012, w1013);
  FullAdder U309 (w1013, w1000, IN44[2], w1014, w1015);
  FullAdder U310 (w1015, w1002, IN45[1], w1016, w1017);
  FullAdder U311 (w1017, w1003, IN46[0], w1018, w1019);
  HalfAdder U312 (w1006, IN40[7], Out1[40], w1021);
  FullAdder U313 (w1021, w1008, IN41[6], w1022, w1023);
  FullAdder U314 (w1023, w1010, IN42[5], w1024, w1025);
  FullAdder U315 (w1025, w1012, IN43[4], w1026, w1027);
  FullAdder U316 (w1027, w1014, IN44[3], w1028, w1029);
  FullAdder U317 (w1029, w1016, IN45[2], w1030, w1031);
  FullAdder U318 (w1031, w1018, IN46[1], w1032, w1033);
  FullAdder U319 (w1033, w1019, IN47[0], w1034, w1035);
  HalfAdder U320 (w1022, IN41[7], Out1[41], w1037);
  FullAdder U321 (w1037, w1024, IN42[6], w1038, w1039);
  FullAdder U322 (w1039, w1026, IN43[5], w1040, w1041);
  FullAdder U323 (w1041, w1028, IN44[4], w1042, w1043);
  FullAdder U324 (w1043, w1030, IN45[3], w1044, w1045);
  FullAdder U325 (w1045, w1032, IN46[2], w1046, w1047);
  FullAdder U326 (w1047, w1034, IN47[1], w1048, w1049);
  FullAdder U327 (w1049, w1035, IN48[0], w1050, w1051);
  HalfAdder U328 (w1038, IN42[7], Out1[42], w1053);
  FullAdder U329 (w1053, w1040, IN43[6], w1054, w1055);
  FullAdder U330 (w1055, w1042, IN44[5], w1056, w1057);
  FullAdder U331 (w1057, w1044, IN45[4], w1058, w1059);
  FullAdder U332 (w1059, w1046, IN46[3], w1060, w1061);
  FullAdder U333 (w1061, w1048, IN47[2], w1062, w1063);
  FullAdder U334 (w1063, w1050, IN48[1], w1064, w1065);
  FullAdder U335 (w1065, w1051, IN49[0], w1066, w1067);
  HalfAdder U336 (w1054, IN43[7], Out1[43], w1069);
  FullAdder U337 (w1069, w1056, IN44[6], Out1[44], w1071);
  FullAdder U338 (w1071, w1058, IN45[5], Out1[45], w1073);
  FullAdder U339 (w1073, w1060, IN46[4], Out1[46], w1075);
  FullAdder U340 (w1075, w1062, IN47[3], Out1[47], w1077);
  FullAdder U341 (w1077, w1064, IN48[2], Out1[48], w1079);
  FullAdder U342 (w1079, w1066, IN49[1], Out1[49], w1081);
  FullAdder U343 (w1081, w1067, IN50[0], Out1[50], Out1[51]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN9[8];
  assign Out2[1] = IN10[8];
  assign Out2[2] = IN11[8];
  assign Out2[3] = IN12[8];
  assign Out2[4] = IN13[8];
  assign Out2[5] = IN14[8];
  assign Out2[6] = IN15[8];
  assign Out2[7] = IN16[8];
  assign Out2[8] = IN17[8];
  assign Out2[9] = IN18[8];
  assign Out2[10] = IN19[8];
  assign Out2[11] = IN20[8];
  assign Out2[12] = IN21[8];
  assign Out2[13] = IN22[8];
  assign Out2[14] = IN23[8];
  assign Out2[15] = IN24[8];
  assign Out2[16] = IN25[8];
  assign Out2[17] = IN26[8];
  assign Out2[18] = IN27[8];
  assign Out2[19] = IN28[8];
  assign Out2[20] = IN29[8];
  assign Out2[21] = IN30[8];
  assign Out2[22] = IN31[8];
  assign Out2[23] = IN32[8];
  assign Out2[24] = IN33[8];
  assign Out2[25] = IN34[8];
  assign Out2[26] = IN35[8];
  assign Out2[27] = IN36[8];
  assign Out2[28] = IN37[8];
  assign Out2[29] = IN38[8];
  assign Out2[30] = IN39[8];
  assign Out2[31] = IN40[8];
  assign Out2[32] = IN41[8];
  assign Out2[33] = IN42[8];
  assign Out2[34] = IN43[8];
  assign Out2[35] = IN44[7];
  assign Out2[36] = IN45[6];
  assign Out2[37] = IN46[5];
  assign Out2[38] = IN47[4];
  assign Out2[39] = IN48[3];
  assign Out2[40] = IN49[2];
  assign Out2[41] = IN50[1];
  assign Out2[42] = IN51[0];

endmodule
module RC_43_43(IN1, IN2, Out);
  input [42:0] IN1;
  input [42:0] IN2;
  output [43:0] Out;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w87);
  FullAdder U1 (IN1[1], IN2[1], w87, Out[1], w89);
  FullAdder U2 (IN1[2], IN2[2], w89, Out[2], w91);
  FullAdder U3 (IN1[3], IN2[3], w91, Out[3], w93);
  FullAdder U4 (IN1[4], IN2[4], w93, Out[4], w95);
  FullAdder U5 (IN1[5], IN2[5], w95, Out[5], w97);
  FullAdder U6 (IN1[6], IN2[6], w97, Out[6], w99);
  FullAdder U7 (IN1[7], IN2[7], w99, Out[7], w101);
  FullAdder U8 (IN1[8], IN2[8], w101, Out[8], w103);
  FullAdder U9 (IN1[9], IN2[9], w103, Out[9], w105);
  FullAdder U10 (IN1[10], IN2[10], w105, Out[10], w107);
  FullAdder U11 (IN1[11], IN2[11], w107, Out[11], w109);
  FullAdder U12 (IN1[12], IN2[12], w109, Out[12], w111);
  FullAdder U13 (IN1[13], IN2[13], w111, Out[13], w113);
  FullAdder U14 (IN1[14], IN2[14], w113, Out[14], w115);
  FullAdder U15 (IN1[15], IN2[15], w115, Out[15], w117);
  FullAdder U16 (IN1[16], IN2[16], w117, Out[16], w119);
  FullAdder U17 (IN1[17], IN2[17], w119, Out[17], w121);
  FullAdder U18 (IN1[18], IN2[18], w121, Out[18], w123);
  FullAdder U19 (IN1[19], IN2[19], w123, Out[19], w125);
  FullAdder U20 (IN1[20], IN2[20], w125, Out[20], w127);
  FullAdder U21 (IN1[21], IN2[21], w127, Out[21], w129);
  FullAdder U22 (IN1[22], IN2[22], w129, Out[22], w131);
  FullAdder U23 (IN1[23], IN2[23], w131, Out[23], w133);
  FullAdder U24 (IN1[24], IN2[24], w133, Out[24], w135);
  FullAdder U25 (IN1[25], IN2[25], w135, Out[25], w137);
  FullAdder U26 (IN1[26], IN2[26], w137, Out[26], w139);
  FullAdder U27 (IN1[27], IN2[27], w139, Out[27], w141);
  FullAdder U28 (IN1[28], IN2[28], w141, Out[28], w143);
  FullAdder U29 (IN1[29], IN2[29], w143, Out[29], w145);
  FullAdder U30 (IN1[30], IN2[30], w145, Out[30], w147);
  FullAdder U31 (IN1[31], IN2[31], w147, Out[31], w149);
  FullAdder U32 (IN1[32], IN2[32], w149, Out[32], w151);
  FullAdder U33 (IN1[33], IN2[33], w151, Out[33], w153);
  FullAdder U34 (IN1[34], IN2[34], w153, Out[34], w155);
  FullAdder U35 (IN1[35], IN2[35], w155, Out[35], w157);
  FullAdder U36 (IN1[36], IN2[36], w157, Out[36], w159);
  FullAdder U37 (IN1[37], IN2[37], w159, Out[37], w161);
  FullAdder U38 (IN1[38], IN2[38], w161, Out[38], w163);
  FullAdder U39 (IN1[39], IN2[39], w163, Out[39], w165);
  FullAdder U40 (IN1[40], IN2[40], w165, Out[40], w167);
  FullAdder U41 (IN1[41], IN2[41], w167, Out[41], w169);
  FullAdder U42 (IN1[42], IN2[42], w169, Out[42], Out[43]);

endmodule
module NR_9_44(IN1, IN2, Out);
  input [8:0] IN1;
  input [43:0] IN2;
  output [52:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [8:0] P9;
  wire [8:0] P10;
  wire [8:0] P11;
  wire [8:0] P12;
  wire [8:0] P13;
  wire [8:0] P14;
  wire [8:0] P15;
  wire [8:0] P16;
  wire [8:0] P17;
  wire [8:0] P18;
  wire [8:0] P19;
  wire [8:0] P20;
  wire [8:0] P21;
  wire [8:0] P22;
  wire [8:0] P23;
  wire [8:0] P24;
  wire [8:0] P25;
  wire [8:0] P26;
  wire [8:0] P27;
  wire [8:0] P28;
  wire [8:0] P29;
  wire [8:0] P30;
  wire [8:0] P31;
  wire [8:0] P32;
  wire [8:0] P33;
  wire [8:0] P34;
  wire [8:0] P35;
  wire [8:0] P36;
  wire [8:0] P37;
  wire [8:0] P38;
  wire [8:0] P39;
  wire [8:0] P40;
  wire [8:0] P41;
  wire [8:0] P42;
  wire [8:0] P43;
  wire [7:0] P44;
  wire [6:0] P45;
  wire [5:0] P46;
  wire [4:0] P47;
  wire [3:0] P48;
  wire [2:0] P49;
  wire [1:0] P50;
  wire [0:0] P51;
  wire [51:0] R1;
  wire [42:0] R2;
  wire [52:0] aOut;
  U_SP_9_44 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, R1, R2);
  RC_43_43 S2 (R1[51:9], R2, aOut[52:9]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign Out = aOut[52:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
