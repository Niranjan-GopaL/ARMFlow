//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 21
  second input length: 43
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_21_43(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  input [20:0] IN1;
  input [42:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [20:0] P21;
  output [20:0] P22;
  output [20:0] P23;
  output [20:0] P24;
  output [20:0] P25;
  output [20:0] P26;
  output [20:0] P27;
  output [20:0] P28;
  output [20:0] P29;
  output [20:0] P30;
  output [20:0] P31;
  output [20:0] P32;
  output [20:0] P33;
  output [20:0] P34;
  output [20:0] P35;
  output [20:0] P36;
  output [20:0] P37;
  output [20:0] P38;
  output [20:0] P39;
  output [20:0] P40;
  output [20:0] P41;
  output [20:0] P42;
  output [19:0] P43;
  output [18:0] P44;
  output [17:0] P45;
  output [16:0] P46;
  output [15:0] P47;
  output [14:0] P48;
  output [13:0] P49;
  output [12:0] P50;
  output [11:0] P51;
  output [10:0] P52;
  output [9:0] P53;
  output [8:0] P54;
  output [7:0] P55;
  output [6:0] P56;
  output [5:0] P57;
  output [4:0] P58;
  output [3:0] P59;
  output [2:0] P60;
  output [1:0] P61;
  output [0:0] P62;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[0] = IN1[1]&IN2[42];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[1] = IN1[2]&IN2[41];
  assign P44[0] = IN1[2]&IN2[42];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[2] = IN1[3]&IN2[40];
  assign P44[1] = IN1[3]&IN2[41];
  assign P45[0] = IN1[3]&IN2[42];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[3] = IN1[4]&IN2[39];
  assign P44[2] = IN1[4]&IN2[40];
  assign P45[1] = IN1[4]&IN2[41];
  assign P46[0] = IN1[4]&IN2[42];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[4] = IN1[5]&IN2[38];
  assign P44[3] = IN1[5]&IN2[39];
  assign P45[2] = IN1[5]&IN2[40];
  assign P46[1] = IN1[5]&IN2[41];
  assign P47[0] = IN1[5]&IN2[42];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[5] = IN1[6]&IN2[37];
  assign P44[4] = IN1[6]&IN2[38];
  assign P45[3] = IN1[6]&IN2[39];
  assign P46[2] = IN1[6]&IN2[40];
  assign P47[1] = IN1[6]&IN2[41];
  assign P48[0] = IN1[6]&IN2[42];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[6] = IN1[7]&IN2[36];
  assign P44[5] = IN1[7]&IN2[37];
  assign P45[4] = IN1[7]&IN2[38];
  assign P46[3] = IN1[7]&IN2[39];
  assign P47[2] = IN1[7]&IN2[40];
  assign P48[1] = IN1[7]&IN2[41];
  assign P49[0] = IN1[7]&IN2[42];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[7] = IN1[8]&IN2[35];
  assign P44[6] = IN1[8]&IN2[36];
  assign P45[5] = IN1[8]&IN2[37];
  assign P46[4] = IN1[8]&IN2[38];
  assign P47[3] = IN1[8]&IN2[39];
  assign P48[2] = IN1[8]&IN2[40];
  assign P49[1] = IN1[8]&IN2[41];
  assign P50[0] = IN1[8]&IN2[42];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[8] = IN1[9]&IN2[34];
  assign P44[7] = IN1[9]&IN2[35];
  assign P45[6] = IN1[9]&IN2[36];
  assign P46[5] = IN1[9]&IN2[37];
  assign P47[4] = IN1[9]&IN2[38];
  assign P48[3] = IN1[9]&IN2[39];
  assign P49[2] = IN1[9]&IN2[40];
  assign P50[1] = IN1[9]&IN2[41];
  assign P51[0] = IN1[9]&IN2[42];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[9] = IN1[10]&IN2[33];
  assign P44[8] = IN1[10]&IN2[34];
  assign P45[7] = IN1[10]&IN2[35];
  assign P46[6] = IN1[10]&IN2[36];
  assign P47[5] = IN1[10]&IN2[37];
  assign P48[4] = IN1[10]&IN2[38];
  assign P49[3] = IN1[10]&IN2[39];
  assign P50[2] = IN1[10]&IN2[40];
  assign P51[1] = IN1[10]&IN2[41];
  assign P52[0] = IN1[10]&IN2[42];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[10] = IN1[11]&IN2[32];
  assign P44[9] = IN1[11]&IN2[33];
  assign P45[8] = IN1[11]&IN2[34];
  assign P46[7] = IN1[11]&IN2[35];
  assign P47[6] = IN1[11]&IN2[36];
  assign P48[5] = IN1[11]&IN2[37];
  assign P49[4] = IN1[11]&IN2[38];
  assign P50[3] = IN1[11]&IN2[39];
  assign P51[2] = IN1[11]&IN2[40];
  assign P52[1] = IN1[11]&IN2[41];
  assign P53[0] = IN1[11]&IN2[42];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[11] = IN1[12]&IN2[31];
  assign P44[10] = IN1[12]&IN2[32];
  assign P45[9] = IN1[12]&IN2[33];
  assign P46[8] = IN1[12]&IN2[34];
  assign P47[7] = IN1[12]&IN2[35];
  assign P48[6] = IN1[12]&IN2[36];
  assign P49[5] = IN1[12]&IN2[37];
  assign P50[4] = IN1[12]&IN2[38];
  assign P51[3] = IN1[12]&IN2[39];
  assign P52[2] = IN1[12]&IN2[40];
  assign P53[1] = IN1[12]&IN2[41];
  assign P54[0] = IN1[12]&IN2[42];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[12] = IN1[13]&IN2[30];
  assign P44[11] = IN1[13]&IN2[31];
  assign P45[10] = IN1[13]&IN2[32];
  assign P46[9] = IN1[13]&IN2[33];
  assign P47[8] = IN1[13]&IN2[34];
  assign P48[7] = IN1[13]&IN2[35];
  assign P49[6] = IN1[13]&IN2[36];
  assign P50[5] = IN1[13]&IN2[37];
  assign P51[4] = IN1[13]&IN2[38];
  assign P52[3] = IN1[13]&IN2[39];
  assign P53[2] = IN1[13]&IN2[40];
  assign P54[1] = IN1[13]&IN2[41];
  assign P55[0] = IN1[13]&IN2[42];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[14] = IN1[14]&IN2[24];
  assign P39[14] = IN1[14]&IN2[25];
  assign P40[14] = IN1[14]&IN2[26];
  assign P41[14] = IN1[14]&IN2[27];
  assign P42[14] = IN1[14]&IN2[28];
  assign P43[13] = IN1[14]&IN2[29];
  assign P44[12] = IN1[14]&IN2[30];
  assign P45[11] = IN1[14]&IN2[31];
  assign P46[10] = IN1[14]&IN2[32];
  assign P47[9] = IN1[14]&IN2[33];
  assign P48[8] = IN1[14]&IN2[34];
  assign P49[7] = IN1[14]&IN2[35];
  assign P50[6] = IN1[14]&IN2[36];
  assign P51[5] = IN1[14]&IN2[37];
  assign P52[4] = IN1[14]&IN2[38];
  assign P53[3] = IN1[14]&IN2[39];
  assign P54[2] = IN1[14]&IN2[40];
  assign P55[1] = IN1[14]&IN2[41];
  assign P56[0] = IN1[14]&IN2[42];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[15] = IN1[15]&IN2[23];
  assign P39[15] = IN1[15]&IN2[24];
  assign P40[15] = IN1[15]&IN2[25];
  assign P41[15] = IN1[15]&IN2[26];
  assign P42[15] = IN1[15]&IN2[27];
  assign P43[14] = IN1[15]&IN2[28];
  assign P44[13] = IN1[15]&IN2[29];
  assign P45[12] = IN1[15]&IN2[30];
  assign P46[11] = IN1[15]&IN2[31];
  assign P47[10] = IN1[15]&IN2[32];
  assign P48[9] = IN1[15]&IN2[33];
  assign P49[8] = IN1[15]&IN2[34];
  assign P50[7] = IN1[15]&IN2[35];
  assign P51[6] = IN1[15]&IN2[36];
  assign P52[5] = IN1[15]&IN2[37];
  assign P53[4] = IN1[15]&IN2[38];
  assign P54[3] = IN1[15]&IN2[39];
  assign P55[2] = IN1[15]&IN2[40];
  assign P56[1] = IN1[15]&IN2[41];
  assign P57[0] = IN1[15]&IN2[42];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[16] = IN1[16]&IN2[22];
  assign P39[16] = IN1[16]&IN2[23];
  assign P40[16] = IN1[16]&IN2[24];
  assign P41[16] = IN1[16]&IN2[25];
  assign P42[16] = IN1[16]&IN2[26];
  assign P43[15] = IN1[16]&IN2[27];
  assign P44[14] = IN1[16]&IN2[28];
  assign P45[13] = IN1[16]&IN2[29];
  assign P46[12] = IN1[16]&IN2[30];
  assign P47[11] = IN1[16]&IN2[31];
  assign P48[10] = IN1[16]&IN2[32];
  assign P49[9] = IN1[16]&IN2[33];
  assign P50[8] = IN1[16]&IN2[34];
  assign P51[7] = IN1[16]&IN2[35];
  assign P52[6] = IN1[16]&IN2[36];
  assign P53[5] = IN1[16]&IN2[37];
  assign P54[4] = IN1[16]&IN2[38];
  assign P55[3] = IN1[16]&IN2[39];
  assign P56[2] = IN1[16]&IN2[40];
  assign P57[1] = IN1[16]&IN2[41];
  assign P58[0] = IN1[16]&IN2[42];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[17] = IN1[17]&IN2[21];
  assign P39[17] = IN1[17]&IN2[22];
  assign P40[17] = IN1[17]&IN2[23];
  assign P41[17] = IN1[17]&IN2[24];
  assign P42[17] = IN1[17]&IN2[25];
  assign P43[16] = IN1[17]&IN2[26];
  assign P44[15] = IN1[17]&IN2[27];
  assign P45[14] = IN1[17]&IN2[28];
  assign P46[13] = IN1[17]&IN2[29];
  assign P47[12] = IN1[17]&IN2[30];
  assign P48[11] = IN1[17]&IN2[31];
  assign P49[10] = IN1[17]&IN2[32];
  assign P50[9] = IN1[17]&IN2[33];
  assign P51[8] = IN1[17]&IN2[34];
  assign P52[7] = IN1[17]&IN2[35];
  assign P53[6] = IN1[17]&IN2[36];
  assign P54[5] = IN1[17]&IN2[37];
  assign P55[4] = IN1[17]&IN2[38];
  assign P56[3] = IN1[17]&IN2[39];
  assign P57[2] = IN1[17]&IN2[40];
  assign P58[1] = IN1[17]&IN2[41];
  assign P59[0] = IN1[17]&IN2[42];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[18] = IN1[18]&IN2[20];
  assign P39[18] = IN1[18]&IN2[21];
  assign P40[18] = IN1[18]&IN2[22];
  assign P41[18] = IN1[18]&IN2[23];
  assign P42[18] = IN1[18]&IN2[24];
  assign P43[17] = IN1[18]&IN2[25];
  assign P44[16] = IN1[18]&IN2[26];
  assign P45[15] = IN1[18]&IN2[27];
  assign P46[14] = IN1[18]&IN2[28];
  assign P47[13] = IN1[18]&IN2[29];
  assign P48[12] = IN1[18]&IN2[30];
  assign P49[11] = IN1[18]&IN2[31];
  assign P50[10] = IN1[18]&IN2[32];
  assign P51[9] = IN1[18]&IN2[33];
  assign P52[8] = IN1[18]&IN2[34];
  assign P53[7] = IN1[18]&IN2[35];
  assign P54[6] = IN1[18]&IN2[36];
  assign P55[5] = IN1[18]&IN2[37];
  assign P56[4] = IN1[18]&IN2[38];
  assign P57[3] = IN1[18]&IN2[39];
  assign P58[2] = IN1[18]&IN2[40];
  assign P59[1] = IN1[18]&IN2[41];
  assign P60[0] = IN1[18]&IN2[42];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[19] = IN1[19]&IN2[19];
  assign P39[19] = IN1[19]&IN2[20];
  assign P40[19] = IN1[19]&IN2[21];
  assign P41[19] = IN1[19]&IN2[22];
  assign P42[19] = IN1[19]&IN2[23];
  assign P43[18] = IN1[19]&IN2[24];
  assign P44[17] = IN1[19]&IN2[25];
  assign P45[16] = IN1[19]&IN2[26];
  assign P46[15] = IN1[19]&IN2[27];
  assign P47[14] = IN1[19]&IN2[28];
  assign P48[13] = IN1[19]&IN2[29];
  assign P49[12] = IN1[19]&IN2[30];
  assign P50[11] = IN1[19]&IN2[31];
  assign P51[10] = IN1[19]&IN2[32];
  assign P52[9] = IN1[19]&IN2[33];
  assign P53[8] = IN1[19]&IN2[34];
  assign P54[7] = IN1[19]&IN2[35];
  assign P55[6] = IN1[19]&IN2[36];
  assign P56[5] = IN1[19]&IN2[37];
  assign P57[4] = IN1[19]&IN2[38];
  assign P58[3] = IN1[19]&IN2[39];
  assign P59[2] = IN1[19]&IN2[40];
  assign P60[1] = IN1[19]&IN2[41];
  assign P61[0] = IN1[19]&IN2[42];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[20] = IN1[20]&IN2[18];
  assign P39[20] = IN1[20]&IN2[19];
  assign P40[20] = IN1[20]&IN2[20];
  assign P41[20] = IN1[20]&IN2[21];
  assign P42[20] = IN1[20]&IN2[22];
  assign P43[19] = IN1[20]&IN2[23];
  assign P44[18] = IN1[20]&IN2[24];
  assign P45[17] = IN1[20]&IN2[25];
  assign P46[16] = IN1[20]&IN2[26];
  assign P47[15] = IN1[20]&IN2[27];
  assign P48[14] = IN1[20]&IN2[28];
  assign P49[13] = IN1[20]&IN2[29];
  assign P50[12] = IN1[20]&IN2[30];
  assign P51[11] = IN1[20]&IN2[31];
  assign P52[10] = IN1[20]&IN2[32];
  assign P53[9] = IN1[20]&IN2[33];
  assign P54[8] = IN1[20]&IN2[34];
  assign P55[7] = IN1[20]&IN2[35];
  assign P56[6] = IN1[20]&IN2[36];
  assign P57[5] = IN1[20]&IN2[37];
  assign P58[4] = IN1[20]&IN2[38];
  assign P59[3] = IN1[20]&IN2[39];
  assign P60[2] = IN1[20]&IN2[40];
  assign P61[1] = IN1[20]&IN2[41];
  assign P62[0] = IN1[20]&IN2[42];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [20:0] IN21;
  input [20:0] IN22;
  input [20:0] IN23;
  input [20:0] IN24;
  input [20:0] IN25;
  input [20:0] IN26;
  input [20:0] IN27;
  input [20:0] IN28;
  input [20:0] IN29;
  input [20:0] IN30;
  input [20:0] IN31;
  input [20:0] IN32;
  input [20:0] IN33;
  input [20:0] IN34;
  input [20:0] IN35;
  input [20:0] IN36;
  input [20:0] IN37;
  input [20:0] IN38;
  input [20:0] IN39;
  input [20:0] IN40;
  input [20:0] IN41;
  input [20:0] IN42;
  input [19:0] IN43;
  input [18:0] IN44;
  input [17:0] IN45;
  input [16:0] IN46;
  input [15:0] IN47;
  input [14:0] IN48;
  input [13:0] IN49;
  input [12:0] IN50;
  input [11:0] IN51;
  input [10:0] IN52;
  input [9:0] IN53;
  input [8:0] IN54;
  input [7:0] IN55;
  input [6:0] IN56;
  input [5:0] IN57;
  input [4:0] IN58;
  input [3:0] IN59;
  input [2:0] IN60;
  input [1:0] IN61;
  input [0:0] IN62;
  output [62:0] Out1;
  output [41:0] Out2;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1984;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2050;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2088;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2140;
  wire w2141;
  wire w2142;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2544;
  wire w2546;
  wire w2548;
  wire w2550;
  wire w2552;
  wire w2554;
  wire w2556;
  wire w2558;
  wire w2560;
  wire w2562;
  wire w2564;
  wire w2566;
  wire w2568;
  wire w2570;
  wire w2572;
  wire w2574;
  wire w2576;
  wire w2578;
  wire w2580;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w904);
  FullAdder U1 (w904, IN2[0], IN2[1], w905, w906);
  FullAdder U2 (w906, IN3[0], IN3[1], w907, w908);
  FullAdder U3 (w908, IN4[0], IN4[1], w909, w910);
  FullAdder U4 (w910, IN5[0], IN5[1], w911, w912);
  FullAdder U5 (w912, IN6[0], IN6[1], w913, w914);
  FullAdder U6 (w914, IN7[0], IN7[1], w915, w916);
  FullAdder U7 (w916, IN8[0], IN8[1], w917, w918);
  FullAdder U8 (w918, IN9[0], IN9[1], w919, w920);
  FullAdder U9 (w920, IN10[0], IN10[1], w921, w922);
  FullAdder U10 (w922, IN11[0], IN11[1], w923, w924);
  FullAdder U11 (w924, IN12[0], IN12[1], w925, w926);
  FullAdder U12 (w926, IN13[0], IN13[1], w927, w928);
  FullAdder U13 (w928, IN14[0], IN14[1], w929, w930);
  FullAdder U14 (w930, IN15[0], IN15[1], w931, w932);
  FullAdder U15 (w932, IN16[0], IN16[1], w933, w934);
  FullAdder U16 (w934, IN17[0], IN17[1], w935, w936);
  FullAdder U17 (w936, IN18[0], IN18[1], w937, w938);
  FullAdder U18 (w938, IN19[0], IN19[1], w939, w940);
  FullAdder U19 (w940, IN20[0], IN20[1], w941, w942);
  HalfAdder U20 (w905, IN2[2], Out1[2], w944);
  FullAdder U21 (w944, w907, IN3[2], w945, w946);
  FullAdder U22 (w946, w909, IN4[2], w947, w948);
  FullAdder U23 (w948, w911, IN5[2], w949, w950);
  FullAdder U24 (w950, w913, IN6[2], w951, w952);
  FullAdder U25 (w952, w915, IN7[2], w953, w954);
  FullAdder U26 (w954, w917, IN8[2], w955, w956);
  FullAdder U27 (w956, w919, IN9[2], w957, w958);
  FullAdder U28 (w958, w921, IN10[2], w959, w960);
  FullAdder U29 (w960, w923, IN11[2], w961, w962);
  FullAdder U30 (w962, w925, IN12[2], w963, w964);
  FullAdder U31 (w964, w927, IN13[2], w965, w966);
  FullAdder U32 (w966, w929, IN14[2], w967, w968);
  FullAdder U33 (w968, w931, IN15[2], w969, w970);
  FullAdder U34 (w970, w933, IN16[2], w971, w972);
  FullAdder U35 (w972, w935, IN17[2], w973, w974);
  FullAdder U36 (w974, w937, IN18[2], w975, w976);
  FullAdder U37 (w976, w939, IN19[2], w977, w978);
  FullAdder U38 (w978, w941, IN20[2], w979, w980);
  FullAdder U39 (w980, w942, IN21[0], w981, w982);
  HalfAdder U40 (w945, IN3[3], Out1[3], w984);
  FullAdder U41 (w984, w947, IN4[3], w985, w986);
  FullAdder U42 (w986, w949, IN5[3], w987, w988);
  FullAdder U43 (w988, w951, IN6[3], w989, w990);
  FullAdder U44 (w990, w953, IN7[3], w991, w992);
  FullAdder U45 (w992, w955, IN8[3], w993, w994);
  FullAdder U46 (w994, w957, IN9[3], w995, w996);
  FullAdder U47 (w996, w959, IN10[3], w997, w998);
  FullAdder U48 (w998, w961, IN11[3], w999, w1000);
  FullAdder U49 (w1000, w963, IN12[3], w1001, w1002);
  FullAdder U50 (w1002, w965, IN13[3], w1003, w1004);
  FullAdder U51 (w1004, w967, IN14[3], w1005, w1006);
  FullAdder U52 (w1006, w969, IN15[3], w1007, w1008);
  FullAdder U53 (w1008, w971, IN16[3], w1009, w1010);
  FullAdder U54 (w1010, w973, IN17[3], w1011, w1012);
  FullAdder U55 (w1012, w975, IN18[3], w1013, w1014);
  FullAdder U56 (w1014, w977, IN19[3], w1015, w1016);
  FullAdder U57 (w1016, w979, IN20[3], w1017, w1018);
  FullAdder U58 (w1018, w981, IN21[1], w1019, w1020);
  FullAdder U59 (w1020, w982, IN22[0], w1021, w1022);
  HalfAdder U60 (w985, IN4[4], Out1[4], w1024);
  FullAdder U61 (w1024, w987, IN5[4], w1025, w1026);
  FullAdder U62 (w1026, w989, IN6[4], w1027, w1028);
  FullAdder U63 (w1028, w991, IN7[4], w1029, w1030);
  FullAdder U64 (w1030, w993, IN8[4], w1031, w1032);
  FullAdder U65 (w1032, w995, IN9[4], w1033, w1034);
  FullAdder U66 (w1034, w997, IN10[4], w1035, w1036);
  FullAdder U67 (w1036, w999, IN11[4], w1037, w1038);
  FullAdder U68 (w1038, w1001, IN12[4], w1039, w1040);
  FullAdder U69 (w1040, w1003, IN13[4], w1041, w1042);
  FullAdder U70 (w1042, w1005, IN14[4], w1043, w1044);
  FullAdder U71 (w1044, w1007, IN15[4], w1045, w1046);
  FullAdder U72 (w1046, w1009, IN16[4], w1047, w1048);
  FullAdder U73 (w1048, w1011, IN17[4], w1049, w1050);
  FullAdder U74 (w1050, w1013, IN18[4], w1051, w1052);
  FullAdder U75 (w1052, w1015, IN19[4], w1053, w1054);
  FullAdder U76 (w1054, w1017, IN20[4], w1055, w1056);
  FullAdder U77 (w1056, w1019, IN21[2], w1057, w1058);
  FullAdder U78 (w1058, w1021, IN22[1], w1059, w1060);
  FullAdder U79 (w1060, w1022, IN23[0], w1061, w1062);
  HalfAdder U80 (w1025, IN5[5], Out1[5], w1064);
  FullAdder U81 (w1064, w1027, IN6[5], w1065, w1066);
  FullAdder U82 (w1066, w1029, IN7[5], w1067, w1068);
  FullAdder U83 (w1068, w1031, IN8[5], w1069, w1070);
  FullAdder U84 (w1070, w1033, IN9[5], w1071, w1072);
  FullAdder U85 (w1072, w1035, IN10[5], w1073, w1074);
  FullAdder U86 (w1074, w1037, IN11[5], w1075, w1076);
  FullAdder U87 (w1076, w1039, IN12[5], w1077, w1078);
  FullAdder U88 (w1078, w1041, IN13[5], w1079, w1080);
  FullAdder U89 (w1080, w1043, IN14[5], w1081, w1082);
  FullAdder U90 (w1082, w1045, IN15[5], w1083, w1084);
  FullAdder U91 (w1084, w1047, IN16[5], w1085, w1086);
  FullAdder U92 (w1086, w1049, IN17[5], w1087, w1088);
  FullAdder U93 (w1088, w1051, IN18[5], w1089, w1090);
  FullAdder U94 (w1090, w1053, IN19[5], w1091, w1092);
  FullAdder U95 (w1092, w1055, IN20[5], w1093, w1094);
  FullAdder U96 (w1094, w1057, IN21[3], w1095, w1096);
  FullAdder U97 (w1096, w1059, IN22[2], w1097, w1098);
  FullAdder U98 (w1098, w1061, IN23[1], w1099, w1100);
  FullAdder U99 (w1100, w1062, IN24[0], w1101, w1102);
  HalfAdder U100 (w1065, IN6[6], Out1[6], w1104);
  FullAdder U101 (w1104, w1067, IN7[6], w1105, w1106);
  FullAdder U102 (w1106, w1069, IN8[6], w1107, w1108);
  FullAdder U103 (w1108, w1071, IN9[6], w1109, w1110);
  FullAdder U104 (w1110, w1073, IN10[6], w1111, w1112);
  FullAdder U105 (w1112, w1075, IN11[6], w1113, w1114);
  FullAdder U106 (w1114, w1077, IN12[6], w1115, w1116);
  FullAdder U107 (w1116, w1079, IN13[6], w1117, w1118);
  FullAdder U108 (w1118, w1081, IN14[6], w1119, w1120);
  FullAdder U109 (w1120, w1083, IN15[6], w1121, w1122);
  FullAdder U110 (w1122, w1085, IN16[6], w1123, w1124);
  FullAdder U111 (w1124, w1087, IN17[6], w1125, w1126);
  FullAdder U112 (w1126, w1089, IN18[6], w1127, w1128);
  FullAdder U113 (w1128, w1091, IN19[6], w1129, w1130);
  FullAdder U114 (w1130, w1093, IN20[6], w1131, w1132);
  FullAdder U115 (w1132, w1095, IN21[4], w1133, w1134);
  FullAdder U116 (w1134, w1097, IN22[3], w1135, w1136);
  FullAdder U117 (w1136, w1099, IN23[2], w1137, w1138);
  FullAdder U118 (w1138, w1101, IN24[1], w1139, w1140);
  FullAdder U119 (w1140, w1102, IN25[0], w1141, w1142);
  HalfAdder U120 (w1105, IN7[7], Out1[7], w1144);
  FullAdder U121 (w1144, w1107, IN8[7], w1145, w1146);
  FullAdder U122 (w1146, w1109, IN9[7], w1147, w1148);
  FullAdder U123 (w1148, w1111, IN10[7], w1149, w1150);
  FullAdder U124 (w1150, w1113, IN11[7], w1151, w1152);
  FullAdder U125 (w1152, w1115, IN12[7], w1153, w1154);
  FullAdder U126 (w1154, w1117, IN13[7], w1155, w1156);
  FullAdder U127 (w1156, w1119, IN14[7], w1157, w1158);
  FullAdder U128 (w1158, w1121, IN15[7], w1159, w1160);
  FullAdder U129 (w1160, w1123, IN16[7], w1161, w1162);
  FullAdder U130 (w1162, w1125, IN17[7], w1163, w1164);
  FullAdder U131 (w1164, w1127, IN18[7], w1165, w1166);
  FullAdder U132 (w1166, w1129, IN19[7], w1167, w1168);
  FullAdder U133 (w1168, w1131, IN20[7], w1169, w1170);
  FullAdder U134 (w1170, w1133, IN21[5], w1171, w1172);
  FullAdder U135 (w1172, w1135, IN22[4], w1173, w1174);
  FullAdder U136 (w1174, w1137, IN23[3], w1175, w1176);
  FullAdder U137 (w1176, w1139, IN24[2], w1177, w1178);
  FullAdder U138 (w1178, w1141, IN25[1], w1179, w1180);
  FullAdder U139 (w1180, w1142, IN26[0], w1181, w1182);
  HalfAdder U140 (w1145, IN8[8], Out1[8], w1184);
  FullAdder U141 (w1184, w1147, IN9[8], w1185, w1186);
  FullAdder U142 (w1186, w1149, IN10[8], w1187, w1188);
  FullAdder U143 (w1188, w1151, IN11[8], w1189, w1190);
  FullAdder U144 (w1190, w1153, IN12[8], w1191, w1192);
  FullAdder U145 (w1192, w1155, IN13[8], w1193, w1194);
  FullAdder U146 (w1194, w1157, IN14[8], w1195, w1196);
  FullAdder U147 (w1196, w1159, IN15[8], w1197, w1198);
  FullAdder U148 (w1198, w1161, IN16[8], w1199, w1200);
  FullAdder U149 (w1200, w1163, IN17[8], w1201, w1202);
  FullAdder U150 (w1202, w1165, IN18[8], w1203, w1204);
  FullAdder U151 (w1204, w1167, IN19[8], w1205, w1206);
  FullAdder U152 (w1206, w1169, IN20[8], w1207, w1208);
  FullAdder U153 (w1208, w1171, IN21[6], w1209, w1210);
  FullAdder U154 (w1210, w1173, IN22[5], w1211, w1212);
  FullAdder U155 (w1212, w1175, IN23[4], w1213, w1214);
  FullAdder U156 (w1214, w1177, IN24[3], w1215, w1216);
  FullAdder U157 (w1216, w1179, IN25[2], w1217, w1218);
  FullAdder U158 (w1218, w1181, IN26[1], w1219, w1220);
  FullAdder U159 (w1220, w1182, IN27[0], w1221, w1222);
  HalfAdder U160 (w1185, IN9[9], Out1[9], w1224);
  FullAdder U161 (w1224, w1187, IN10[9], w1225, w1226);
  FullAdder U162 (w1226, w1189, IN11[9], w1227, w1228);
  FullAdder U163 (w1228, w1191, IN12[9], w1229, w1230);
  FullAdder U164 (w1230, w1193, IN13[9], w1231, w1232);
  FullAdder U165 (w1232, w1195, IN14[9], w1233, w1234);
  FullAdder U166 (w1234, w1197, IN15[9], w1235, w1236);
  FullAdder U167 (w1236, w1199, IN16[9], w1237, w1238);
  FullAdder U168 (w1238, w1201, IN17[9], w1239, w1240);
  FullAdder U169 (w1240, w1203, IN18[9], w1241, w1242);
  FullAdder U170 (w1242, w1205, IN19[9], w1243, w1244);
  FullAdder U171 (w1244, w1207, IN20[9], w1245, w1246);
  FullAdder U172 (w1246, w1209, IN21[7], w1247, w1248);
  FullAdder U173 (w1248, w1211, IN22[6], w1249, w1250);
  FullAdder U174 (w1250, w1213, IN23[5], w1251, w1252);
  FullAdder U175 (w1252, w1215, IN24[4], w1253, w1254);
  FullAdder U176 (w1254, w1217, IN25[3], w1255, w1256);
  FullAdder U177 (w1256, w1219, IN26[2], w1257, w1258);
  FullAdder U178 (w1258, w1221, IN27[1], w1259, w1260);
  FullAdder U179 (w1260, w1222, IN28[0], w1261, w1262);
  HalfAdder U180 (w1225, IN10[10], Out1[10], w1264);
  FullAdder U181 (w1264, w1227, IN11[10], w1265, w1266);
  FullAdder U182 (w1266, w1229, IN12[10], w1267, w1268);
  FullAdder U183 (w1268, w1231, IN13[10], w1269, w1270);
  FullAdder U184 (w1270, w1233, IN14[10], w1271, w1272);
  FullAdder U185 (w1272, w1235, IN15[10], w1273, w1274);
  FullAdder U186 (w1274, w1237, IN16[10], w1275, w1276);
  FullAdder U187 (w1276, w1239, IN17[10], w1277, w1278);
  FullAdder U188 (w1278, w1241, IN18[10], w1279, w1280);
  FullAdder U189 (w1280, w1243, IN19[10], w1281, w1282);
  FullAdder U190 (w1282, w1245, IN20[10], w1283, w1284);
  FullAdder U191 (w1284, w1247, IN21[8], w1285, w1286);
  FullAdder U192 (w1286, w1249, IN22[7], w1287, w1288);
  FullAdder U193 (w1288, w1251, IN23[6], w1289, w1290);
  FullAdder U194 (w1290, w1253, IN24[5], w1291, w1292);
  FullAdder U195 (w1292, w1255, IN25[4], w1293, w1294);
  FullAdder U196 (w1294, w1257, IN26[3], w1295, w1296);
  FullAdder U197 (w1296, w1259, IN27[2], w1297, w1298);
  FullAdder U198 (w1298, w1261, IN28[1], w1299, w1300);
  FullAdder U199 (w1300, w1262, IN29[0], w1301, w1302);
  HalfAdder U200 (w1265, IN11[11], Out1[11], w1304);
  FullAdder U201 (w1304, w1267, IN12[11], w1305, w1306);
  FullAdder U202 (w1306, w1269, IN13[11], w1307, w1308);
  FullAdder U203 (w1308, w1271, IN14[11], w1309, w1310);
  FullAdder U204 (w1310, w1273, IN15[11], w1311, w1312);
  FullAdder U205 (w1312, w1275, IN16[11], w1313, w1314);
  FullAdder U206 (w1314, w1277, IN17[11], w1315, w1316);
  FullAdder U207 (w1316, w1279, IN18[11], w1317, w1318);
  FullAdder U208 (w1318, w1281, IN19[11], w1319, w1320);
  FullAdder U209 (w1320, w1283, IN20[11], w1321, w1322);
  FullAdder U210 (w1322, w1285, IN21[9], w1323, w1324);
  FullAdder U211 (w1324, w1287, IN22[8], w1325, w1326);
  FullAdder U212 (w1326, w1289, IN23[7], w1327, w1328);
  FullAdder U213 (w1328, w1291, IN24[6], w1329, w1330);
  FullAdder U214 (w1330, w1293, IN25[5], w1331, w1332);
  FullAdder U215 (w1332, w1295, IN26[4], w1333, w1334);
  FullAdder U216 (w1334, w1297, IN27[3], w1335, w1336);
  FullAdder U217 (w1336, w1299, IN28[2], w1337, w1338);
  FullAdder U218 (w1338, w1301, IN29[1], w1339, w1340);
  FullAdder U219 (w1340, w1302, IN30[0], w1341, w1342);
  HalfAdder U220 (w1305, IN12[12], Out1[12], w1344);
  FullAdder U221 (w1344, w1307, IN13[12], w1345, w1346);
  FullAdder U222 (w1346, w1309, IN14[12], w1347, w1348);
  FullAdder U223 (w1348, w1311, IN15[12], w1349, w1350);
  FullAdder U224 (w1350, w1313, IN16[12], w1351, w1352);
  FullAdder U225 (w1352, w1315, IN17[12], w1353, w1354);
  FullAdder U226 (w1354, w1317, IN18[12], w1355, w1356);
  FullAdder U227 (w1356, w1319, IN19[12], w1357, w1358);
  FullAdder U228 (w1358, w1321, IN20[12], w1359, w1360);
  FullAdder U229 (w1360, w1323, IN21[10], w1361, w1362);
  FullAdder U230 (w1362, w1325, IN22[9], w1363, w1364);
  FullAdder U231 (w1364, w1327, IN23[8], w1365, w1366);
  FullAdder U232 (w1366, w1329, IN24[7], w1367, w1368);
  FullAdder U233 (w1368, w1331, IN25[6], w1369, w1370);
  FullAdder U234 (w1370, w1333, IN26[5], w1371, w1372);
  FullAdder U235 (w1372, w1335, IN27[4], w1373, w1374);
  FullAdder U236 (w1374, w1337, IN28[3], w1375, w1376);
  FullAdder U237 (w1376, w1339, IN29[2], w1377, w1378);
  FullAdder U238 (w1378, w1341, IN30[1], w1379, w1380);
  FullAdder U239 (w1380, w1342, IN31[0], w1381, w1382);
  HalfAdder U240 (w1345, IN13[13], Out1[13], w1384);
  FullAdder U241 (w1384, w1347, IN14[13], w1385, w1386);
  FullAdder U242 (w1386, w1349, IN15[13], w1387, w1388);
  FullAdder U243 (w1388, w1351, IN16[13], w1389, w1390);
  FullAdder U244 (w1390, w1353, IN17[13], w1391, w1392);
  FullAdder U245 (w1392, w1355, IN18[13], w1393, w1394);
  FullAdder U246 (w1394, w1357, IN19[13], w1395, w1396);
  FullAdder U247 (w1396, w1359, IN20[13], w1397, w1398);
  FullAdder U248 (w1398, w1361, IN21[11], w1399, w1400);
  FullAdder U249 (w1400, w1363, IN22[10], w1401, w1402);
  FullAdder U250 (w1402, w1365, IN23[9], w1403, w1404);
  FullAdder U251 (w1404, w1367, IN24[8], w1405, w1406);
  FullAdder U252 (w1406, w1369, IN25[7], w1407, w1408);
  FullAdder U253 (w1408, w1371, IN26[6], w1409, w1410);
  FullAdder U254 (w1410, w1373, IN27[5], w1411, w1412);
  FullAdder U255 (w1412, w1375, IN28[4], w1413, w1414);
  FullAdder U256 (w1414, w1377, IN29[3], w1415, w1416);
  FullAdder U257 (w1416, w1379, IN30[2], w1417, w1418);
  FullAdder U258 (w1418, w1381, IN31[1], w1419, w1420);
  FullAdder U259 (w1420, w1382, IN32[0], w1421, w1422);
  HalfAdder U260 (w1385, IN14[14], Out1[14], w1424);
  FullAdder U261 (w1424, w1387, IN15[14], w1425, w1426);
  FullAdder U262 (w1426, w1389, IN16[14], w1427, w1428);
  FullAdder U263 (w1428, w1391, IN17[14], w1429, w1430);
  FullAdder U264 (w1430, w1393, IN18[14], w1431, w1432);
  FullAdder U265 (w1432, w1395, IN19[14], w1433, w1434);
  FullAdder U266 (w1434, w1397, IN20[14], w1435, w1436);
  FullAdder U267 (w1436, w1399, IN21[12], w1437, w1438);
  FullAdder U268 (w1438, w1401, IN22[11], w1439, w1440);
  FullAdder U269 (w1440, w1403, IN23[10], w1441, w1442);
  FullAdder U270 (w1442, w1405, IN24[9], w1443, w1444);
  FullAdder U271 (w1444, w1407, IN25[8], w1445, w1446);
  FullAdder U272 (w1446, w1409, IN26[7], w1447, w1448);
  FullAdder U273 (w1448, w1411, IN27[6], w1449, w1450);
  FullAdder U274 (w1450, w1413, IN28[5], w1451, w1452);
  FullAdder U275 (w1452, w1415, IN29[4], w1453, w1454);
  FullAdder U276 (w1454, w1417, IN30[3], w1455, w1456);
  FullAdder U277 (w1456, w1419, IN31[2], w1457, w1458);
  FullAdder U278 (w1458, w1421, IN32[1], w1459, w1460);
  FullAdder U279 (w1460, w1422, IN33[0], w1461, w1462);
  HalfAdder U280 (w1425, IN15[15], Out1[15], w1464);
  FullAdder U281 (w1464, w1427, IN16[15], w1465, w1466);
  FullAdder U282 (w1466, w1429, IN17[15], w1467, w1468);
  FullAdder U283 (w1468, w1431, IN18[15], w1469, w1470);
  FullAdder U284 (w1470, w1433, IN19[15], w1471, w1472);
  FullAdder U285 (w1472, w1435, IN20[15], w1473, w1474);
  FullAdder U286 (w1474, w1437, IN21[13], w1475, w1476);
  FullAdder U287 (w1476, w1439, IN22[12], w1477, w1478);
  FullAdder U288 (w1478, w1441, IN23[11], w1479, w1480);
  FullAdder U289 (w1480, w1443, IN24[10], w1481, w1482);
  FullAdder U290 (w1482, w1445, IN25[9], w1483, w1484);
  FullAdder U291 (w1484, w1447, IN26[8], w1485, w1486);
  FullAdder U292 (w1486, w1449, IN27[7], w1487, w1488);
  FullAdder U293 (w1488, w1451, IN28[6], w1489, w1490);
  FullAdder U294 (w1490, w1453, IN29[5], w1491, w1492);
  FullAdder U295 (w1492, w1455, IN30[4], w1493, w1494);
  FullAdder U296 (w1494, w1457, IN31[3], w1495, w1496);
  FullAdder U297 (w1496, w1459, IN32[2], w1497, w1498);
  FullAdder U298 (w1498, w1461, IN33[1], w1499, w1500);
  FullAdder U299 (w1500, w1462, IN34[0], w1501, w1502);
  HalfAdder U300 (w1465, IN16[16], Out1[16], w1504);
  FullAdder U301 (w1504, w1467, IN17[16], w1505, w1506);
  FullAdder U302 (w1506, w1469, IN18[16], w1507, w1508);
  FullAdder U303 (w1508, w1471, IN19[16], w1509, w1510);
  FullAdder U304 (w1510, w1473, IN20[16], w1511, w1512);
  FullAdder U305 (w1512, w1475, IN21[14], w1513, w1514);
  FullAdder U306 (w1514, w1477, IN22[13], w1515, w1516);
  FullAdder U307 (w1516, w1479, IN23[12], w1517, w1518);
  FullAdder U308 (w1518, w1481, IN24[11], w1519, w1520);
  FullAdder U309 (w1520, w1483, IN25[10], w1521, w1522);
  FullAdder U310 (w1522, w1485, IN26[9], w1523, w1524);
  FullAdder U311 (w1524, w1487, IN27[8], w1525, w1526);
  FullAdder U312 (w1526, w1489, IN28[7], w1527, w1528);
  FullAdder U313 (w1528, w1491, IN29[6], w1529, w1530);
  FullAdder U314 (w1530, w1493, IN30[5], w1531, w1532);
  FullAdder U315 (w1532, w1495, IN31[4], w1533, w1534);
  FullAdder U316 (w1534, w1497, IN32[3], w1535, w1536);
  FullAdder U317 (w1536, w1499, IN33[2], w1537, w1538);
  FullAdder U318 (w1538, w1501, IN34[1], w1539, w1540);
  FullAdder U319 (w1540, w1502, IN35[0], w1541, w1542);
  HalfAdder U320 (w1505, IN17[17], Out1[17], w1544);
  FullAdder U321 (w1544, w1507, IN18[17], w1545, w1546);
  FullAdder U322 (w1546, w1509, IN19[17], w1547, w1548);
  FullAdder U323 (w1548, w1511, IN20[17], w1549, w1550);
  FullAdder U324 (w1550, w1513, IN21[15], w1551, w1552);
  FullAdder U325 (w1552, w1515, IN22[14], w1553, w1554);
  FullAdder U326 (w1554, w1517, IN23[13], w1555, w1556);
  FullAdder U327 (w1556, w1519, IN24[12], w1557, w1558);
  FullAdder U328 (w1558, w1521, IN25[11], w1559, w1560);
  FullAdder U329 (w1560, w1523, IN26[10], w1561, w1562);
  FullAdder U330 (w1562, w1525, IN27[9], w1563, w1564);
  FullAdder U331 (w1564, w1527, IN28[8], w1565, w1566);
  FullAdder U332 (w1566, w1529, IN29[7], w1567, w1568);
  FullAdder U333 (w1568, w1531, IN30[6], w1569, w1570);
  FullAdder U334 (w1570, w1533, IN31[5], w1571, w1572);
  FullAdder U335 (w1572, w1535, IN32[4], w1573, w1574);
  FullAdder U336 (w1574, w1537, IN33[3], w1575, w1576);
  FullAdder U337 (w1576, w1539, IN34[2], w1577, w1578);
  FullAdder U338 (w1578, w1541, IN35[1], w1579, w1580);
  FullAdder U339 (w1580, w1542, IN36[0], w1581, w1582);
  HalfAdder U340 (w1545, IN18[18], Out1[18], w1584);
  FullAdder U341 (w1584, w1547, IN19[18], w1585, w1586);
  FullAdder U342 (w1586, w1549, IN20[18], w1587, w1588);
  FullAdder U343 (w1588, w1551, IN21[16], w1589, w1590);
  FullAdder U344 (w1590, w1553, IN22[15], w1591, w1592);
  FullAdder U345 (w1592, w1555, IN23[14], w1593, w1594);
  FullAdder U346 (w1594, w1557, IN24[13], w1595, w1596);
  FullAdder U347 (w1596, w1559, IN25[12], w1597, w1598);
  FullAdder U348 (w1598, w1561, IN26[11], w1599, w1600);
  FullAdder U349 (w1600, w1563, IN27[10], w1601, w1602);
  FullAdder U350 (w1602, w1565, IN28[9], w1603, w1604);
  FullAdder U351 (w1604, w1567, IN29[8], w1605, w1606);
  FullAdder U352 (w1606, w1569, IN30[7], w1607, w1608);
  FullAdder U353 (w1608, w1571, IN31[6], w1609, w1610);
  FullAdder U354 (w1610, w1573, IN32[5], w1611, w1612);
  FullAdder U355 (w1612, w1575, IN33[4], w1613, w1614);
  FullAdder U356 (w1614, w1577, IN34[3], w1615, w1616);
  FullAdder U357 (w1616, w1579, IN35[2], w1617, w1618);
  FullAdder U358 (w1618, w1581, IN36[1], w1619, w1620);
  FullAdder U359 (w1620, w1582, IN37[0], w1621, w1622);
  HalfAdder U360 (w1585, IN19[19], Out1[19], w1624);
  FullAdder U361 (w1624, w1587, IN20[19], w1625, w1626);
  FullAdder U362 (w1626, w1589, IN21[17], w1627, w1628);
  FullAdder U363 (w1628, w1591, IN22[16], w1629, w1630);
  FullAdder U364 (w1630, w1593, IN23[15], w1631, w1632);
  FullAdder U365 (w1632, w1595, IN24[14], w1633, w1634);
  FullAdder U366 (w1634, w1597, IN25[13], w1635, w1636);
  FullAdder U367 (w1636, w1599, IN26[12], w1637, w1638);
  FullAdder U368 (w1638, w1601, IN27[11], w1639, w1640);
  FullAdder U369 (w1640, w1603, IN28[10], w1641, w1642);
  FullAdder U370 (w1642, w1605, IN29[9], w1643, w1644);
  FullAdder U371 (w1644, w1607, IN30[8], w1645, w1646);
  FullAdder U372 (w1646, w1609, IN31[7], w1647, w1648);
  FullAdder U373 (w1648, w1611, IN32[6], w1649, w1650);
  FullAdder U374 (w1650, w1613, IN33[5], w1651, w1652);
  FullAdder U375 (w1652, w1615, IN34[4], w1653, w1654);
  FullAdder U376 (w1654, w1617, IN35[3], w1655, w1656);
  FullAdder U377 (w1656, w1619, IN36[2], w1657, w1658);
  FullAdder U378 (w1658, w1621, IN37[1], w1659, w1660);
  FullAdder U379 (w1660, w1622, IN38[0], w1661, w1662);
  HalfAdder U380 (w1625, IN20[20], Out1[20], w1664);
  FullAdder U381 (w1664, w1627, IN21[18], w1665, w1666);
  FullAdder U382 (w1666, w1629, IN22[17], w1667, w1668);
  FullAdder U383 (w1668, w1631, IN23[16], w1669, w1670);
  FullAdder U384 (w1670, w1633, IN24[15], w1671, w1672);
  FullAdder U385 (w1672, w1635, IN25[14], w1673, w1674);
  FullAdder U386 (w1674, w1637, IN26[13], w1675, w1676);
  FullAdder U387 (w1676, w1639, IN27[12], w1677, w1678);
  FullAdder U388 (w1678, w1641, IN28[11], w1679, w1680);
  FullAdder U389 (w1680, w1643, IN29[10], w1681, w1682);
  FullAdder U390 (w1682, w1645, IN30[9], w1683, w1684);
  FullAdder U391 (w1684, w1647, IN31[8], w1685, w1686);
  FullAdder U392 (w1686, w1649, IN32[7], w1687, w1688);
  FullAdder U393 (w1688, w1651, IN33[6], w1689, w1690);
  FullAdder U394 (w1690, w1653, IN34[5], w1691, w1692);
  FullAdder U395 (w1692, w1655, IN35[4], w1693, w1694);
  FullAdder U396 (w1694, w1657, IN36[3], w1695, w1696);
  FullAdder U397 (w1696, w1659, IN37[2], w1697, w1698);
  FullAdder U398 (w1698, w1661, IN38[1], w1699, w1700);
  FullAdder U399 (w1700, w1662, IN39[0], w1701, w1702);
  HalfAdder U400 (w1665, IN21[19], Out1[21], w1704);
  FullAdder U401 (w1704, w1667, IN22[18], w1705, w1706);
  FullAdder U402 (w1706, w1669, IN23[17], w1707, w1708);
  FullAdder U403 (w1708, w1671, IN24[16], w1709, w1710);
  FullAdder U404 (w1710, w1673, IN25[15], w1711, w1712);
  FullAdder U405 (w1712, w1675, IN26[14], w1713, w1714);
  FullAdder U406 (w1714, w1677, IN27[13], w1715, w1716);
  FullAdder U407 (w1716, w1679, IN28[12], w1717, w1718);
  FullAdder U408 (w1718, w1681, IN29[11], w1719, w1720);
  FullAdder U409 (w1720, w1683, IN30[10], w1721, w1722);
  FullAdder U410 (w1722, w1685, IN31[9], w1723, w1724);
  FullAdder U411 (w1724, w1687, IN32[8], w1725, w1726);
  FullAdder U412 (w1726, w1689, IN33[7], w1727, w1728);
  FullAdder U413 (w1728, w1691, IN34[6], w1729, w1730);
  FullAdder U414 (w1730, w1693, IN35[5], w1731, w1732);
  FullAdder U415 (w1732, w1695, IN36[4], w1733, w1734);
  FullAdder U416 (w1734, w1697, IN37[3], w1735, w1736);
  FullAdder U417 (w1736, w1699, IN38[2], w1737, w1738);
  FullAdder U418 (w1738, w1701, IN39[1], w1739, w1740);
  FullAdder U419 (w1740, w1702, IN40[0], w1741, w1742);
  HalfAdder U420 (w1705, IN22[19], Out1[22], w1744);
  FullAdder U421 (w1744, w1707, IN23[18], w1745, w1746);
  FullAdder U422 (w1746, w1709, IN24[17], w1747, w1748);
  FullAdder U423 (w1748, w1711, IN25[16], w1749, w1750);
  FullAdder U424 (w1750, w1713, IN26[15], w1751, w1752);
  FullAdder U425 (w1752, w1715, IN27[14], w1753, w1754);
  FullAdder U426 (w1754, w1717, IN28[13], w1755, w1756);
  FullAdder U427 (w1756, w1719, IN29[12], w1757, w1758);
  FullAdder U428 (w1758, w1721, IN30[11], w1759, w1760);
  FullAdder U429 (w1760, w1723, IN31[10], w1761, w1762);
  FullAdder U430 (w1762, w1725, IN32[9], w1763, w1764);
  FullAdder U431 (w1764, w1727, IN33[8], w1765, w1766);
  FullAdder U432 (w1766, w1729, IN34[7], w1767, w1768);
  FullAdder U433 (w1768, w1731, IN35[6], w1769, w1770);
  FullAdder U434 (w1770, w1733, IN36[5], w1771, w1772);
  FullAdder U435 (w1772, w1735, IN37[4], w1773, w1774);
  FullAdder U436 (w1774, w1737, IN38[3], w1775, w1776);
  FullAdder U437 (w1776, w1739, IN39[2], w1777, w1778);
  FullAdder U438 (w1778, w1741, IN40[1], w1779, w1780);
  FullAdder U439 (w1780, w1742, IN41[0], w1781, w1782);
  HalfAdder U440 (w1745, IN23[19], Out1[23], w1784);
  FullAdder U441 (w1784, w1747, IN24[18], w1785, w1786);
  FullAdder U442 (w1786, w1749, IN25[17], w1787, w1788);
  FullAdder U443 (w1788, w1751, IN26[16], w1789, w1790);
  FullAdder U444 (w1790, w1753, IN27[15], w1791, w1792);
  FullAdder U445 (w1792, w1755, IN28[14], w1793, w1794);
  FullAdder U446 (w1794, w1757, IN29[13], w1795, w1796);
  FullAdder U447 (w1796, w1759, IN30[12], w1797, w1798);
  FullAdder U448 (w1798, w1761, IN31[11], w1799, w1800);
  FullAdder U449 (w1800, w1763, IN32[10], w1801, w1802);
  FullAdder U450 (w1802, w1765, IN33[9], w1803, w1804);
  FullAdder U451 (w1804, w1767, IN34[8], w1805, w1806);
  FullAdder U452 (w1806, w1769, IN35[7], w1807, w1808);
  FullAdder U453 (w1808, w1771, IN36[6], w1809, w1810);
  FullAdder U454 (w1810, w1773, IN37[5], w1811, w1812);
  FullAdder U455 (w1812, w1775, IN38[4], w1813, w1814);
  FullAdder U456 (w1814, w1777, IN39[3], w1815, w1816);
  FullAdder U457 (w1816, w1779, IN40[2], w1817, w1818);
  FullAdder U458 (w1818, w1781, IN41[1], w1819, w1820);
  FullAdder U459 (w1820, w1782, IN42[0], w1821, w1822);
  HalfAdder U460 (w1785, IN24[19], Out1[24], w1824);
  FullAdder U461 (w1824, w1787, IN25[18], w1825, w1826);
  FullAdder U462 (w1826, w1789, IN26[17], w1827, w1828);
  FullAdder U463 (w1828, w1791, IN27[16], w1829, w1830);
  FullAdder U464 (w1830, w1793, IN28[15], w1831, w1832);
  FullAdder U465 (w1832, w1795, IN29[14], w1833, w1834);
  FullAdder U466 (w1834, w1797, IN30[13], w1835, w1836);
  FullAdder U467 (w1836, w1799, IN31[12], w1837, w1838);
  FullAdder U468 (w1838, w1801, IN32[11], w1839, w1840);
  FullAdder U469 (w1840, w1803, IN33[10], w1841, w1842);
  FullAdder U470 (w1842, w1805, IN34[9], w1843, w1844);
  FullAdder U471 (w1844, w1807, IN35[8], w1845, w1846);
  FullAdder U472 (w1846, w1809, IN36[7], w1847, w1848);
  FullAdder U473 (w1848, w1811, IN37[6], w1849, w1850);
  FullAdder U474 (w1850, w1813, IN38[5], w1851, w1852);
  FullAdder U475 (w1852, w1815, IN39[4], w1853, w1854);
  FullAdder U476 (w1854, w1817, IN40[3], w1855, w1856);
  FullAdder U477 (w1856, w1819, IN41[2], w1857, w1858);
  FullAdder U478 (w1858, w1821, IN42[1], w1859, w1860);
  FullAdder U479 (w1860, w1822, IN43[0], w1861, w1862);
  HalfAdder U480 (w1825, IN25[19], Out1[25], w1864);
  FullAdder U481 (w1864, w1827, IN26[18], w1865, w1866);
  FullAdder U482 (w1866, w1829, IN27[17], w1867, w1868);
  FullAdder U483 (w1868, w1831, IN28[16], w1869, w1870);
  FullAdder U484 (w1870, w1833, IN29[15], w1871, w1872);
  FullAdder U485 (w1872, w1835, IN30[14], w1873, w1874);
  FullAdder U486 (w1874, w1837, IN31[13], w1875, w1876);
  FullAdder U487 (w1876, w1839, IN32[12], w1877, w1878);
  FullAdder U488 (w1878, w1841, IN33[11], w1879, w1880);
  FullAdder U489 (w1880, w1843, IN34[10], w1881, w1882);
  FullAdder U490 (w1882, w1845, IN35[9], w1883, w1884);
  FullAdder U491 (w1884, w1847, IN36[8], w1885, w1886);
  FullAdder U492 (w1886, w1849, IN37[7], w1887, w1888);
  FullAdder U493 (w1888, w1851, IN38[6], w1889, w1890);
  FullAdder U494 (w1890, w1853, IN39[5], w1891, w1892);
  FullAdder U495 (w1892, w1855, IN40[4], w1893, w1894);
  FullAdder U496 (w1894, w1857, IN41[3], w1895, w1896);
  FullAdder U497 (w1896, w1859, IN42[2], w1897, w1898);
  FullAdder U498 (w1898, w1861, IN43[1], w1899, w1900);
  FullAdder U499 (w1900, w1862, IN44[0], w1901, w1902);
  HalfAdder U500 (w1865, IN26[19], Out1[26], w1904);
  FullAdder U501 (w1904, w1867, IN27[18], w1905, w1906);
  FullAdder U502 (w1906, w1869, IN28[17], w1907, w1908);
  FullAdder U503 (w1908, w1871, IN29[16], w1909, w1910);
  FullAdder U504 (w1910, w1873, IN30[15], w1911, w1912);
  FullAdder U505 (w1912, w1875, IN31[14], w1913, w1914);
  FullAdder U506 (w1914, w1877, IN32[13], w1915, w1916);
  FullAdder U507 (w1916, w1879, IN33[12], w1917, w1918);
  FullAdder U508 (w1918, w1881, IN34[11], w1919, w1920);
  FullAdder U509 (w1920, w1883, IN35[10], w1921, w1922);
  FullAdder U510 (w1922, w1885, IN36[9], w1923, w1924);
  FullAdder U511 (w1924, w1887, IN37[8], w1925, w1926);
  FullAdder U512 (w1926, w1889, IN38[7], w1927, w1928);
  FullAdder U513 (w1928, w1891, IN39[6], w1929, w1930);
  FullAdder U514 (w1930, w1893, IN40[5], w1931, w1932);
  FullAdder U515 (w1932, w1895, IN41[4], w1933, w1934);
  FullAdder U516 (w1934, w1897, IN42[3], w1935, w1936);
  FullAdder U517 (w1936, w1899, IN43[2], w1937, w1938);
  FullAdder U518 (w1938, w1901, IN44[1], w1939, w1940);
  FullAdder U519 (w1940, w1902, IN45[0], w1941, w1942);
  HalfAdder U520 (w1905, IN27[19], Out1[27], w1944);
  FullAdder U521 (w1944, w1907, IN28[18], w1945, w1946);
  FullAdder U522 (w1946, w1909, IN29[17], w1947, w1948);
  FullAdder U523 (w1948, w1911, IN30[16], w1949, w1950);
  FullAdder U524 (w1950, w1913, IN31[15], w1951, w1952);
  FullAdder U525 (w1952, w1915, IN32[14], w1953, w1954);
  FullAdder U526 (w1954, w1917, IN33[13], w1955, w1956);
  FullAdder U527 (w1956, w1919, IN34[12], w1957, w1958);
  FullAdder U528 (w1958, w1921, IN35[11], w1959, w1960);
  FullAdder U529 (w1960, w1923, IN36[10], w1961, w1962);
  FullAdder U530 (w1962, w1925, IN37[9], w1963, w1964);
  FullAdder U531 (w1964, w1927, IN38[8], w1965, w1966);
  FullAdder U532 (w1966, w1929, IN39[7], w1967, w1968);
  FullAdder U533 (w1968, w1931, IN40[6], w1969, w1970);
  FullAdder U534 (w1970, w1933, IN41[5], w1971, w1972);
  FullAdder U535 (w1972, w1935, IN42[4], w1973, w1974);
  FullAdder U536 (w1974, w1937, IN43[3], w1975, w1976);
  FullAdder U537 (w1976, w1939, IN44[2], w1977, w1978);
  FullAdder U538 (w1978, w1941, IN45[1], w1979, w1980);
  FullAdder U539 (w1980, w1942, IN46[0], w1981, w1982);
  HalfAdder U540 (w1945, IN28[19], Out1[28], w1984);
  FullAdder U541 (w1984, w1947, IN29[18], w1985, w1986);
  FullAdder U542 (w1986, w1949, IN30[17], w1987, w1988);
  FullAdder U543 (w1988, w1951, IN31[16], w1989, w1990);
  FullAdder U544 (w1990, w1953, IN32[15], w1991, w1992);
  FullAdder U545 (w1992, w1955, IN33[14], w1993, w1994);
  FullAdder U546 (w1994, w1957, IN34[13], w1995, w1996);
  FullAdder U547 (w1996, w1959, IN35[12], w1997, w1998);
  FullAdder U548 (w1998, w1961, IN36[11], w1999, w2000);
  FullAdder U549 (w2000, w1963, IN37[10], w2001, w2002);
  FullAdder U550 (w2002, w1965, IN38[9], w2003, w2004);
  FullAdder U551 (w2004, w1967, IN39[8], w2005, w2006);
  FullAdder U552 (w2006, w1969, IN40[7], w2007, w2008);
  FullAdder U553 (w2008, w1971, IN41[6], w2009, w2010);
  FullAdder U554 (w2010, w1973, IN42[5], w2011, w2012);
  FullAdder U555 (w2012, w1975, IN43[4], w2013, w2014);
  FullAdder U556 (w2014, w1977, IN44[3], w2015, w2016);
  FullAdder U557 (w2016, w1979, IN45[2], w2017, w2018);
  FullAdder U558 (w2018, w1981, IN46[1], w2019, w2020);
  FullAdder U559 (w2020, w1982, IN47[0], w2021, w2022);
  HalfAdder U560 (w1985, IN29[19], Out1[29], w2024);
  FullAdder U561 (w2024, w1987, IN30[18], w2025, w2026);
  FullAdder U562 (w2026, w1989, IN31[17], w2027, w2028);
  FullAdder U563 (w2028, w1991, IN32[16], w2029, w2030);
  FullAdder U564 (w2030, w1993, IN33[15], w2031, w2032);
  FullAdder U565 (w2032, w1995, IN34[14], w2033, w2034);
  FullAdder U566 (w2034, w1997, IN35[13], w2035, w2036);
  FullAdder U567 (w2036, w1999, IN36[12], w2037, w2038);
  FullAdder U568 (w2038, w2001, IN37[11], w2039, w2040);
  FullAdder U569 (w2040, w2003, IN38[10], w2041, w2042);
  FullAdder U570 (w2042, w2005, IN39[9], w2043, w2044);
  FullAdder U571 (w2044, w2007, IN40[8], w2045, w2046);
  FullAdder U572 (w2046, w2009, IN41[7], w2047, w2048);
  FullAdder U573 (w2048, w2011, IN42[6], w2049, w2050);
  FullAdder U574 (w2050, w2013, IN43[5], w2051, w2052);
  FullAdder U575 (w2052, w2015, IN44[4], w2053, w2054);
  FullAdder U576 (w2054, w2017, IN45[3], w2055, w2056);
  FullAdder U577 (w2056, w2019, IN46[2], w2057, w2058);
  FullAdder U578 (w2058, w2021, IN47[1], w2059, w2060);
  FullAdder U579 (w2060, w2022, IN48[0], w2061, w2062);
  HalfAdder U580 (w2025, IN30[19], Out1[30], w2064);
  FullAdder U581 (w2064, w2027, IN31[18], w2065, w2066);
  FullAdder U582 (w2066, w2029, IN32[17], w2067, w2068);
  FullAdder U583 (w2068, w2031, IN33[16], w2069, w2070);
  FullAdder U584 (w2070, w2033, IN34[15], w2071, w2072);
  FullAdder U585 (w2072, w2035, IN35[14], w2073, w2074);
  FullAdder U586 (w2074, w2037, IN36[13], w2075, w2076);
  FullAdder U587 (w2076, w2039, IN37[12], w2077, w2078);
  FullAdder U588 (w2078, w2041, IN38[11], w2079, w2080);
  FullAdder U589 (w2080, w2043, IN39[10], w2081, w2082);
  FullAdder U590 (w2082, w2045, IN40[9], w2083, w2084);
  FullAdder U591 (w2084, w2047, IN41[8], w2085, w2086);
  FullAdder U592 (w2086, w2049, IN42[7], w2087, w2088);
  FullAdder U593 (w2088, w2051, IN43[6], w2089, w2090);
  FullAdder U594 (w2090, w2053, IN44[5], w2091, w2092);
  FullAdder U595 (w2092, w2055, IN45[4], w2093, w2094);
  FullAdder U596 (w2094, w2057, IN46[3], w2095, w2096);
  FullAdder U597 (w2096, w2059, IN47[2], w2097, w2098);
  FullAdder U598 (w2098, w2061, IN48[1], w2099, w2100);
  FullAdder U599 (w2100, w2062, IN49[0], w2101, w2102);
  HalfAdder U600 (w2065, IN31[19], Out1[31], w2104);
  FullAdder U601 (w2104, w2067, IN32[18], w2105, w2106);
  FullAdder U602 (w2106, w2069, IN33[17], w2107, w2108);
  FullAdder U603 (w2108, w2071, IN34[16], w2109, w2110);
  FullAdder U604 (w2110, w2073, IN35[15], w2111, w2112);
  FullAdder U605 (w2112, w2075, IN36[14], w2113, w2114);
  FullAdder U606 (w2114, w2077, IN37[13], w2115, w2116);
  FullAdder U607 (w2116, w2079, IN38[12], w2117, w2118);
  FullAdder U608 (w2118, w2081, IN39[11], w2119, w2120);
  FullAdder U609 (w2120, w2083, IN40[10], w2121, w2122);
  FullAdder U610 (w2122, w2085, IN41[9], w2123, w2124);
  FullAdder U611 (w2124, w2087, IN42[8], w2125, w2126);
  FullAdder U612 (w2126, w2089, IN43[7], w2127, w2128);
  FullAdder U613 (w2128, w2091, IN44[6], w2129, w2130);
  FullAdder U614 (w2130, w2093, IN45[5], w2131, w2132);
  FullAdder U615 (w2132, w2095, IN46[4], w2133, w2134);
  FullAdder U616 (w2134, w2097, IN47[3], w2135, w2136);
  FullAdder U617 (w2136, w2099, IN48[2], w2137, w2138);
  FullAdder U618 (w2138, w2101, IN49[1], w2139, w2140);
  FullAdder U619 (w2140, w2102, IN50[0], w2141, w2142);
  HalfAdder U620 (w2105, IN32[19], Out1[32], w2144);
  FullAdder U621 (w2144, w2107, IN33[18], w2145, w2146);
  FullAdder U622 (w2146, w2109, IN34[17], w2147, w2148);
  FullAdder U623 (w2148, w2111, IN35[16], w2149, w2150);
  FullAdder U624 (w2150, w2113, IN36[15], w2151, w2152);
  FullAdder U625 (w2152, w2115, IN37[14], w2153, w2154);
  FullAdder U626 (w2154, w2117, IN38[13], w2155, w2156);
  FullAdder U627 (w2156, w2119, IN39[12], w2157, w2158);
  FullAdder U628 (w2158, w2121, IN40[11], w2159, w2160);
  FullAdder U629 (w2160, w2123, IN41[10], w2161, w2162);
  FullAdder U630 (w2162, w2125, IN42[9], w2163, w2164);
  FullAdder U631 (w2164, w2127, IN43[8], w2165, w2166);
  FullAdder U632 (w2166, w2129, IN44[7], w2167, w2168);
  FullAdder U633 (w2168, w2131, IN45[6], w2169, w2170);
  FullAdder U634 (w2170, w2133, IN46[5], w2171, w2172);
  FullAdder U635 (w2172, w2135, IN47[4], w2173, w2174);
  FullAdder U636 (w2174, w2137, IN48[3], w2175, w2176);
  FullAdder U637 (w2176, w2139, IN49[2], w2177, w2178);
  FullAdder U638 (w2178, w2141, IN50[1], w2179, w2180);
  FullAdder U639 (w2180, w2142, IN51[0], w2181, w2182);
  HalfAdder U640 (w2145, IN33[19], Out1[33], w2184);
  FullAdder U641 (w2184, w2147, IN34[18], w2185, w2186);
  FullAdder U642 (w2186, w2149, IN35[17], w2187, w2188);
  FullAdder U643 (w2188, w2151, IN36[16], w2189, w2190);
  FullAdder U644 (w2190, w2153, IN37[15], w2191, w2192);
  FullAdder U645 (w2192, w2155, IN38[14], w2193, w2194);
  FullAdder U646 (w2194, w2157, IN39[13], w2195, w2196);
  FullAdder U647 (w2196, w2159, IN40[12], w2197, w2198);
  FullAdder U648 (w2198, w2161, IN41[11], w2199, w2200);
  FullAdder U649 (w2200, w2163, IN42[10], w2201, w2202);
  FullAdder U650 (w2202, w2165, IN43[9], w2203, w2204);
  FullAdder U651 (w2204, w2167, IN44[8], w2205, w2206);
  FullAdder U652 (w2206, w2169, IN45[7], w2207, w2208);
  FullAdder U653 (w2208, w2171, IN46[6], w2209, w2210);
  FullAdder U654 (w2210, w2173, IN47[5], w2211, w2212);
  FullAdder U655 (w2212, w2175, IN48[4], w2213, w2214);
  FullAdder U656 (w2214, w2177, IN49[3], w2215, w2216);
  FullAdder U657 (w2216, w2179, IN50[2], w2217, w2218);
  FullAdder U658 (w2218, w2181, IN51[1], w2219, w2220);
  FullAdder U659 (w2220, w2182, IN52[0], w2221, w2222);
  HalfAdder U660 (w2185, IN34[19], Out1[34], w2224);
  FullAdder U661 (w2224, w2187, IN35[18], w2225, w2226);
  FullAdder U662 (w2226, w2189, IN36[17], w2227, w2228);
  FullAdder U663 (w2228, w2191, IN37[16], w2229, w2230);
  FullAdder U664 (w2230, w2193, IN38[15], w2231, w2232);
  FullAdder U665 (w2232, w2195, IN39[14], w2233, w2234);
  FullAdder U666 (w2234, w2197, IN40[13], w2235, w2236);
  FullAdder U667 (w2236, w2199, IN41[12], w2237, w2238);
  FullAdder U668 (w2238, w2201, IN42[11], w2239, w2240);
  FullAdder U669 (w2240, w2203, IN43[10], w2241, w2242);
  FullAdder U670 (w2242, w2205, IN44[9], w2243, w2244);
  FullAdder U671 (w2244, w2207, IN45[8], w2245, w2246);
  FullAdder U672 (w2246, w2209, IN46[7], w2247, w2248);
  FullAdder U673 (w2248, w2211, IN47[6], w2249, w2250);
  FullAdder U674 (w2250, w2213, IN48[5], w2251, w2252);
  FullAdder U675 (w2252, w2215, IN49[4], w2253, w2254);
  FullAdder U676 (w2254, w2217, IN50[3], w2255, w2256);
  FullAdder U677 (w2256, w2219, IN51[2], w2257, w2258);
  FullAdder U678 (w2258, w2221, IN52[1], w2259, w2260);
  FullAdder U679 (w2260, w2222, IN53[0], w2261, w2262);
  HalfAdder U680 (w2225, IN35[19], Out1[35], w2264);
  FullAdder U681 (w2264, w2227, IN36[18], w2265, w2266);
  FullAdder U682 (w2266, w2229, IN37[17], w2267, w2268);
  FullAdder U683 (w2268, w2231, IN38[16], w2269, w2270);
  FullAdder U684 (w2270, w2233, IN39[15], w2271, w2272);
  FullAdder U685 (w2272, w2235, IN40[14], w2273, w2274);
  FullAdder U686 (w2274, w2237, IN41[13], w2275, w2276);
  FullAdder U687 (w2276, w2239, IN42[12], w2277, w2278);
  FullAdder U688 (w2278, w2241, IN43[11], w2279, w2280);
  FullAdder U689 (w2280, w2243, IN44[10], w2281, w2282);
  FullAdder U690 (w2282, w2245, IN45[9], w2283, w2284);
  FullAdder U691 (w2284, w2247, IN46[8], w2285, w2286);
  FullAdder U692 (w2286, w2249, IN47[7], w2287, w2288);
  FullAdder U693 (w2288, w2251, IN48[6], w2289, w2290);
  FullAdder U694 (w2290, w2253, IN49[5], w2291, w2292);
  FullAdder U695 (w2292, w2255, IN50[4], w2293, w2294);
  FullAdder U696 (w2294, w2257, IN51[3], w2295, w2296);
  FullAdder U697 (w2296, w2259, IN52[2], w2297, w2298);
  FullAdder U698 (w2298, w2261, IN53[1], w2299, w2300);
  FullAdder U699 (w2300, w2262, IN54[0], w2301, w2302);
  HalfAdder U700 (w2265, IN36[19], Out1[36], w2304);
  FullAdder U701 (w2304, w2267, IN37[18], w2305, w2306);
  FullAdder U702 (w2306, w2269, IN38[17], w2307, w2308);
  FullAdder U703 (w2308, w2271, IN39[16], w2309, w2310);
  FullAdder U704 (w2310, w2273, IN40[15], w2311, w2312);
  FullAdder U705 (w2312, w2275, IN41[14], w2313, w2314);
  FullAdder U706 (w2314, w2277, IN42[13], w2315, w2316);
  FullAdder U707 (w2316, w2279, IN43[12], w2317, w2318);
  FullAdder U708 (w2318, w2281, IN44[11], w2319, w2320);
  FullAdder U709 (w2320, w2283, IN45[10], w2321, w2322);
  FullAdder U710 (w2322, w2285, IN46[9], w2323, w2324);
  FullAdder U711 (w2324, w2287, IN47[8], w2325, w2326);
  FullAdder U712 (w2326, w2289, IN48[7], w2327, w2328);
  FullAdder U713 (w2328, w2291, IN49[6], w2329, w2330);
  FullAdder U714 (w2330, w2293, IN50[5], w2331, w2332);
  FullAdder U715 (w2332, w2295, IN51[4], w2333, w2334);
  FullAdder U716 (w2334, w2297, IN52[3], w2335, w2336);
  FullAdder U717 (w2336, w2299, IN53[2], w2337, w2338);
  FullAdder U718 (w2338, w2301, IN54[1], w2339, w2340);
  FullAdder U719 (w2340, w2302, IN55[0], w2341, w2342);
  HalfAdder U720 (w2305, IN37[19], Out1[37], w2344);
  FullAdder U721 (w2344, w2307, IN38[18], w2345, w2346);
  FullAdder U722 (w2346, w2309, IN39[17], w2347, w2348);
  FullAdder U723 (w2348, w2311, IN40[16], w2349, w2350);
  FullAdder U724 (w2350, w2313, IN41[15], w2351, w2352);
  FullAdder U725 (w2352, w2315, IN42[14], w2353, w2354);
  FullAdder U726 (w2354, w2317, IN43[13], w2355, w2356);
  FullAdder U727 (w2356, w2319, IN44[12], w2357, w2358);
  FullAdder U728 (w2358, w2321, IN45[11], w2359, w2360);
  FullAdder U729 (w2360, w2323, IN46[10], w2361, w2362);
  FullAdder U730 (w2362, w2325, IN47[9], w2363, w2364);
  FullAdder U731 (w2364, w2327, IN48[8], w2365, w2366);
  FullAdder U732 (w2366, w2329, IN49[7], w2367, w2368);
  FullAdder U733 (w2368, w2331, IN50[6], w2369, w2370);
  FullAdder U734 (w2370, w2333, IN51[5], w2371, w2372);
  FullAdder U735 (w2372, w2335, IN52[4], w2373, w2374);
  FullAdder U736 (w2374, w2337, IN53[3], w2375, w2376);
  FullAdder U737 (w2376, w2339, IN54[2], w2377, w2378);
  FullAdder U738 (w2378, w2341, IN55[1], w2379, w2380);
  FullAdder U739 (w2380, w2342, IN56[0], w2381, w2382);
  HalfAdder U740 (w2345, IN38[19], Out1[38], w2384);
  FullAdder U741 (w2384, w2347, IN39[18], w2385, w2386);
  FullAdder U742 (w2386, w2349, IN40[17], w2387, w2388);
  FullAdder U743 (w2388, w2351, IN41[16], w2389, w2390);
  FullAdder U744 (w2390, w2353, IN42[15], w2391, w2392);
  FullAdder U745 (w2392, w2355, IN43[14], w2393, w2394);
  FullAdder U746 (w2394, w2357, IN44[13], w2395, w2396);
  FullAdder U747 (w2396, w2359, IN45[12], w2397, w2398);
  FullAdder U748 (w2398, w2361, IN46[11], w2399, w2400);
  FullAdder U749 (w2400, w2363, IN47[10], w2401, w2402);
  FullAdder U750 (w2402, w2365, IN48[9], w2403, w2404);
  FullAdder U751 (w2404, w2367, IN49[8], w2405, w2406);
  FullAdder U752 (w2406, w2369, IN50[7], w2407, w2408);
  FullAdder U753 (w2408, w2371, IN51[6], w2409, w2410);
  FullAdder U754 (w2410, w2373, IN52[5], w2411, w2412);
  FullAdder U755 (w2412, w2375, IN53[4], w2413, w2414);
  FullAdder U756 (w2414, w2377, IN54[3], w2415, w2416);
  FullAdder U757 (w2416, w2379, IN55[2], w2417, w2418);
  FullAdder U758 (w2418, w2381, IN56[1], w2419, w2420);
  FullAdder U759 (w2420, w2382, IN57[0], w2421, w2422);
  HalfAdder U760 (w2385, IN39[19], Out1[39], w2424);
  FullAdder U761 (w2424, w2387, IN40[18], w2425, w2426);
  FullAdder U762 (w2426, w2389, IN41[17], w2427, w2428);
  FullAdder U763 (w2428, w2391, IN42[16], w2429, w2430);
  FullAdder U764 (w2430, w2393, IN43[15], w2431, w2432);
  FullAdder U765 (w2432, w2395, IN44[14], w2433, w2434);
  FullAdder U766 (w2434, w2397, IN45[13], w2435, w2436);
  FullAdder U767 (w2436, w2399, IN46[12], w2437, w2438);
  FullAdder U768 (w2438, w2401, IN47[11], w2439, w2440);
  FullAdder U769 (w2440, w2403, IN48[10], w2441, w2442);
  FullAdder U770 (w2442, w2405, IN49[9], w2443, w2444);
  FullAdder U771 (w2444, w2407, IN50[8], w2445, w2446);
  FullAdder U772 (w2446, w2409, IN51[7], w2447, w2448);
  FullAdder U773 (w2448, w2411, IN52[6], w2449, w2450);
  FullAdder U774 (w2450, w2413, IN53[5], w2451, w2452);
  FullAdder U775 (w2452, w2415, IN54[4], w2453, w2454);
  FullAdder U776 (w2454, w2417, IN55[3], w2455, w2456);
  FullAdder U777 (w2456, w2419, IN56[2], w2457, w2458);
  FullAdder U778 (w2458, w2421, IN57[1], w2459, w2460);
  FullAdder U779 (w2460, w2422, IN58[0], w2461, w2462);
  HalfAdder U780 (w2425, IN40[19], Out1[40], w2464);
  FullAdder U781 (w2464, w2427, IN41[18], w2465, w2466);
  FullAdder U782 (w2466, w2429, IN42[17], w2467, w2468);
  FullAdder U783 (w2468, w2431, IN43[16], w2469, w2470);
  FullAdder U784 (w2470, w2433, IN44[15], w2471, w2472);
  FullAdder U785 (w2472, w2435, IN45[14], w2473, w2474);
  FullAdder U786 (w2474, w2437, IN46[13], w2475, w2476);
  FullAdder U787 (w2476, w2439, IN47[12], w2477, w2478);
  FullAdder U788 (w2478, w2441, IN48[11], w2479, w2480);
  FullAdder U789 (w2480, w2443, IN49[10], w2481, w2482);
  FullAdder U790 (w2482, w2445, IN50[9], w2483, w2484);
  FullAdder U791 (w2484, w2447, IN51[8], w2485, w2486);
  FullAdder U792 (w2486, w2449, IN52[7], w2487, w2488);
  FullAdder U793 (w2488, w2451, IN53[6], w2489, w2490);
  FullAdder U794 (w2490, w2453, IN54[5], w2491, w2492);
  FullAdder U795 (w2492, w2455, IN55[4], w2493, w2494);
  FullAdder U796 (w2494, w2457, IN56[3], w2495, w2496);
  FullAdder U797 (w2496, w2459, IN57[2], w2497, w2498);
  FullAdder U798 (w2498, w2461, IN58[1], w2499, w2500);
  FullAdder U799 (w2500, w2462, IN59[0], w2501, w2502);
  HalfAdder U800 (w2465, IN41[19], Out1[41], w2504);
  FullAdder U801 (w2504, w2467, IN42[18], w2505, w2506);
  FullAdder U802 (w2506, w2469, IN43[17], w2507, w2508);
  FullAdder U803 (w2508, w2471, IN44[16], w2509, w2510);
  FullAdder U804 (w2510, w2473, IN45[15], w2511, w2512);
  FullAdder U805 (w2512, w2475, IN46[14], w2513, w2514);
  FullAdder U806 (w2514, w2477, IN47[13], w2515, w2516);
  FullAdder U807 (w2516, w2479, IN48[12], w2517, w2518);
  FullAdder U808 (w2518, w2481, IN49[11], w2519, w2520);
  FullAdder U809 (w2520, w2483, IN50[10], w2521, w2522);
  FullAdder U810 (w2522, w2485, IN51[9], w2523, w2524);
  FullAdder U811 (w2524, w2487, IN52[8], w2525, w2526);
  FullAdder U812 (w2526, w2489, IN53[7], w2527, w2528);
  FullAdder U813 (w2528, w2491, IN54[6], w2529, w2530);
  FullAdder U814 (w2530, w2493, IN55[5], w2531, w2532);
  FullAdder U815 (w2532, w2495, IN56[4], w2533, w2534);
  FullAdder U816 (w2534, w2497, IN57[3], w2535, w2536);
  FullAdder U817 (w2536, w2499, IN58[2], w2537, w2538);
  FullAdder U818 (w2538, w2501, IN59[1], w2539, w2540);
  FullAdder U819 (w2540, w2502, IN60[0], w2541, w2542);
  HalfAdder U820 (w2505, IN42[19], Out1[42], w2544);
  FullAdder U821 (w2544, w2507, IN43[18], Out1[43], w2546);
  FullAdder U822 (w2546, w2509, IN44[17], Out1[44], w2548);
  FullAdder U823 (w2548, w2511, IN45[16], Out1[45], w2550);
  FullAdder U824 (w2550, w2513, IN46[15], Out1[46], w2552);
  FullAdder U825 (w2552, w2515, IN47[14], Out1[47], w2554);
  FullAdder U826 (w2554, w2517, IN48[13], Out1[48], w2556);
  FullAdder U827 (w2556, w2519, IN49[12], Out1[49], w2558);
  FullAdder U828 (w2558, w2521, IN50[11], Out1[50], w2560);
  FullAdder U829 (w2560, w2523, IN51[10], Out1[51], w2562);
  FullAdder U830 (w2562, w2525, IN52[9], Out1[52], w2564);
  FullAdder U831 (w2564, w2527, IN53[8], Out1[53], w2566);
  FullAdder U832 (w2566, w2529, IN54[7], Out1[54], w2568);
  FullAdder U833 (w2568, w2531, IN55[6], Out1[55], w2570);
  FullAdder U834 (w2570, w2533, IN56[5], Out1[56], w2572);
  FullAdder U835 (w2572, w2535, IN57[4], Out1[57], w2574);
  FullAdder U836 (w2574, w2537, IN58[3], Out1[58], w2576);
  FullAdder U837 (w2576, w2539, IN59[2], Out1[59], w2578);
  FullAdder U838 (w2578, w2541, IN60[1], Out1[60], w2580);
  FullAdder U839 (w2580, w2542, IN61[0], Out1[61], Out1[62]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN21[20];
  assign Out2[1] = IN22[20];
  assign Out2[2] = IN23[20];
  assign Out2[3] = IN24[20];
  assign Out2[4] = IN25[20];
  assign Out2[5] = IN26[20];
  assign Out2[6] = IN27[20];
  assign Out2[7] = IN28[20];
  assign Out2[8] = IN29[20];
  assign Out2[9] = IN30[20];
  assign Out2[10] = IN31[20];
  assign Out2[11] = IN32[20];
  assign Out2[12] = IN33[20];
  assign Out2[13] = IN34[20];
  assign Out2[14] = IN35[20];
  assign Out2[15] = IN36[20];
  assign Out2[16] = IN37[20];
  assign Out2[17] = IN38[20];
  assign Out2[18] = IN39[20];
  assign Out2[19] = IN40[20];
  assign Out2[20] = IN41[20];
  assign Out2[21] = IN42[20];
  assign Out2[22] = IN43[19];
  assign Out2[23] = IN44[18];
  assign Out2[24] = IN45[17];
  assign Out2[25] = IN46[16];
  assign Out2[26] = IN47[15];
  assign Out2[27] = IN48[14];
  assign Out2[28] = IN49[13];
  assign Out2[29] = IN50[12];
  assign Out2[30] = IN51[11];
  assign Out2[31] = IN52[10];
  assign Out2[32] = IN53[9];
  assign Out2[33] = IN54[8];
  assign Out2[34] = IN55[7];
  assign Out2[35] = IN56[6];
  assign Out2[36] = IN57[5];
  assign Out2[37] = IN58[4];
  assign Out2[38] = IN59[3];
  assign Out2[39] = IN60[2];
  assign Out2[40] = IN61[1];
  assign Out2[41] = IN62[0];

endmodule
module RC_42_42(IN1, IN2, Out);
  input [41:0] IN1;
  input [41:0] IN2;
  output [42:0] Out;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w85);
  FullAdder U1 (IN1[1], IN2[1], w85, Out[1], w87);
  FullAdder U2 (IN1[2], IN2[2], w87, Out[2], w89);
  FullAdder U3 (IN1[3], IN2[3], w89, Out[3], w91);
  FullAdder U4 (IN1[4], IN2[4], w91, Out[4], w93);
  FullAdder U5 (IN1[5], IN2[5], w93, Out[5], w95);
  FullAdder U6 (IN1[6], IN2[6], w95, Out[6], w97);
  FullAdder U7 (IN1[7], IN2[7], w97, Out[7], w99);
  FullAdder U8 (IN1[8], IN2[8], w99, Out[8], w101);
  FullAdder U9 (IN1[9], IN2[9], w101, Out[9], w103);
  FullAdder U10 (IN1[10], IN2[10], w103, Out[10], w105);
  FullAdder U11 (IN1[11], IN2[11], w105, Out[11], w107);
  FullAdder U12 (IN1[12], IN2[12], w107, Out[12], w109);
  FullAdder U13 (IN1[13], IN2[13], w109, Out[13], w111);
  FullAdder U14 (IN1[14], IN2[14], w111, Out[14], w113);
  FullAdder U15 (IN1[15], IN2[15], w113, Out[15], w115);
  FullAdder U16 (IN1[16], IN2[16], w115, Out[16], w117);
  FullAdder U17 (IN1[17], IN2[17], w117, Out[17], w119);
  FullAdder U18 (IN1[18], IN2[18], w119, Out[18], w121);
  FullAdder U19 (IN1[19], IN2[19], w121, Out[19], w123);
  FullAdder U20 (IN1[20], IN2[20], w123, Out[20], w125);
  FullAdder U21 (IN1[21], IN2[21], w125, Out[21], w127);
  FullAdder U22 (IN1[22], IN2[22], w127, Out[22], w129);
  FullAdder U23 (IN1[23], IN2[23], w129, Out[23], w131);
  FullAdder U24 (IN1[24], IN2[24], w131, Out[24], w133);
  FullAdder U25 (IN1[25], IN2[25], w133, Out[25], w135);
  FullAdder U26 (IN1[26], IN2[26], w135, Out[26], w137);
  FullAdder U27 (IN1[27], IN2[27], w137, Out[27], w139);
  FullAdder U28 (IN1[28], IN2[28], w139, Out[28], w141);
  FullAdder U29 (IN1[29], IN2[29], w141, Out[29], w143);
  FullAdder U30 (IN1[30], IN2[30], w143, Out[30], w145);
  FullAdder U31 (IN1[31], IN2[31], w145, Out[31], w147);
  FullAdder U32 (IN1[32], IN2[32], w147, Out[32], w149);
  FullAdder U33 (IN1[33], IN2[33], w149, Out[33], w151);
  FullAdder U34 (IN1[34], IN2[34], w151, Out[34], w153);
  FullAdder U35 (IN1[35], IN2[35], w153, Out[35], w155);
  FullAdder U36 (IN1[36], IN2[36], w155, Out[36], w157);
  FullAdder U37 (IN1[37], IN2[37], w157, Out[37], w159);
  FullAdder U38 (IN1[38], IN2[38], w159, Out[38], w161);
  FullAdder U39 (IN1[39], IN2[39], w161, Out[39], w163);
  FullAdder U40 (IN1[40], IN2[40], w163, Out[40], w165);
  FullAdder U41 (IN1[41], IN2[41], w165, Out[41], Out[42]);

endmodule
module NR_21_43(IN1, IN2, Out);
  input [20:0] IN1;
  input [42:0] IN2;
  output [63:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [20:0] P21;
  wire [20:0] P22;
  wire [20:0] P23;
  wire [20:0] P24;
  wire [20:0] P25;
  wire [20:0] P26;
  wire [20:0] P27;
  wire [20:0] P28;
  wire [20:0] P29;
  wire [20:0] P30;
  wire [20:0] P31;
  wire [20:0] P32;
  wire [20:0] P33;
  wire [20:0] P34;
  wire [20:0] P35;
  wire [20:0] P36;
  wire [20:0] P37;
  wire [20:0] P38;
  wire [20:0] P39;
  wire [20:0] P40;
  wire [20:0] P41;
  wire [20:0] P42;
  wire [19:0] P43;
  wire [18:0] P44;
  wire [17:0] P45;
  wire [16:0] P46;
  wire [15:0] P47;
  wire [14:0] P48;
  wire [13:0] P49;
  wire [12:0] P50;
  wire [11:0] P51;
  wire [10:0] P52;
  wire [9:0] P53;
  wire [8:0] P54;
  wire [7:0] P55;
  wire [6:0] P56;
  wire [5:0] P57;
  wire [4:0] P58;
  wire [3:0] P59;
  wire [2:0] P60;
  wire [1:0] P61;
  wire [0:0] P62;
  wire [62:0] R1;
  wire [41:0] R2;
  wire [63:0] aOut;
  U_SP_21_43 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, R1, R2);
  RC_42_42 S2 (R1[62:21], R2, aOut[63:21]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign Out = aOut[63:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
