
module customAdder57_0(
    input [56 : 0] A,
    input [56 : 0] B,
    output [57 : 0] Sum
);

    assign Sum = A+B;

endmodule
