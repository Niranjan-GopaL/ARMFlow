//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 46
  second input length: 25
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_46_25(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69);
  input [45:0] IN1;
  input [24:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [24:0] P25;
  output [24:0] P26;
  output [24:0] P27;
  output [24:0] P28;
  output [24:0] P29;
  output [24:0] P30;
  output [24:0] P31;
  output [24:0] P32;
  output [24:0] P33;
  output [24:0] P34;
  output [24:0] P35;
  output [24:0] P36;
  output [24:0] P37;
  output [24:0] P38;
  output [24:0] P39;
  output [24:0] P40;
  output [24:0] P41;
  output [24:0] P42;
  output [24:0] P43;
  output [24:0] P44;
  output [24:0] P45;
  output [23:0] P46;
  output [22:0] P47;
  output [21:0] P48;
  output [20:0] P49;
  output [19:0] P50;
  output [18:0] P51;
  output [17:0] P52;
  output [16:0] P53;
  output [15:0] P54;
  output [14:0] P55;
  output [13:0] P56;
  output [12:0] P57;
  output [11:0] P58;
  output [10:0] P59;
  output [9:0] P60;
  output [8:0] P61;
  output [7:0] P62;
  output [6:0] P63;
  output [5:0] P64;
  output [4:0] P65;
  output [3:0] P66;
  output [2:0] P67;
  output [1:0] P68;
  output [0:0] P69;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[0] = IN1[1]&IN2[24];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[1] = IN1[2]&IN2[23];
  assign P26[0] = IN1[2]&IN2[24];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[2] = IN1[3]&IN2[22];
  assign P26[1] = IN1[3]&IN2[23];
  assign P27[0] = IN1[3]&IN2[24];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[3] = IN1[4]&IN2[21];
  assign P26[2] = IN1[4]&IN2[22];
  assign P27[1] = IN1[4]&IN2[23];
  assign P28[0] = IN1[4]&IN2[24];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[4] = IN1[5]&IN2[20];
  assign P26[3] = IN1[5]&IN2[21];
  assign P27[2] = IN1[5]&IN2[22];
  assign P28[1] = IN1[5]&IN2[23];
  assign P29[0] = IN1[5]&IN2[24];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[5] = IN1[6]&IN2[19];
  assign P26[4] = IN1[6]&IN2[20];
  assign P27[3] = IN1[6]&IN2[21];
  assign P28[2] = IN1[6]&IN2[22];
  assign P29[1] = IN1[6]&IN2[23];
  assign P30[0] = IN1[6]&IN2[24];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[6] = IN1[7]&IN2[18];
  assign P26[5] = IN1[7]&IN2[19];
  assign P27[4] = IN1[7]&IN2[20];
  assign P28[3] = IN1[7]&IN2[21];
  assign P29[2] = IN1[7]&IN2[22];
  assign P30[1] = IN1[7]&IN2[23];
  assign P31[0] = IN1[7]&IN2[24];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[7] = IN1[8]&IN2[17];
  assign P26[6] = IN1[8]&IN2[18];
  assign P27[5] = IN1[8]&IN2[19];
  assign P28[4] = IN1[8]&IN2[20];
  assign P29[3] = IN1[8]&IN2[21];
  assign P30[2] = IN1[8]&IN2[22];
  assign P31[1] = IN1[8]&IN2[23];
  assign P32[0] = IN1[8]&IN2[24];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[8] = IN1[9]&IN2[16];
  assign P26[7] = IN1[9]&IN2[17];
  assign P27[6] = IN1[9]&IN2[18];
  assign P28[5] = IN1[9]&IN2[19];
  assign P29[4] = IN1[9]&IN2[20];
  assign P30[3] = IN1[9]&IN2[21];
  assign P31[2] = IN1[9]&IN2[22];
  assign P32[1] = IN1[9]&IN2[23];
  assign P33[0] = IN1[9]&IN2[24];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[9] = IN1[10]&IN2[15];
  assign P26[8] = IN1[10]&IN2[16];
  assign P27[7] = IN1[10]&IN2[17];
  assign P28[6] = IN1[10]&IN2[18];
  assign P29[5] = IN1[10]&IN2[19];
  assign P30[4] = IN1[10]&IN2[20];
  assign P31[3] = IN1[10]&IN2[21];
  assign P32[2] = IN1[10]&IN2[22];
  assign P33[1] = IN1[10]&IN2[23];
  assign P34[0] = IN1[10]&IN2[24];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[10] = IN1[11]&IN2[14];
  assign P26[9] = IN1[11]&IN2[15];
  assign P27[8] = IN1[11]&IN2[16];
  assign P28[7] = IN1[11]&IN2[17];
  assign P29[6] = IN1[11]&IN2[18];
  assign P30[5] = IN1[11]&IN2[19];
  assign P31[4] = IN1[11]&IN2[20];
  assign P32[3] = IN1[11]&IN2[21];
  assign P33[2] = IN1[11]&IN2[22];
  assign P34[1] = IN1[11]&IN2[23];
  assign P35[0] = IN1[11]&IN2[24];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[11] = IN1[12]&IN2[13];
  assign P26[10] = IN1[12]&IN2[14];
  assign P27[9] = IN1[12]&IN2[15];
  assign P28[8] = IN1[12]&IN2[16];
  assign P29[7] = IN1[12]&IN2[17];
  assign P30[6] = IN1[12]&IN2[18];
  assign P31[5] = IN1[12]&IN2[19];
  assign P32[4] = IN1[12]&IN2[20];
  assign P33[3] = IN1[12]&IN2[21];
  assign P34[2] = IN1[12]&IN2[22];
  assign P35[1] = IN1[12]&IN2[23];
  assign P36[0] = IN1[12]&IN2[24];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[12] = IN1[13]&IN2[12];
  assign P26[11] = IN1[13]&IN2[13];
  assign P27[10] = IN1[13]&IN2[14];
  assign P28[9] = IN1[13]&IN2[15];
  assign P29[8] = IN1[13]&IN2[16];
  assign P30[7] = IN1[13]&IN2[17];
  assign P31[6] = IN1[13]&IN2[18];
  assign P32[5] = IN1[13]&IN2[19];
  assign P33[4] = IN1[13]&IN2[20];
  assign P34[3] = IN1[13]&IN2[21];
  assign P35[2] = IN1[13]&IN2[22];
  assign P36[1] = IN1[13]&IN2[23];
  assign P37[0] = IN1[13]&IN2[24];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[13] = IN1[14]&IN2[11];
  assign P26[12] = IN1[14]&IN2[12];
  assign P27[11] = IN1[14]&IN2[13];
  assign P28[10] = IN1[14]&IN2[14];
  assign P29[9] = IN1[14]&IN2[15];
  assign P30[8] = IN1[14]&IN2[16];
  assign P31[7] = IN1[14]&IN2[17];
  assign P32[6] = IN1[14]&IN2[18];
  assign P33[5] = IN1[14]&IN2[19];
  assign P34[4] = IN1[14]&IN2[20];
  assign P35[3] = IN1[14]&IN2[21];
  assign P36[2] = IN1[14]&IN2[22];
  assign P37[1] = IN1[14]&IN2[23];
  assign P38[0] = IN1[14]&IN2[24];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[14] = IN1[15]&IN2[10];
  assign P26[13] = IN1[15]&IN2[11];
  assign P27[12] = IN1[15]&IN2[12];
  assign P28[11] = IN1[15]&IN2[13];
  assign P29[10] = IN1[15]&IN2[14];
  assign P30[9] = IN1[15]&IN2[15];
  assign P31[8] = IN1[15]&IN2[16];
  assign P32[7] = IN1[15]&IN2[17];
  assign P33[6] = IN1[15]&IN2[18];
  assign P34[5] = IN1[15]&IN2[19];
  assign P35[4] = IN1[15]&IN2[20];
  assign P36[3] = IN1[15]&IN2[21];
  assign P37[2] = IN1[15]&IN2[22];
  assign P38[1] = IN1[15]&IN2[23];
  assign P39[0] = IN1[15]&IN2[24];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[15] = IN1[16]&IN2[9];
  assign P26[14] = IN1[16]&IN2[10];
  assign P27[13] = IN1[16]&IN2[11];
  assign P28[12] = IN1[16]&IN2[12];
  assign P29[11] = IN1[16]&IN2[13];
  assign P30[10] = IN1[16]&IN2[14];
  assign P31[9] = IN1[16]&IN2[15];
  assign P32[8] = IN1[16]&IN2[16];
  assign P33[7] = IN1[16]&IN2[17];
  assign P34[6] = IN1[16]&IN2[18];
  assign P35[5] = IN1[16]&IN2[19];
  assign P36[4] = IN1[16]&IN2[20];
  assign P37[3] = IN1[16]&IN2[21];
  assign P38[2] = IN1[16]&IN2[22];
  assign P39[1] = IN1[16]&IN2[23];
  assign P40[0] = IN1[16]&IN2[24];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[16] = IN1[17]&IN2[8];
  assign P26[15] = IN1[17]&IN2[9];
  assign P27[14] = IN1[17]&IN2[10];
  assign P28[13] = IN1[17]&IN2[11];
  assign P29[12] = IN1[17]&IN2[12];
  assign P30[11] = IN1[17]&IN2[13];
  assign P31[10] = IN1[17]&IN2[14];
  assign P32[9] = IN1[17]&IN2[15];
  assign P33[8] = IN1[17]&IN2[16];
  assign P34[7] = IN1[17]&IN2[17];
  assign P35[6] = IN1[17]&IN2[18];
  assign P36[5] = IN1[17]&IN2[19];
  assign P37[4] = IN1[17]&IN2[20];
  assign P38[3] = IN1[17]&IN2[21];
  assign P39[2] = IN1[17]&IN2[22];
  assign P40[1] = IN1[17]&IN2[23];
  assign P41[0] = IN1[17]&IN2[24];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[17] = IN1[18]&IN2[7];
  assign P26[16] = IN1[18]&IN2[8];
  assign P27[15] = IN1[18]&IN2[9];
  assign P28[14] = IN1[18]&IN2[10];
  assign P29[13] = IN1[18]&IN2[11];
  assign P30[12] = IN1[18]&IN2[12];
  assign P31[11] = IN1[18]&IN2[13];
  assign P32[10] = IN1[18]&IN2[14];
  assign P33[9] = IN1[18]&IN2[15];
  assign P34[8] = IN1[18]&IN2[16];
  assign P35[7] = IN1[18]&IN2[17];
  assign P36[6] = IN1[18]&IN2[18];
  assign P37[5] = IN1[18]&IN2[19];
  assign P38[4] = IN1[18]&IN2[20];
  assign P39[3] = IN1[18]&IN2[21];
  assign P40[2] = IN1[18]&IN2[22];
  assign P41[1] = IN1[18]&IN2[23];
  assign P42[0] = IN1[18]&IN2[24];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[18] = IN1[19]&IN2[6];
  assign P26[17] = IN1[19]&IN2[7];
  assign P27[16] = IN1[19]&IN2[8];
  assign P28[15] = IN1[19]&IN2[9];
  assign P29[14] = IN1[19]&IN2[10];
  assign P30[13] = IN1[19]&IN2[11];
  assign P31[12] = IN1[19]&IN2[12];
  assign P32[11] = IN1[19]&IN2[13];
  assign P33[10] = IN1[19]&IN2[14];
  assign P34[9] = IN1[19]&IN2[15];
  assign P35[8] = IN1[19]&IN2[16];
  assign P36[7] = IN1[19]&IN2[17];
  assign P37[6] = IN1[19]&IN2[18];
  assign P38[5] = IN1[19]&IN2[19];
  assign P39[4] = IN1[19]&IN2[20];
  assign P40[3] = IN1[19]&IN2[21];
  assign P41[2] = IN1[19]&IN2[22];
  assign P42[1] = IN1[19]&IN2[23];
  assign P43[0] = IN1[19]&IN2[24];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[19] = IN1[20]&IN2[5];
  assign P26[18] = IN1[20]&IN2[6];
  assign P27[17] = IN1[20]&IN2[7];
  assign P28[16] = IN1[20]&IN2[8];
  assign P29[15] = IN1[20]&IN2[9];
  assign P30[14] = IN1[20]&IN2[10];
  assign P31[13] = IN1[20]&IN2[11];
  assign P32[12] = IN1[20]&IN2[12];
  assign P33[11] = IN1[20]&IN2[13];
  assign P34[10] = IN1[20]&IN2[14];
  assign P35[9] = IN1[20]&IN2[15];
  assign P36[8] = IN1[20]&IN2[16];
  assign P37[7] = IN1[20]&IN2[17];
  assign P38[6] = IN1[20]&IN2[18];
  assign P39[5] = IN1[20]&IN2[19];
  assign P40[4] = IN1[20]&IN2[20];
  assign P41[3] = IN1[20]&IN2[21];
  assign P42[2] = IN1[20]&IN2[22];
  assign P43[1] = IN1[20]&IN2[23];
  assign P44[0] = IN1[20]&IN2[24];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[20] = IN1[21]&IN2[4];
  assign P26[19] = IN1[21]&IN2[5];
  assign P27[18] = IN1[21]&IN2[6];
  assign P28[17] = IN1[21]&IN2[7];
  assign P29[16] = IN1[21]&IN2[8];
  assign P30[15] = IN1[21]&IN2[9];
  assign P31[14] = IN1[21]&IN2[10];
  assign P32[13] = IN1[21]&IN2[11];
  assign P33[12] = IN1[21]&IN2[12];
  assign P34[11] = IN1[21]&IN2[13];
  assign P35[10] = IN1[21]&IN2[14];
  assign P36[9] = IN1[21]&IN2[15];
  assign P37[8] = IN1[21]&IN2[16];
  assign P38[7] = IN1[21]&IN2[17];
  assign P39[6] = IN1[21]&IN2[18];
  assign P40[5] = IN1[21]&IN2[19];
  assign P41[4] = IN1[21]&IN2[20];
  assign P42[3] = IN1[21]&IN2[21];
  assign P43[2] = IN1[21]&IN2[22];
  assign P44[1] = IN1[21]&IN2[23];
  assign P45[0] = IN1[21]&IN2[24];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[21] = IN1[22]&IN2[3];
  assign P26[20] = IN1[22]&IN2[4];
  assign P27[19] = IN1[22]&IN2[5];
  assign P28[18] = IN1[22]&IN2[6];
  assign P29[17] = IN1[22]&IN2[7];
  assign P30[16] = IN1[22]&IN2[8];
  assign P31[15] = IN1[22]&IN2[9];
  assign P32[14] = IN1[22]&IN2[10];
  assign P33[13] = IN1[22]&IN2[11];
  assign P34[12] = IN1[22]&IN2[12];
  assign P35[11] = IN1[22]&IN2[13];
  assign P36[10] = IN1[22]&IN2[14];
  assign P37[9] = IN1[22]&IN2[15];
  assign P38[8] = IN1[22]&IN2[16];
  assign P39[7] = IN1[22]&IN2[17];
  assign P40[6] = IN1[22]&IN2[18];
  assign P41[5] = IN1[22]&IN2[19];
  assign P42[4] = IN1[22]&IN2[20];
  assign P43[3] = IN1[22]&IN2[21];
  assign P44[2] = IN1[22]&IN2[22];
  assign P45[1] = IN1[22]&IN2[23];
  assign P46[0] = IN1[22]&IN2[24];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[22] = IN1[23]&IN2[2];
  assign P26[21] = IN1[23]&IN2[3];
  assign P27[20] = IN1[23]&IN2[4];
  assign P28[19] = IN1[23]&IN2[5];
  assign P29[18] = IN1[23]&IN2[6];
  assign P30[17] = IN1[23]&IN2[7];
  assign P31[16] = IN1[23]&IN2[8];
  assign P32[15] = IN1[23]&IN2[9];
  assign P33[14] = IN1[23]&IN2[10];
  assign P34[13] = IN1[23]&IN2[11];
  assign P35[12] = IN1[23]&IN2[12];
  assign P36[11] = IN1[23]&IN2[13];
  assign P37[10] = IN1[23]&IN2[14];
  assign P38[9] = IN1[23]&IN2[15];
  assign P39[8] = IN1[23]&IN2[16];
  assign P40[7] = IN1[23]&IN2[17];
  assign P41[6] = IN1[23]&IN2[18];
  assign P42[5] = IN1[23]&IN2[19];
  assign P43[4] = IN1[23]&IN2[20];
  assign P44[3] = IN1[23]&IN2[21];
  assign P45[2] = IN1[23]&IN2[22];
  assign P46[1] = IN1[23]&IN2[23];
  assign P47[0] = IN1[23]&IN2[24];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[23] = IN1[24]&IN2[1];
  assign P26[22] = IN1[24]&IN2[2];
  assign P27[21] = IN1[24]&IN2[3];
  assign P28[20] = IN1[24]&IN2[4];
  assign P29[19] = IN1[24]&IN2[5];
  assign P30[18] = IN1[24]&IN2[6];
  assign P31[17] = IN1[24]&IN2[7];
  assign P32[16] = IN1[24]&IN2[8];
  assign P33[15] = IN1[24]&IN2[9];
  assign P34[14] = IN1[24]&IN2[10];
  assign P35[13] = IN1[24]&IN2[11];
  assign P36[12] = IN1[24]&IN2[12];
  assign P37[11] = IN1[24]&IN2[13];
  assign P38[10] = IN1[24]&IN2[14];
  assign P39[9] = IN1[24]&IN2[15];
  assign P40[8] = IN1[24]&IN2[16];
  assign P41[7] = IN1[24]&IN2[17];
  assign P42[6] = IN1[24]&IN2[18];
  assign P43[5] = IN1[24]&IN2[19];
  assign P44[4] = IN1[24]&IN2[20];
  assign P45[3] = IN1[24]&IN2[21];
  assign P46[2] = IN1[24]&IN2[22];
  assign P47[1] = IN1[24]&IN2[23];
  assign P48[0] = IN1[24]&IN2[24];
  assign P25[24] = IN1[25]&IN2[0];
  assign P26[23] = IN1[25]&IN2[1];
  assign P27[22] = IN1[25]&IN2[2];
  assign P28[21] = IN1[25]&IN2[3];
  assign P29[20] = IN1[25]&IN2[4];
  assign P30[19] = IN1[25]&IN2[5];
  assign P31[18] = IN1[25]&IN2[6];
  assign P32[17] = IN1[25]&IN2[7];
  assign P33[16] = IN1[25]&IN2[8];
  assign P34[15] = IN1[25]&IN2[9];
  assign P35[14] = IN1[25]&IN2[10];
  assign P36[13] = IN1[25]&IN2[11];
  assign P37[12] = IN1[25]&IN2[12];
  assign P38[11] = IN1[25]&IN2[13];
  assign P39[10] = IN1[25]&IN2[14];
  assign P40[9] = IN1[25]&IN2[15];
  assign P41[8] = IN1[25]&IN2[16];
  assign P42[7] = IN1[25]&IN2[17];
  assign P43[6] = IN1[25]&IN2[18];
  assign P44[5] = IN1[25]&IN2[19];
  assign P45[4] = IN1[25]&IN2[20];
  assign P46[3] = IN1[25]&IN2[21];
  assign P47[2] = IN1[25]&IN2[22];
  assign P48[1] = IN1[25]&IN2[23];
  assign P49[0] = IN1[25]&IN2[24];
  assign P26[24] = IN1[26]&IN2[0];
  assign P27[23] = IN1[26]&IN2[1];
  assign P28[22] = IN1[26]&IN2[2];
  assign P29[21] = IN1[26]&IN2[3];
  assign P30[20] = IN1[26]&IN2[4];
  assign P31[19] = IN1[26]&IN2[5];
  assign P32[18] = IN1[26]&IN2[6];
  assign P33[17] = IN1[26]&IN2[7];
  assign P34[16] = IN1[26]&IN2[8];
  assign P35[15] = IN1[26]&IN2[9];
  assign P36[14] = IN1[26]&IN2[10];
  assign P37[13] = IN1[26]&IN2[11];
  assign P38[12] = IN1[26]&IN2[12];
  assign P39[11] = IN1[26]&IN2[13];
  assign P40[10] = IN1[26]&IN2[14];
  assign P41[9] = IN1[26]&IN2[15];
  assign P42[8] = IN1[26]&IN2[16];
  assign P43[7] = IN1[26]&IN2[17];
  assign P44[6] = IN1[26]&IN2[18];
  assign P45[5] = IN1[26]&IN2[19];
  assign P46[4] = IN1[26]&IN2[20];
  assign P47[3] = IN1[26]&IN2[21];
  assign P48[2] = IN1[26]&IN2[22];
  assign P49[1] = IN1[26]&IN2[23];
  assign P50[0] = IN1[26]&IN2[24];
  assign P27[24] = IN1[27]&IN2[0];
  assign P28[23] = IN1[27]&IN2[1];
  assign P29[22] = IN1[27]&IN2[2];
  assign P30[21] = IN1[27]&IN2[3];
  assign P31[20] = IN1[27]&IN2[4];
  assign P32[19] = IN1[27]&IN2[5];
  assign P33[18] = IN1[27]&IN2[6];
  assign P34[17] = IN1[27]&IN2[7];
  assign P35[16] = IN1[27]&IN2[8];
  assign P36[15] = IN1[27]&IN2[9];
  assign P37[14] = IN1[27]&IN2[10];
  assign P38[13] = IN1[27]&IN2[11];
  assign P39[12] = IN1[27]&IN2[12];
  assign P40[11] = IN1[27]&IN2[13];
  assign P41[10] = IN1[27]&IN2[14];
  assign P42[9] = IN1[27]&IN2[15];
  assign P43[8] = IN1[27]&IN2[16];
  assign P44[7] = IN1[27]&IN2[17];
  assign P45[6] = IN1[27]&IN2[18];
  assign P46[5] = IN1[27]&IN2[19];
  assign P47[4] = IN1[27]&IN2[20];
  assign P48[3] = IN1[27]&IN2[21];
  assign P49[2] = IN1[27]&IN2[22];
  assign P50[1] = IN1[27]&IN2[23];
  assign P51[0] = IN1[27]&IN2[24];
  assign P28[24] = IN1[28]&IN2[0];
  assign P29[23] = IN1[28]&IN2[1];
  assign P30[22] = IN1[28]&IN2[2];
  assign P31[21] = IN1[28]&IN2[3];
  assign P32[20] = IN1[28]&IN2[4];
  assign P33[19] = IN1[28]&IN2[5];
  assign P34[18] = IN1[28]&IN2[6];
  assign P35[17] = IN1[28]&IN2[7];
  assign P36[16] = IN1[28]&IN2[8];
  assign P37[15] = IN1[28]&IN2[9];
  assign P38[14] = IN1[28]&IN2[10];
  assign P39[13] = IN1[28]&IN2[11];
  assign P40[12] = IN1[28]&IN2[12];
  assign P41[11] = IN1[28]&IN2[13];
  assign P42[10] = IN1[28]&IN2[14];
  assign P43[9] = IN1[28]&IN2[15];
  assign P44[8] = IN1[28]&IN2[16];
  assign P45[7] = IN1[28]&IN2[17];
  assign P46[6] = IN1[28]&IN2[18];
  assign P47[5] = IN1[28]&IN2[19];
  assign P48[4] = IN1[28]&IN2[20];
  assign P49[3] = IN1[28]&IN2[21];
  assign P50[2] = IN1[28]&IN2[22];
  assign P51[1] = IN1[28]&IN2[23];
  assign P52[0] = IN1[28]&IN2[24];
  assign P29[24] = IN1[29]&IN2[0];
  assign P30[23] = IN1[29]&IN2[1];
  assign P31[22] = IN1[29]&IN2[2];
  assign P32[21] = IN1[29]&IN2[3];
  assign P33[20] = IN1[29]&IN2[4];
  assign P34[19] = IN1[29]&IN2[5];
  assign P35[18] = IN1[29]&IN2[6];
  assign P36[17] = IN1[29]&IN2[7];
  assign P37[16] = IN1[29]&IN2[8];
  assign P38[15] = IN1[29]&IN2[9];
  assign P39[14] = IN1[29]&IN2[10];
  assign P40[13] = IN1[29]&IN2[11];
  assign P41[12] = IN1[29]&IN2[12];
  assign P42[11] = IN1[29]&IN2[13];
  assign P43[10] = IN1[29]&IN2[14];
  assign P44[9] = IN1[29]&IN2[15];
  assign P45[8] = IN1[29]&IN2[16];
  assign P46[7] = IN1[29]&IN2[17];
  assign P47[6] = IN1[29]&IN2[18];
  assign P48[5] = IN1[29]&IN2[19];
  assign P49[4] = IN1[29]&IN2[20];
  assign P50[3] = IN1[29]&IN2[21];
  assign P51[2] = IN1[29]&IN2[22];
  assign P52[1] = IN1[29]&IN2[23];
  assign P53[0] = IN1[29]&IN2[24];
  assign P30[24] = IN1[30]&IN2[0];
  assign P31[23] = IN1[30]&IN2[1];
  assign P32[22] = IN1[30]&IN2[2];
  assign P33[21] = IN1[30]&IN2[3];
  assign P34[20] = IN1[30]&IN2[4];
  assign P35[19] = IN1[30]&IN2[5];
  assign P36[18] = IN1[30]&IN2[6];
  assign P37[17] = IN1[30]&IN2[7];
  assign P38[16] = IN1[30]&IN2[8];
  assign P39[15] = IN1[30]&IN2[9];
  assign P40[14] = IN1[30]&IN2[10];
  assign P41[13] = IN1[30]&IN2[11];
  assign P42[12] = IN1[30]&IN2[12];
  assign P43[11] = IN1[30]&IN2[13];
  assign P44[10] = IN1[30]&IN2[14];
  assign P45[9] = IN1[30]&IN2[15];
  assign P46[8] = IN1[30]&IN2[16];
  assign P47[7] = IN1[30]&IN2[17];
  assign P48[6] = IN1[30]&IN2[18];
  assign P49[5] = IN1[30]&IN2[19];
  assign P50[4] = IN1[30]&IN2[20];
  assign P51[3] = IN1[30]&IN2[21];
  assign P52[2] = IN1[30]&IN2[22];
  assign P53[1] = IN1[30]&IN2[23];
  assign P54[0] = IN1[30]&IN2[24];
  assign P31[24] = IN1[31]&IN2[0];
  assign P32[23] = IN1[31]&IN2[1];
  assign P33[22] = IN1[31]&IN2[2];
  assign P34[21] = IN1[31]&IN2[3];
  assign P35[20] = IN1[31]&IN2[4];
  assign P36[19] = IN1[31]&IN2[5];
  assign P37[18] = IN1[31]&IN2[6];
  assign P38[17] = IN1[31]&IN2[7];
  assign P39[16] = IN1[31]&IN2[8];
  assign P40[15] = IN1[31]&IN2[9];
  assign P41[14] = IN1[31]&IN2[10];
  assign P42[13] = IN1[31]&IN2[11];
  assign P43[12] = IN1[31]&IN2[12];
  assign P44[11] = IN1[31]&IN2[13];
  assign P45[10] = IN1[31]&IN2[14];
  assign P46[9] = IN1[31]&IN2[15];
  assign P47[8] = IN1[31]&IN2[16];
  assign P48[7] = IN1[31]&IN2[17];
  assign P49[6] = IN1[31]&IN2[18];
  assign P50[5] = IN1[31]&IN2[19];
  assign P51[4] = IN1[31]&IN2[20];
  assign P52[3] = IN1[31]&IN2[21];
  assign P53[2] = IN1[31]&IN2[22];
  assign P54[1] = IN1[31]&IN2[23];
  assign P55[0] = IN1[31]&IN2[24];
  assign P32[24] = IN1[32]&IN2[0];
  assign P33[23] = IN1[32]&IN2[1];
  assign P34[22] = IN1[32]&IN2[2];
  assign P35[21] = IN1[32]&IN2[3];
  assign P36[20] = IN1[32]&IN2[4];
  assign P37[19] = IN1[32]&IN2[5];
  assign P38[18] = IN1[32]&IN2[6];
  assign P39[17] = IN1[32]&IN2[7];
  assign P40[16] = IN1[32]&IN2[8];
  assign P41[15] = IN1[32]&IN2[9];
  assign P42[14] = IN1[32]&IN2[10];
  assign P43[13] = IN1[32]&IN2[11];
  assign P44[12] = IN1[32]&IN2[12];
  assign P45[11] = IN1[32]&IN2[13];
  assign P46[10] = IN1[32]&IN2[14];
  assign P47[9] = IN1[32]&IN2[15];
  assign P48[8] = IN1[32]&IN2[16];
  assign P49[7] = IN1[32]&IN2[17];
  assign P50[6] = IN1[32]&IN2[18];
  assign P51[5] = IN1[32]&IN2[19];
  assign P52[4] = IN1[32]&IN2[20];
  assign P53[3] = IN1[32]&IN2[21];
  assign P54[2] = IN1[32]&IN2[22];
  assign P55[1] = IN1[32]&IN2[23];
  assign P56[0] = IN1[32]&IN2[24];
  assign P33[24] = IN1[33]&IN2[0];
  assign P34[23] = IN1[33]&IN2[1];
  assign P35[22] = IN1[33]&IN2[2];
  assign P36[21] = IN1[33]&IN2[3];
  assign P37[20] = IN1[33]&IN2[4];
  assign P38[19] = IN1[33]&IN2[5];
  assign P39[18] = IN1[33]&IN2[6];
  assign P40[17] = IN1[33]&IN2[7];
  assign P41[16] = IN1[33]&IN2[8];
  assign P42[15] = IN1[33]&IN2[9];
  assign P43[14] = IN1[33]&IN2[10];
  assign P44[13] = IN1[33]&IN2[11];
  assign P45[12] = IN1[33]&IN2[12];
  assign P46[11] = IN1[33]&IN2[13];
  assign P47[10] = IN1[33]&IN2[14];
  assign P48[9] = IN1[33]&IN2[15];
  assign P49[8] = IN1[33]&IN2[16];
  assign P50[7] = IN1[33]&IN2[17];
  assign P51[6] = IN1[33]&IN2[18];
  assign P52[5] = IN1[33]&IN2[19];
  assign P53[4] = IN1[33]&IN2[20];
  assign P54[3] = IN1[33]&IN2[21];
  assign P55[2] = IN1[33]&IN2[22];
  assign P56[1] = IN1[33]&IN2[23];
  assign P57[0] = IN1[33]&IN2[24];
  assign P34[24] = IN1[34]&IN2[0];
  assign P35[23] = IN1[34]&IN2[1];
  assign P36[22] = IN1[34]&IN2[2];
  assign P37[21] = IN1[34]&IN2[3];
  assign P38[20] = IN1[34]&IN2[4];
  assign P39[19] = IN1[34]&IN2[5];
  assign P40[18] = IN1[34]&IN2[6];
  assign P41[17] = IN1[34]&IN2[7];
  assign P42[16] = IN1[34]&IN2[8];
  assign P43[15] = IN1[34]&IN2[9];
  assign P44[14] = IN1[34]&IN2[10];
  assign P45[13] = IN1[34]&IN2[11];
  assign P46[12] = IN1[34]&IN2[12];
  assign P47[11] = IN1[34]&IN2[13];
  assign P48[10] = IN1[34]&IN2[14];
  assign P49[9] = IN1[34]&IN2[15];
  assign P50[8] = IN1[34]&IN2[16];
  assign P51[7] = IN1[34]&IN2[17];
  assign P52[6] = IN1[34]&IN2[18];
  assign P53[5] = IN1[34]&IN2[19];
  assign P54[4] = IN1[34]&IN2[20];
  assign P55[3] = IN1[34]&IN2[21];
  assign P56[2] = IN1[34]&IN2[22];
  assign P57[1] = IN1[34]&IN2[23];
  assign P58[0] = IN1[34]&IN2[24];
  assign P35[24] = IN1[35]&IN2[0];
  assign P36[23] = IN1[35]&IN2[1];
  assign P37[22] = IN1[35]&IN2[2];
  assign P38[21] = IN1[35]&IN2[3];
  assign P39[20] = IN1[35]&IN2[4];
  assign P40[19] = IN1[35]&IN2[5];
  assign P41[18] = IN1[35]&IN2[6];
  assign P42[17] = IN1[35]&IN2[7];
  assign P43[16] = IN1[35]&IN2[8];
  assign P44[15] = IN1[35]&IN2[9];
  assign P45[14] = IN1[35]&IN2[10];
  assign P46[13] = IN1[35]&IN2[11];
  assign P47[12] = IN1[35]&IN2[12];
  assign P48[11] = IN1[35]&IN2[13];
  assign P49[10] = IN1[35]&IN2[14];
  assign P50[9] = IN1[35]&IN2[15];
  assign P51[8] = IN1[35]&IN2[16];
  assign P52[7] = IN1[35]&IN2[17];
  assign P53[6] = IN1[35]&IN2[18];
  assign P54[5] = IN1[35]&IN2[19];
  assign P55[4] = IN1[35]&IN2[20];
  assign P56[3] = IN1[35]&IN2[21];
  assign P57[2] = IN1[35]&IN2[22];
  assign P58[1] = IN1[35]&IN2[23];
  assign P59[0] = IN1[35]&IN2[24];
  assign P36[24] = IN1[36]&IN2[0];
  assign P37[23] = IN1[36]&IN2[1];
  assign P38[22] = IN1[36]&IN2[2];
  assign P39[21] = IN1[36]&IN2[3];
  assign P40[20] = IN1[36]&IN2[4];
  assign P41[19] = IN1[36]&IN2[5];
  assign P42[18] = IN1[36]&IN2[6];
  assign P43[17] = IN1[36]&IN2[7];
  assign P44[16] = IN1[36]&IN2[8];
  assign P45[15] = IN1[36]&IN2[9];
  assign P46[14] = IN1[36]&IN2[10];
  assign P47[13] = IN1[36]&IN2[11];
  assign P48[12] = IN1[36]&IN2[12];
  assign P49[11] = IN1[36]&IN2[13];
  assign P50[10] = IN1[36]&IN2[14];
  assign P51[9] = IN1[36]&IN2[15];
  assign P52[8] = IN1[36]&IN2[16];
  assign P53[7] = IN1[36]&IN2[17];
  assign P54[6] = IN1[36]&IN2[18];
  assign P55[5] = IN1[36]&IN2[19];
  assign P56[4] = IN1[36]&IN2[20];
  assign P57[3] = IN1[36]&IN2[21];
  assign P58[2] = IN1[36]&IN2[22];
  assign P59[1] = IN1[36]&IN2[23];
  assign P60[0] = IN1[36]&IN2[24];
  assign P37[24] = IN1[37]&IN2[0];
  assign P38[23] = IN1[37]&IN2[1];
  assign P39[22] = IN1[37]&IN2[2];
  assign P40[21] = IN1[37]&IN2[3];
  assign P41[20] = IN1[37]&IN2[4];
  assign P42[19] = IN1[37]&IN2[5];
  assign P43[18] = IN1[37]&IN2[6];
  assign P44[17] = IN1[37]&IN2[7];
  assign P45[16] = IN1[37]&IN2[8];
  assign P46[15] = IN1[37]&IN2[9];
  assign P47[14] = IN1[37]&IN2[10];
  assign P48[13] = IN1[37]&IN2[11];
  assign P49[12] = IN1[37]&IN2[12];
  assign P50[11] = IN1[37]&IN2[13];
  assign P51[10] = IN1[37]&IN2[14];
  assign P52[9] = IN1[37]&IN2[15];
  assign P53[8] = IN1[37]&IN2[16];
  assign P54[7] = IN1[37]&IN2[17];
  assign P55[6] = IN1[37]&IN2[18];
  assign P56[5] = IN1[37]&IN2[19];
  assign P57[4] = IN1[37]&IN2[20];
  assign P58[3] = IN1[37]&IN2[21];
  assign P59[2] = IN1[37]&IN2[22];
  assign P60[1] = IN1[37]&IN2[23];
  assign P61[0] = IN1[37]&IN2[24];
  assign P38[24] = IN1[38]&IN2[0];
  assign P39[23] = IN1[38]&IN2[1];
  assign P40[22] = IN1[38]&IN2[2];
  assign P41[21] = IN1[38]&IN2[3];
  assign P42[20] = IN1[38]&IN2[4];
  assign P43[19] = IN1[38]&IN2[5];
  assign P44[18] = IN1[38]&IN2[6];
  assign P45[17] = IN1[38]&IN2[7];
  assign P46[16] = IN1[38]&IN2[8];
  assign P47[15] = IN1[38]&IN2[9];
  assign P48[14] = IN1[38]&IN2[10];
  assign P49[13] = IN1[38]&IN2[11];
  assign P50[12] = IN1[38]&IN2[12];
  assign P51[11] = IN1[38]&IN2[13];
  assign P52[10] = IN1[38]&IN2[14];
  assign P53[9] = IN1[38]&IN2[15];
  assign P54[8] = IN1[38]&IN2[16];
  assign P55[7] = IN1[38]&IN2[17];
  assign P56[6] = IN1[38]&IN2[18];
  assign P57[5] = IN1[38]&IN2[19];
  assign P58[4] = IN1[38]&IN2[20];
  assign P59[3] = IN1[38]&IN2[21];
  assign P60[2] = IN1[38]&IN2[22];
  assign P61[1] = IN1[38]&IN2[23];
  assign P62[0] = IN1[38]&IN2[24];
  assign P39[24] = IN1[39]&IN2[0];
  assign P40[23] = IN1[39]&IN2[1];
  assign P41[22] = IN1[39]&IN2[2];
  assign P42[21] = IN1[39]&IN2[3];
  assign P43[20] = IN1[39]&IN2[4];
  assign P44[19] = IN1[39]&IN2[5];
  assign P45[18] = IN1[39]&IN2[6];
  assign P46[17] = IN1[39]&IN2[7];
  assign P47[16] = IN1[39]&IN2[8];
  assign P48[15] = IN1[39]&IN2[9];
  assign P49[14] = IN1[39]&IN2[10];
  assign P50[13] = IN1[39]&IN2[11];
  assign P51[12] = IN1[39]&IN2[12];
  assign P52[11] = IN1[39]&IN2[13];
  assign P53[10] = IN1[39]&IN2[14];
  assign P54[9] = IN1[39]&IN2[15];
  assign P55[8] = IN1[39]&IN2[16];
  assign P56[7] = IN1[39]&IN2[17];
  assign P57[6] = IN1[39]&IN2[18];
  assign P58[5] = IN1[39]&IN2[19];
  assign P59[4] = IN1[39]&IN2[20];
  assign P60[3] = IN1[39]&IN2[21];
  assign P61[2] = IN1[39]&IN2[22];
  assign P62[1] = IN1[39]&IN2[23];
  assign P63[0] = IN1[39]&IN2[24];
  assign P40[24] = IN1[40]&IN2[0];
  assign P41[23] = IN1[40]&IN2[1];
  assign P42[22] = IN1[40]&IN2[2];
  assign P43[21] = IN1[40]&IN2[3];
  assign P44[20] = IN1[40]&IN2[4];
  assign P45[19] = IN1[40]&IN2[5];
  assign P46[18] = IN1[40]&IN2[6];
  assign P47[17] = IN1[40]&IN2[7];
  assign P48[16] = IN1[40]&IN2[8];
  assign P49[15] = IN1[40]&IN2[9];
  assign P50[14] = IN1[40]&IN2[10];
  assign P51[13] = IN1[40]&IN2[11];
  assign P52[12] = IN1[40]&IN2[12];
  assign P53[11] = IN1[40]&IN2[13];
  assign P54[10] = IN1[40]&IN2[14];
  assign P55[9] = IN1[40]&IN2[15];
  assign P56[8] = IN1[40]&IN2[16];
  assign P57[7] = IN1[40]&IN2[17];
  assign P58[6] = IN1[40]&IN2[18];
  assign P59[5] = IN1[40]&IN2[19];
  assign P60[4] = IN1[40]&IN2[20];
  assign P61[3] = IN1[40]&IN2[21];
  assign P62[2] = IN1[40]&IN2[22];
  assign P63[1] = IN1[40]&IN2[23];
  assign P64[0] = IN1[40]&IN2[24];
  assign P41[24] = IN1[41]&IN2[0];
  assign P42[23] = IN1[41]&IN2[1];
  assign P43[22] = IN1[41]&IN2[2];
  assign P44[21] = IN1[41]&IN2[3];
  assign P45[20] = IN1[41]&IN2[4];
  assign P46[19] = IN1[41]&IN2[5];
  assign P47[18] = IN1[41]&IN2[6];
  assign P48[17] = IN1[41]&IN2[7];
  assign P49[16] = IN1[41]&IN2[8];
  assign P50[15] = IN1[41]&IN2[9];
  assign P51[14] = IN1[41]&IN2[10];
  assign P52[13] = IN1[41]&IN2[11];
  assign P53[12] = IN1[41]&IN2[12];
  assign P54[11] = IN1[41]&IN2[13];
  assign P55[10] = IN1[41]&IN2[14];
  assign P56[9] = IN1[41]&IN2[15];
  assign P57[8] = IN1[41]&IN2[16];
  assign P58[7] = IN1[41]&IN2[17];
  assign P59[6] = IN1[41]&IN2[18];
  assign P60[5] = IN1[41]&IN2[19];
  assign P61[4] = IN1[41]&IN2[20];
  assign P62[3] = IN1[41]&IN2[21];
  assign P63[2] = IN1[41]&IN2[22];
  assign P64[1] = IN1[41]&IN2[23];
  assign P65[0] = IN1[41]&IN2[24];
  assign P42[24] = IN1[42]&IN2[0];
  assign P43[23] = IN1[42]&IN2[1];
  assign P44[22] = IN1[42]&IN2[2];
  assign P45[21] = IN1[42]&IN2[3];
  assign P46[20] = IN1[42]&IN2[4];
  assign P47[19] = IN1[42]&IN2[5];
  assign P48[18] = IN1[42]&IN2[6];
  assign P49[17] = IN1[42]&IN2[7];
  assign P50[16] = IN1[42]&IN2[8];
  assign P51[15] = IN1[42]&IN2[9];
  assign P52[14] = IN1[42]&IN2[10];
  assign P53[13] = IN1[42]&IN2[11];
  assign P54[12] = IN1[42]&IN2[12];
  assign P55[11] = IN1[42]&IN2[13];
  assign P56[10] = IN1[42]&IN2[14];
  assign P57[9] = IN1[42]&IN2[15];
  assign P58[8] = IN1[42]&IN2[16];
  assign P59[7] = IN1[42]&IN2[17];
  assign P60[6] = IN1[42]&IN2[18];
  assign P61[5] = IN1[42]&IN2[19];
  assign P62[4] = IN1[42]&IN2[20];
  assign P63[3] = IN1[42]&IN2[21];
  assign P64[2] = IN1[42]&IN2[22];
  assign P65[1] = IN1[42]&IN2[23];
  assign P66[0] = IN1[42]&IN2[24];
  assign P43[24] = IN1[43]&IN2[0];
  assign P44[23] = IN1[43]&IN2[1];
  assign P45[22] = IN1[43]&IN2[2];
  assign P46[21] = IN1[43]&IN2[3];
  assign P47[20] = IN1[43]&IN2[4];
  assign P48[19] = IN1[43]&IN2[5];
  assign P49[18] = IN1[43]&IN2[6];
  assign P50[17] = IN1[43]&IN2[7];
  assign P51[16] = IN1[43]&IN2[8];
  assign P52[15] = IN1[43]&IN2[9];
  assign P53[14] = IN1[43]&IN2[10];
  assign P54[13] = IN1[43]&IN2[11];
  assign P55[12] = IN1[43]&IN2[12];
  assign P56[11] = IN1[43]&IN2[13];
  assign P57[10] = IN1[43]&IN2[14];
  assign P58[9] = IN1[43]&IN2[15];
  assign P59[8] = IN1[43]&IN2[16];
  assign P60[7] = IN1[43]&IN2[17];
  assign P61[6] = IN1[43]&IN2[18];
  assign P62[5] = IN1[43]&IN2[19];
  assign P63[4] = IN1[43]&IN2[20];
  assign P64[3] = IN1[43]&IN2[21];
  assign P65[2] = IN1[43]&IN2[22];
  assign P66[1] = IN1[43]&IN2[23];
  assign P67[0] = IN1[43]&IN2[24];
  assign P44[24] = IN1[44]&IN2[0];
  assign P45[23] = IN1[44]&IN2[1];
  assign P46[22] = IN1[44]&IN2[2];
  assign P47[21] = IN1[44]&IN2[3];
  assign P48[20] = IN1[44]&IN2[4];
  assign P49[19] = IN1[44]&IN2[5];
  assign P50[18] = IN1[44]&IN2[6];
  assign P51[17] = IN1[44]&IN2[7];
  assign P52[16] = IN1[44]&IN2[8];
  assign P53[15] = IN1[44]&IN2[9];
  assign P54[14] = IN1[44]&IN2[10];
  assign P55[13] = IN1[44]&IN2[11];
  assign P56[12] = IN1[44]&IN2[12];
  assign P57[11] = IN1[44]&IN2[13];
  assign P58[10] = IN1[44]&IN2[14];
  assign P59[9] = IN1[44]&IN2[15];
  assign P60[8] = IN1[44]&IN2[16];
  assign P61[7] = IN1[44]&IN2[17];
  assign P62[6] = IN1[44]&IN2[18];
  assign P63[5] = IN1[44]&IN2[19];
  assign P64[4] = IN1[44]&IN2[20];
  assign P65[3] = IN1[44]&IN2[21];
  assign P66[2] = IN1[44]&IN2[22];
  assign P67[1] = IN1[44]&IN2[23];
  assign P68[0] = IN1[44]&IN2[24];
  assign P45[24] = IN1[45]&IN2[0];
  assign P46[23] = IN1[45]&IN2[1];
  assign P47[22] = IN1[45]&IN2[2];
  assign P48[21] = IN1[45]&IN2[3];
  assign P49[20] = IN1[45]&IN2[4];
  assign P50[19] = IN1[45]&IN2[5];
  assign P51[18] = IN1[45]&IN2[6];
  assign P52[17] = IN1[45]&IN2[7];
  assign P53[16] = IN1[45]&IN2[8];
  assign P54[15] = IN1[45]&IN2[9];
  assign P55[14] = IN1[45]&IN2[10];
  assign P56[13] = IN1[45]&IN2[11];
  assign P57[12] = IN1[45]&IN2[12];
  assign P58[11] = IN1[45]&IN2[13];
  assign P59[10] = IN1[45]&IN2[14];
  assign P60[9] = IN1[45]&IN2[15];
  assign P61[8] = IN1[45]&IN2[16];
  assign P62[7] = IN1[45]&IN2[17];
  assign P63[6] = IN1[45]&IN2[18];
  assign P64[5] = IN1[45]&IN2[19];
  assign P65[4] = IN1[45]&IN2[20];
  assign P66[3] = IN1[45]&IN2[21];
  assign P67[2] = IN1[45]&IN2[22];
  assign P68[1] = IN1[45]&IN2[23];
  assign P69[0] = IN1[45]&IN2[24];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [24:0] IN25;
  input [24:0] IN26;
  input [24:0] IN27;
  input [24:0] IN28;
  input [24:0] IN29;
  input [24:0] IN30;
  input [24:0] IN31;
  input [24:0] IN32;
  input [24:0] IN33;
  input [24:0] IN34;
  input [24:0] IN35;
  input [24:0] IN36;
  input [24:0] IN37;
  input [24:0] IN38;
  input [24:0] IN39;
  input [24:0] IN40;
  input [24:0] IN41;
  input [24:0] IN42;
  input [24:0] IN43;
  input [24:0] IN44;
  input [24:0] IN45;
  input [23:0] IN46;
  input [22:0] IN47;
  input [21:0] IN48;
  input [20:0] IN49;
  input [19:0] IN50;
  input [18:0] IN51;
  input [17:0] IN52;
  input [16:0] IN53;
  input [15:0] IN54;
  input [14:0] IN55;
  input [13:0] IN56;
  input [12:0] IN57;
  input [11:0] IN58;
  input [10:0] IN59;
  input [9:0] IN60;
  input [8:0] IN61;
  input [7:0] IN62;
  input [6:0] IN63;
  input [5:0] IN64;
  input [4:0] IN65;
  input [3:0] IN66;
  input [2:0] IN67;
  input [1:0] IN68;
  input [0:0] IN69;
  output [69:0] Out1;
  output [23:0] Out2;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1984;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2088;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2585;
  wire w2586;
  wire w2587;
  wire w2588;
  wire w2589;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2614;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2631;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2638;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2685;
  wire w2686;
  wire w2687;
  wire w2688;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2694;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2708;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2738;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2747;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2774;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2785;
  wire w2786;
  wire w2787;
  wire w2788;
  wire w2789;
  wire w2790;
  wire w2791;
  wire w2792;
  wire w2793;
  wire w2794;
  wire w2795;
  wire w2796;
  wire w2797;
  wire w2798;
  wire w2799;
  wire w2800;
  wire w2801;
  wire w2802;
  wire w2803;
  wire w2804;
  wire w2805;
  wire w2806;
  wire w2807;
  wire w2808;
  wire w2809;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2854;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2861;
  wire w2862;
  wire w2863;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2885;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2896;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2913;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2934;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2979;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2985;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2990;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3014;
  wire w3015;
  wire w3016;
  wire w3017;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3084;
  wire w3085;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3094;
  wire w3095;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3121;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3221;
  wire w3223;
  wire w3225;
  wire w3227;
  wire w3229;
  wire w3231;
  wire w3233;
  wire w3235;
  wire w3237;
  wire w3239;
  wire w3241;
  wire w3243;
  wire w3245;
  wire w3247;
  wire w3249;
  wire w3251;
  wire w3253;
  wire w3255;
  wire w3257;
  wire w3259;
  wire w3261;
  wire w3263;
  wire w3265;
  wire w3267;
  wire w3269;
  wire w3271;
  wire w3273;
  wire w3275;
  wire w3277;
  wire w3279;
  wire w3281;
  wire w3283;
  wire w3285;
  wire w3287;
  wire w3289;
  wire w3291;
  wire w3293;
  wire w3295;
  wire w3297;
  wire w3299;
  wire w3301;
  wire w3303;
  wire w3305;
  wire w3307;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w1151);
  FullAdder U1 (w1151, IN2[0], IN2[1], w1152, w1153);
  FullAdder U2 (w1153, IN3[0], IN3[1], w1154, w1155);
  FullAdder U3 (w1155, IN4[0], IN4[1], w1156, w1157);
  FullAdder U4 (w1157, IN5[0], IN5[1], w1158, w1159);
  FullAdder U5 (w1159, IN6[0], IN6[1], w1160, w1161);
  FullAdder U6 (w1161, IN7[0], IN7[1], w1162, w1163);
  FullAdder U7 (w1163, IN8[0], IN8[1], w1164, w1165);
  FullAdder U8 (w1165, IN9[0], IN9[1], w1166, w1167);
  FullAdder U9 (w1167, IN10[0], IN10[1], w1168, w1169);
  FullAdder U10 (w1169, IN11[0], IN11[1], w1170, w1171);
  FullAdder U11 (w1171, IN12[0], IN12[1], w1172, w1173);
  FullAdder U12 (w1173, IN13[0], IN13[1], w1174, w1175);
  FullAdder U13 (w1175, IN14[0], IN14[1], w1176, w1177);
  FullAdder U14 (w1177, IN15[0], IN15[1], w1178, w1179);
  FullAdder U15 (w1179, IN16[0], IN16[1], w1180, w1181);
  FullAdder U16 (w1181, IN17[0], IN17[1], w1182, w1183);
  FullAdder U17 (w1183, IN18[0], IN18[1], w1184, w1185);
  FullAdder U18 (w1185, IN19[0], IN19[1], w1186, w1187);
  FullAdder U19 (w1187, IN20[0], IN20[1], w1188, w1189);
  FullAdder U20 (w1189, IN21[0], IN21[1], w1190, w1191);
  FullAdder U21 (w1191, IN22[0], IN22[1], w1192, w1193);
  FullAdder U22 (w1193, IN23[0], IN23[1], w1194, w1195);
  FullAdder U23 (w1195, IN24[0], IN24[1], w1196, w1197);
  FullAdder U24 (w1197, IN25[0], IN25[1], w1198, w1199);
  FullAdder U25 (w1199, IN26[0], IN26[1], w1200, w1201);
  FullAdder U26 (w1201, IN27[0], IN27[1], w1202, w1203);
  FullAdder U27 (w1203, IN28[0], IN28[1], w1204, w1205);
  FullAdder U28 (w1205, IN29[0], IN29[1], w1206, w1207);
  FullAdder U29 (w1207, IN30[0], IN30[1], w1208, w1209);
  FullAdder U30 (w1209, IN31[0], IN31[1], w1210, w1211);
  FullAdder U31 (w1211, IN32[0], IN32[1], w1212, w1213);
  FullAdder U32 (w1213, IN33[0], IN33[1], w1214, w1215);
  FullAdder U33 (w1215, IN34[0], IN34[1], w1216, w1217);
  FullAdder U34 (w1217, IN35[0], IN35[1], w1218, w1219);
  FullAdder U35 (w1219, IN36[0], IN36[1], w1220, w1221);
  FullAdder U36 (w1221, IN37[0], IN37[1], w1222, w1223);
  FullAdder U37 (w1223, IN38[0], IN38[1], w1224, w1225);
  FullAdder U38 (w1225, IN39[0], IN39[1], w1226, w1227);
  FullAdder U39 (w1227, IN40[0], IN40[1], w1228, w1229);
  FullAdder U40 (w1229, IN41[0], IN41[1], w1230, w1231);
  FullAdder U41 (w1231, IN42[0], IN42[1], w1232, w1233);
  FullAdder U42 (w1233, IN43[0], IN43[1], w1234, w1235);
  FullAdder U43 (w1235, IN44[0], IN44[1], w1236, w1237);
  FullAdder U44 (w1237, IN45[0], IN45[1], w1238, w1239);
  HalfAdder U45 (w1152, IN2[2], Out1[2], w1241);
  FullAdder U46 (w1241, w1154, IN3[2], w1242, w1243);
  FullAdder U47 (w1243, w1156, IN4[2], w1244, w1245);
  FullAdder U48 (w1245, w1158, IN5[2], w1246, w1247);
  FullAdder U49 (w1247, w1160, IN6[2], w1248, w1249);
  FullAdder U50 (w1249, w1162, IN7[2], w1250, w1251);
  FullAdder U51 (w1251, w1164, IN8[2], w1252, w1253);
  FullAdder U52 (w1253, w1166, IN9[2], w1254, w1255);
  FullAdder U53 (w1255, w1168, IN10[2], w1256, w1257);
  FullAdder U54 (w1257, w1170, IN11[2], w1258, w1259);
  FullAdder U55 (w1259, w1172, IN12[2], w1260, w1261);
  FullAdder U56 (w1261, w1174, IN13[2], w1262, w1263);
  FullAdder U57 (w1263, w1176, IN14[2], w1264, w1265);
  FullAdder U58 (w1265, w1178, IN15[2], w1266, w1267);
  FullAdder U59 (w1267, w1180, IN16[2], w1268, w1269);
  FullAdder U60 (w1269, w1182, IN17[2], w1270, w1271);
  FullAdder U61 (w1271, w1184, IN18[2], w1272, w1273);
  FullAdder U62 (w1273, w1186, IN19[2], w1274, w1275);
  FullAdder U63 (w1275, w1188, IN20[2], w1276, w1277);
  FullAdder U64 (w1277, w1190, IN21[2], w1278, w1279);
  FullAdder U65 (w1279, w1192, IN22[2], w1280, w1281);
  FullAdder U66 (w1281, w1194, IN23[2], w1282, w1283);
  FullAdder U67 (w1283, w1196, IN24[2], w1284, w1285);
  FullAdder U68 (w1285, w1198, IN25[2], w1286, w1287);
  FullAdder U69 (w1287, w1200, IN26[2], w1288, w1289);
  FullAdder U70 (w1289, w1202, IN27[2], w1290, w1291);
  FullAdder U71 (w1291, w1204, IN28[2], w1292, w1293);
  FullAdder U72 (w1293, w1206, IN29[2], w1294, w1295);
  FullAdder U73 (w1295, w1208, IN30[2], w1296, w1297);
  FullAdder U74 (w1297, w1210, IN31[2], w1298, w1299);
  FullAdder U75 (w1299, w1212, IN32[2], w1300, w1301);
  FullAdder U76 (w1301, w1214, IN33[2], w1302, w1303);
  FullAdder U77 (w1303, w1216, IN34[2], w1304, w1305);
  FullAdder U78 (w1305, w1218, IN35[2], w1306, w1307);
  FullAdder U79 (w1307, w1220, IN36[2], w1308, w1309);
  FullAdder U80 (w1309, w1222, IN37[2], w1310, w1311);
  FullAdder U81 (w1311, w1224, IN38[2], w1312, w1313);
  FullAdder U82 (w1313, w1226, IN39[2], w1314, w1315);
  FullAdder U83 (w1315, w1228, IN40[2], w1316, w1317);
  FullAdder U84 (w1317, w1230, IN41[2], w1318, w1319);
  FullAdder U85 (w1319, w1232, IN42[2], w1320, w1321);
  FullAdder U86 (w1321, w1234, IN43[2], w1322, w1323);
  FullAdder U87 (w1323, w1236, IN44[2], w1324, w1325);
  FullAdder U88 (w1325, w1238, IN45[2], w1326, w1327);
  FullAdder U89 (w1327, w1239, IN46[0], w1328, w1329);
  HalfAdder U90 (w1242, IN3[3], Out1[3], w1331);
  FullAdder U91 (w1331, w1244, IN4[3], w1332, w1333);
  FullAdder U92 (w1333, w1246, IN5[3], w1334, w1335);
  FullAdder U93 (w1335, w1248, IN6[3], w1336, w1337);
  FullAdder U94 (w1337, w1250, IN7[3], w1338, w1339);
  FullAdder U95 (w1339, w1252, IN8[3], w1340, w1341);
  FullAdder U96 (w1341, w1254, IN9[3], w1342, w1343);
  FullAdder U97 (w1343, w1256, IN10[3], w1344, w1345);
  FullAdder U98 (w1345, w1258, IN11[3], w1346, w1347);
  FullAdder U99 (w1347, w1260, IN12[3], w1348, w1349);
  FullAdder U100 (w1349, w1262, IN13[3], w1350, w1351);
  FullAdder U101 (w1351, w1264, IN14[3], w1352, w1353);
  FullAdder U102 (w1353, w1266, IN15[3], w1354, w1355);
  FullAdder U103 (w1355, w1268, IN16[3], w1356, w1357);
  FullAdder U104 (w1357, w1270, IN17[3], w1358, w1359);
  FullAdder U105 (w1359, w1272, IN18[3], w1360, w1361);
  FullAdder U106 (w1361, w1274, IN19[3], w1362, w1363);
  FullAdder U107 (w1363, w1276, IN20[3], w1364, w1365);
  FullAdder U108 (w1365, w1278, IN21[3], w1366, w1367);
  FullAdder U109 (w1367, w1280, IN22[3], w1368, w1369);
  FullAdder U110 (w1369, w1282, IN23[3], w1370, w1371);
  FullAdder U111 (w1371, w1284, IN24[3], w1372, w1373);
  FullAdder U112 (w1373, w1286, IN25[3], w1374, w1375);
  FullAdder U113 (w1375, w1288, IN26[3], w1376, w1377);
  FullAdder U114 (w1377, w1290, IN27[3], w1378, w1379);
  FullAdder U115 (w1379, w1292, IN28[3], w1380, w1381);
  FullAdder U116 (w1381, w1294, IN29[3], w1382, w1383);
  FullAdder U117 (w1383, w1296, IN30[3], w1384, w1385);
  FullAdder U118 (w1385, w1298, IN31[3], w1386, w1387);
  FullAdder U119 (w1387, w1300, IN32[3], w1388, w1389);
  FullAdder U120 (w1389, w1302, IN33[3], w1390, w1391);
  FullAdder U121 (w1391, w1304, IN34[3], w1392, w1393);
  FullAdder U122 (w1393, w1306, IN35[3], w1394, w1395);
  FullAdder U123 (w1395, w1308, IN36[3], w1396, w1397);
  FullAdder U124 (w1397, w1310, IN37[3], w1398, w1399);
  FullAdder U125 (w1399, w1312, IN38[3], w1400, w1401);
  FullAdder U126 (w1401, w1314, IN39[3], w1402, w1403);
  FullAdder U127 (w1403, w1316, IN40[3], w1404, w1405);
  FullAdder U128 (w1405, w1318, IN41[3], w1406, w1407);
  FullAdder U129 (w1407, w1320, IN42[3], w1408, w1409);
  FullAdder U130 (w1409, w1322, IN43[3], w1410, w1411);
  FullAdder U131 (w1411, w1324, IN44[3], w1412, w1413);
  FullAdder U132 (w1413, w1326, IN45[3], w1414, w1415);
  FullAdder U133 (w1415, w1328, IN46[1], w1416, w1417);
  FullAdder U134 (w1417, w1329, IN47[0], w1418, w1419);
  HalfAdder U135 (w1332, IN4[4], Out1[4], w1421);
  FullAdder U136 (w1421, w1334, IN5[4], w1422, w1423);
  FullAdder U137 (w1423, w1336, IN6[4], w1424, w1425);
  FullAdder U138 (w1425, w1338, IN7[4], w1426, w1427);
  FullAdder U139 (w1427, w1340, IN8[4], w1428, w1429);
  FullAdder U140 (w1429, w1342, IN9[4], w1430, w1431);
  FullAdder U141 (w1431, w1344, IN10[4], w1432, w1433);
  FullAdder U142 (w1433, w1346, IN11[4], w1434, w1435);
  FullAdder U143 (w1435, w1348, IN12[4], w1436, w1437);
  FullAdder U144 (w1437, w1350, IN13[4], w1438, w1439);
  FullAdder U145 (w1439, w1352, IN14[4], w1440, w1441);
  FullAdder U146 (w1441, w1354, IN15[4], w1442, w1443);
  FullAdder U147 (w1443, w1356, IN16[4], w1444, w1445);
  FullAdder U148 (w1445, w1358, IN17[4], w1446, w1447);
  FullAdder U149 (w1447, w1360, IN18[4], w1448, w1449);
  FullAdder U150 (w1449, w1362, IN19[4], w1450, w1451);
  FullAdder U151 (w1451, w1364, IN20[4], w1452, w1453);
  FullAdder U152 (w1453, w1366, IN21[4], w1454, w1455);
  FullAdder U153 (w1455, w1368, IN22[4], w1456, w1457);
  FullAdder U154 (w1457, w1370, IN23[4], w1458, w1459);
  FullAdder U155 (w1459, w1372, IN24[4], w1460, w1461);
  FullAdder U156 (w1461, w1374, IN25[4], w1462, w1463);
  FullAdder U157 (w1463, w1376, IN26[4], w1464, w1465);
  FullAdder U158 (w1465, w1378, IN27[4], w1466, w1467);
  FullAdder U159 (w1467, w1380, IN28[4], w1468, w1469);
  FullAdder U160 (w1469, w1382, IN29[4], w1470, w1471);
  FullAdder U161 (w1471, w1384, IN30[4], w1472, w1473);
  FullAdder U162 (w1473, w1386, IN31[4], w1474, w1475);
  FullAdder U163 (w1475, w1388, IN32[4], w1476, w1477);
  FullAdder U164 (w1477, w1390, IN33[4], w1478, w1479);
  FullAdder U165 (w1479, w1392, IN34[4], w1480, w1481);
  FullAdder U166 (w1481, w1394, IN35[4], w1482, w1483);
  FullAdder U167 (w1483, w1396, IN36[4], w1484, w1485);
  FullAdder U168 (w1485, w1398, IN37[4], w1486, w1487);
  FullAdder U169 (w1487, w1400, IN38[4], w1488, w1489);
  FullAdder U170 (w1489, w1402, IN39[4], w1490, w1491);
  FullAdder U171 (w1491, w1404, IN40[4], w1492, w1493);
  FullAdder U172 (w1493, w1406, IN41[4], w1494, w1495);
  FullAdder U173 (w1495, w1408, IN42[4], w1496, w1497);
  FullAdder U174 (w1497, w1410, IN43[4], w1498, w1499);
  FullAdder U175 (w1499, w1412, IN44[4], w1500, w1501);
  FullAdder U176 (w1501, w1414, IN45[4], w1502, w1503);
  FullAdder U177 (w1503, w1416, IN46[2], w1504, w1505);
  FullAdder U178 (w1505, w1418, IN47[1], w1506, w1507);
  FullAdder U179 (w1507, w1419, IN48[0], w1508, w1509);
  HalfAdder U180 (w1422, IN5[5], Out1[5], w1511);
  FullAdder U181 (w1511, w1424, IN6[5], w1512, w1513);
  FullAdder U182 (w1513, w1426, IN7[5], w1514, w1515);
  FullAdder U183 (w1515, w1428, IN8[5], w1516, w1517);
  FullAdder U184 (w1517, w1430, IN9[5], w1518, w1519);
  FullAdder U185 (w1519, w1432, IN10[5], w1520, w1521);
  FullAdder U186 (w1521, w1434, IN11[5], w1522, w1523);
  FullAdder U187 (w1523, w1436, IN12[5], w1524, w1525);
  FullAdder U188 (w1525, w1438, IN13[5], w1526, w1527);
  FullAdder U189 (w1527, w1440, IN14[5], w1528, w1529);
  FullAdder U190 (w1529, w1442, IN15[5], w1530, w1531);
  FullAdder U191 (w1531, w1444, IN16[5], w1532, w1533);
  FullAdder U192 (w1533, w1446, IN17[5], w1534, w1535);
  FullAdder U193 (w1535, w1448, IN18[5], w1536, w1537);
  FullAdder U194 (w1537, w1450, IN19[5], w1538, w1539);
  FullAdder U195 (w1539, w1452, IN20[5], w1540, w1541);
  FullAdder U196 (w1541, w1454, IN21[5], w1542, w1543);
  FullAdder U197 (w1543, w1456, IN22[5], w1544, w1545);
  FullAdder U198 (w1545, w1458, IN23[5], w1546, w1547);
  FullAdder U199 (w1547, w1460, IN24[5], w1548, w1549);
  FullAdder U200 (w1549, w1462, IN25[5], w1550, w1551);
  FullAdder U201 (w1551, w1464, IN26[5], w1552, w1553);
  FullAdder U202 (w1553, w1466, IN27[5], w1554, w1555);
  FullAdder U203 (w1555, w1468, IN28[5], w1556, w1557);
  FullAdder U204 (w1557, w1470, IN29[5], w1558, w1559);
  FullAdder U205 (w1559, w1472, IN30[5], w1560, w1561);
  FullAdder U206 (w1561, w1474, IN31[5], w1562, w1563);
  FullAdder U207 (w1563, w1476, IN32[5], w1564, w1565);
  FullAdder U208 (w1565, w1478, IN33[5], w1566, w1567);
  FullAdder U209 (w1567, w1480, IN34[5], w1568, w1569);
  FullAdder U210 (w1569, w1482, IN35[5], w1570, w1571);
  FullAdder U211 (w1571, w1484, IN36[5], w1572, w1573);
  FullAdder U212 (w1573, w1486, IN37[5], w1574, w1575);
  FullAdder U213 (w1575, w1488, IN38[5], w1576, w1577);
  FullAdder U214 (w1577, w1490, IN39[5], w1578, w1579);
  FullAdder U215 (w1579, w1492, IN40[5], w1580, w1581);
  FullAdder U216 (w1581, w1494, IN41[5], w1582, w1583);
  FullAdder U217 (w1583, w1496, IN42[5], w1584, w1585);
  FullAdder U218 (w1585, w1498, IN43[5], w1586, w1587);
  FullAdder U219 (w1587, w1500, IN44[5], w1588, w1589);
  FullAdder U220 (w1589, w1502, IN45[5], w1590, w1591);
  FullAdder U221 (w1591, w1504, IN46[3], w1592, w1593);
  FullAdder U222 (w1593, w1506, IN47[2], w1594, w1595);
  FullAdder U223 (w1595, w1508, IN48[1], w1596, w1597);
  FullAdder U224 (w1597, w1509, IN49[0], w1598, w1599);
  HalfAdder U225 (w1512, IN6[6], Out1[6], w1601);
  FullAdder U226 (w1601, w1514, IN7[6], w1602, w1603);
  FullAdder U227 (w1603, w1516, IN8[6], w1604, w1605);
  FullAdder U228 (w1605, w1518, IN9[6], w1606, w1607);
  FullAdder U229 (w1607, w1520, IN10[6], w1608, w1609);
  FullAdder U230 (w1609, w1522, IN11[6], w1610, w1611);
  FullAdder U231 (w1611, w1524, IN12[6], w1612, w1613);
  FullAdder U232 (w1613, w1526, IN13[6], w1614, w1615);
  FullAdder U233 (w1615, w1528, IN14[6], w1616, w1617);
  FullAdder U234 (w1617, w1530, IN15[6], w1618, w1619);
  FullAdder U235 (w1619, w1532, IN16[6], w1620, w1621);
  FullAdder U236 (w1621, w1534, IN17[6], w1622, w1623);
  FullAdder U237 (w1623, w1536, IN18[6], w1624, w1625);
  FullAdder U238 (w1625, w1538, IN19[6], w1626, w1627);
  FullAdder U239 (w1627, w1540, IN20[6], w1628, w1629);
  FullAdder U240 (w1629, w1542, IN21[6], w1630, w1631);
  FullAdder U241 (w1631, w1544, IN22[6], w1632, w1633);
  FullAdder U242 (w1633, w1546, IN23[6], w1634, w1635);
  FullAdder U243 (w1635, w1548, IN24[6], w1636, w1637);
  FullAdder U244 (w1637, w1550, IN25[6], w1638, w1639);
  FullAdder U245 (w1639, w1552, IN26[6], w1640, w1641);
  FullAdder U246 (w1641, w1554, IN27[6], w1642, w1643);
  FullAdder U247 (w1643, w1556, IN28[6], w1644, w1645);
  FullAdder U248 (w1645, w1558, IN29[6], w1646, w1647);
  FullAdder U249 (w1647, w1560, IN30[6], w1648, w1649);
  FullAdder U250 (w1649, w1562, IN31[6], w1650, w1651);
  FullAdder U251 (w1651, w1564, IN32[6], w1652, w1653);
  FullAdder U252 (w1653, w1566, IN33[6], w1654, w1655);
  FullAdder U253 (w1655, w1568, IN34[6], w1656, w1657);
  FullAdder U254 (w1657, w1570, IN35[6], w1658, w1659);
  FullAdder U255 (w1659, w1572, IN36[6], w1660, w1661);
  FullAdder U256 (w1661, w1574, IN37[6], w1662, w1663);
  FullAdder U257 (w1663, w1576, IN38[6], w1664, w1665);
  FullAdder U258 (w1665, w1578, IN39[6], w1666, w1667);
  FullAdder U259 (w1667, w1580, IN40[6], w1668, w1669);
  FullAdder U260 (w1669, w1582, IN41[6], w1670, w1671);
  FullAdder U261 (w1671, w1584, IN42[6], w1672, w1673);
  FullAdder U262 (w1673, w1586, IN43[6], w1674, w1675);
  FullAdder U263 (w1675, w1588, IN44[6], w1676, w1677);
  FullAdder U264 (w1677, w1590, IN45[6], w1678, w1679);
  FullAdder U265 (w1679, w1592, IN46[4], w1680, w1681);
  FullAdder U266 (w1681, w1594, IN47[3], w1682, w1683);
  FullAdder U267 (w1683, w1596, IN48[2], w1684, w1685);
  FullAdder U268 (w1685, w1598, IN49[1], w1686, w1687);
  FullAdder U269 (w1687, w1599, IN50[0], w1688, w1689);
  HalfAdder U270 (w1602, IN7[7], Out1[7], w1691);
  FullAdder U271 (w1691, w1604, IN8[7], w1692, w1693);
  FullAdder U272 (w1693, w1606, IN9[7], w1694, w1695);
  FullAdder U273 (w1695, w1608, IN10[7], w1696, w1697);
  FullAdder U274 (w1697, w1610, IN11[7], w1698, w1699);
  FullAdder U275 (w1699, w1612, IN12[7], w1700, w1701);
  FullAdder U276 (w1701, w1614, IN13[7], w1702, w1703);
  FullAdder U277 (w1703, w1616, IN14[7], w1704, w1705);
  FullAdder U278 (w1705, w1618, IN15[7], w1706, w1707);
  FullAdder U279 (w1707, w1620, IN16[7], w1708, w1709);
  FullAdder U280 (w1709, w1622, IN17[7], w1710, w1711);
  FullAdder U281 (w1711, w1624, IN18[7], w1712, w1713);
  FullAdder U282 (w1713, w1626, IN19[7], w1714, w1715);
  FullAdder U283 (w1715, w1628, IN20[7], w1716, w1717);
  FullAdder U284 (w1717, w1630, IN21[7], w1718, w1719);
  FullAdder U285 (w1719, w1632, IN22[7], w1720, w1721);
  FullAdder U286 (w1721, w1634, IN23[7], w1722, w1723);
  FullAdder U287 (w1723, w1636, IN24[7], w1724, w1725);
  FullAdder U288 (w1725, w1638, IN25[7], w1726, w1727);
  FullAdder U289 (w1727, w1640, IN26[7], w1728, w1729);
  FullAdder U290 (w1729, w1642, IN27[7], w1730, w1731);
  FullAdder U291 (w1731, w1644, IN28[7], w1732, w1733);
  FullAdder U292 (w1733, w1646, IN29[7], w1734, w1735);
  FullAdder U293 (w1735, w1648, IN30[7], w1736, w1737);
  FullAdder U294 (w1737, w1650, IN31[7], w1738, w1739);
  FullAdder U295 (w1739, w1652, IN32[7], w1740, w1741);
  FullAdder U296 (w1741, w1654, IN33[7], w1742, w1743);
  FullAdder U297 (w1743, w1656, IN34[7], w1744, w1745);
  FullAdder U298 (w1745, w1658, IN35[7], w1746, w1747);
  FullAdder U299 (w1747, w1660, IN36[7], w1748, w1749);
  FullAdder U300 (w1749, w1662, IN37[7], w1750, w1751);
  FullAdder U301 (w1751, w1664, IN38[7], w1752, w1753);
  FullAdder U302 (w1753, w1666, IN39[7], w1754, w1755);
  FullAdder U303 (w1755, w1668, IN40[7], w1756, w1757);
  FullAdder U304 (w1757, w1670, IN41[7], w1758, w1759);
  FullAdder U305 (w1759, w1672, IN42[7], w1760, w1761);
  FullAdder U306 (w1761, w1674, IN43[7], w1762, w1763);
  FullAdder U307 (w1763, w1676, IN44[7], w1764, w1765);
  FullAdder U308 (w1765, w1678, IN45[7], w1766, w1767);
  FullAdder U309 (w1767, w1680, IN46[5], w1768, w1769);
  FullAdder U310 (w1769, w1682, IN47[4], w1770, w1771);
  FullAdder U311 (w1771, w1684, IN48[3], w1772, w1773);
  FullAdder U312 (w1773, w1686, IN49[2], w1774, w1775);
  FullAdder U313 (w1775, w1688, IN50[1], w1776, w1777);
  FullAdder U314 (w1777, w1689, IN51[0], w1778, w1779);
  HalfAdder U315 (w1692, IN8[8], Out1[8], w1781);
  FullAdder U316 (w1781, w1694, IN9[8], w1782, w1783);
  FullAdder U317 (w1783, w1696, IN10[8], w1784, w1785);
  FullAdder U318 (w1785, w1698, IN11[8], w1786, w1787);
  FullAdder U319 (w1787, w1700, IN12[8], w1788, w1789);
  FullAdder U320 (w1789, w1702, IN13[8], w1790, w1791);
  FullAdder U321 (w1791, w1704, IN14[8], w1792, w1793);
  FullAdder U322 (w1793, w1706, IN15[8], w1794, w1795);
  FullAdder U323 (w1795, w1708, IN16[8], w1796, w1797);
  FullAdder U324 (w1797, w1710, IN17[8], w1798, w1799);
  FullAdder U325 (w1799, w1712, IN18[8], w1800, w1801);
  FullAdder U326 (w1801, w1714, IN19[8], w1802, w1803);
  FullAdder U327 (w1803, w1716, IN20[8], w1804, w1805);
  FullAdder U328 (w1805, w1718, IN21[8], w1806, w1807);
  FullAdder U329 (w1807, w1720, IN22[8], w1808, w1809);
  FullAdder U330 (w1809, w1722, IN23[8], w1810, w1811);
  FullAdder U331 (w1811, w1724, IN24[8], w1812, w1813);
  FullAdder U332 (w1813, w1726, IN25[8], w1814, w1815);
  FullAdder U333 (w1815, w1728, IN26[8], w1816, w1817);
  FullAdder U334 (w1817, w1730, IN27[8], w1818, w1819);
  FullAdder U335 (w1819, w1732, IN28[8], w1820, w1821);
  FullAdder U336 (w1821, w1734, IN29[8], w1822, w1823);
  FullAdder U337 (w1823, w1736, IN30[8], w1824, w1825);
  FullAdder U338 (w1825, w1738, IN31[8], w1826, w1827);
  FullAdder U339 (w1827, w1740, IN32[8], w1828, w1829);
  FullAdder U340 (w1829, w1742, IN33[8], w1830, w1831);
  FullAdder U341 (w1831, w1744, IN34[8], w1832, w1833);
  FullAdder U342 (w1833, w1746, IN35[8], w1834, w1835);
  FullAdder U343 (w1835, w1748, IN36[8], w1836, w1837);
  FullAdder U344 (w1837, w1750, IN37[8], w1838, w1839);
  FullAdder U345 (w1839, w1752, IN38[8], w1840, w1841);
  FullAdder U346 (w1841, w1754, IN39[8], w1842, w1843);
  FullAdder U347 (w1843, w1756, IN40[8], w1844, w1845);
  FullAdder U348 (w1845, w1758, IN41[8], w1846, w1847);
  FullAdder U349 (w1847, w1760, IN42[8], w1848, w1849);
  FullAdder U350 (w1849, w1762, IN43[8], w1850, w1851);
  FullAdder U351 (w1851, w1764, IN44[8], w1852, w1853);
  FullAdder U352 (w1853, w1766, IN45[8], w1854, w1855);
  FullAdder U353 (w1855, w1768, IN46[6], w1856, w1857);
  FullAdder U354 (w1857, w1770, IN47[5], w1858, w1859);
  FullAdder U355 (w1859, w1772, IN48[4], w1860, w1861);
  FullAdder U356 (w1861, w1774, IN49[3], w1862, w1863);
  FullAdder U357 (w1863, w1776, IN50[2], w1864, w1865);
  FullAdder U358 (w1865, w1778, IN51[1], w1866, w1867);
  FullAdder U359 (w1867, w1779, IN52[0], w1868, w1869);
  HalfAdder U360 (w1782, IN9[9], Out1[9], w1871);
  FullAdder U361 (w1871, w1784, IN10[9], w1872, w1873);
  FullAdder U362 (w1873, w1786, IN11[9], w1874, w1875);
  FullAdder U363 (w1875, w1788, IN12[9], w1876, w1877);
  FullAdder U364 (w1877, w1790, IN13[9], w1878, w1879);
  FullAdder U365 (w1879, w1792, IN14[9], w1880, w1881);
  FullAdder U366 (w1881, w1794, IN15[9], w1882, w1883);
  FullAdder U367 (w1883, w1796, IN16[9], w1884, w1885);
  FullAdder U368 (w1885, w1798, IN17[9], w1886, w1887);
  FullAdder U369 (w1887, w1800, IN18[9], w1888, w1889);
  FullAdder U370 (w1889, w1802, IN19[9], w1890, w1891);
  FullAdder U371 (w1891, w1804, IN20[9], w1892, w1893);
  FullAdder U372 (w1893, w1806, IN21[9], w1894, w1895);
  FullAdder U373 (w1895, w1808, IN22[9], w1896, w1897);
  FullAdder U374 (w1897, w1810, IN23[9], w1898, w1899);
  FullAdder U375 (w1899, w1812, IN24[9], w1900, w1901);
  FullAdder U376 (w1901, w1814, IN25[9], w1902, w1903);
  FullAdder U377 (w1903, w1816, IN26[9], w1904, w1905);
  FullAdder U378 (w1905, w1818, IN27[9], w1906, w1907);
  FullAdder U379 (w1907, w1820, IN28[9], w1908, w1909);
  FullAdder U380 (w1909, w1822, IN29[9], w1910, w1911);
  FullAdder U381 (w1911, w1824, IN30[9], w1912, w1913);
  FullAdder U382 (w1913, w1826, IN31[9], w1914, w1915);
  FullAdder U383 (w1915, w1828, IN32[9], w1916, w1917);
  FullAdder U384 (w1917, w1830, IN33[9], w1918, w1919);
  FullAdder U385 (w1919, w1832, IN34[9], w1920, w1921);
  FullAdder U386 (w1921, w1834, IN35[9], w1922, w1923);
  FullAdder U387 (w1923, w1836, IN36[9], w1924, w1925);
  FullAdder U388 (w1925, w1838, IN37[9], w1926, w1927);
  FullAdder U389 (w1927, w1840, IN38[9], w1928, w1929);
  FullAdder U390 (w1929, w1842, IN39[9], w1930, w1931);
  FullAdder U391 (w1931, w1844, IN40[9], w1932, w1933);
  FullAdder U392 (w1933, w1846, IN41[9], w1934, w1935);
  FullAdder U393 (w1935, w1848, IN42[9], w1936, w1937);
  FullAdder U394 (w1937, w1850, IN43[9], w1938, w1939);
  FullAdder U395 (w1939, w1852, IN44[9], w1940, w1941);
  FullAdder U396 (w1941, w1854, IN45[9], w1942, w1943);
  FullAdder U397 (w1943, w1856, IN46[7], w1944, w1945);
  FullAdder U398 (w1945, w1858, IN47[6], w1946, w1947);
  FullAdder U399 (w1947, w1860, IN48[5], w1948, w1949);
  FullAdder U400 (w1949, w1862, IN49[4], w1950, w1951);
  FullAdder U401 (w1951, w1864, IN50[3], w1952, w1953);
  FullAdder U402 (w1953, w1866, IN51[2], w1954, w1955);
  FullAdder U403 (w1955, w1868, IN52[1], w1956, w1957);
  FullAdder U404 (w1957, w1869, IN53[0], w1958, w1959);
  HalfAdder U405 (w1872, IN10[10], Out1[10], w1961);
  FullAdder U406 (w1961, w1874, IN11[10], w1962, w1963);
  FullAdder U407 (w1963, w1876, IN12[10], w1964, w1965);
  FullAdder U408 (w1965, w1878, IN13[10], w1966, w1967);
  FullAdder U409 (w1967, w1880, IN14[10], w1968, w1969);
  FullAdder U410 (w1969, w1882, IN15[10], w1970, w1971);
  FullAdder U411 (w1971, w1884, IN16[10], w1972, w1973);
  FullAdder U412 (w1973, w1886, IN17[10], w1974, w1975);
  FullAdder U413 (w1975, w1888, IN18[10], w1976, w1977);
  FullAdder U414 (w1977, w1890, IN19[10], w1978, w1979);
  FullAdder U415 (w1979, w1892, IN20[10], w1980, w1981);
  FullAdder U416 (w1981, w1894, IN21[10], w1982, w1983);
  FullAdder U417 (w1983, w1896, IN22[10], w1984, w1985);
  FullAdder U418 (w1985, w1898, IN23[10], w1986, w1987);
  FullAdder U419 (w1987, w1900, IN24[10], w1988, w1989);
  FullAdder U420 (w1989, w1902, IN25[10], w1990, w1991);
  FullAdder U421 (w1991, w1904, IN26[10], w1992, w1993);
  FullAdder U422 (w1993, w1906, IN27[10], w1994, w1995);
  FullAdder U423 (w1995, w1908, IN28[10], w1996, w1997);
  FullAdder U424 (w1997, w1910, IN29[10], w1998, w1999);
  FullAdder U425 (w1999, w1912, IN30[10], w2000, w2001);
  FullAdder U426 (w2001, w1914, IN31[10], w2002, w2003);
  FullAdder U427 (w2003, w1916, IN32[10], w2004, w2005);
  FullAdder U428 (w2005, w1918, IN33[10], w2006, w2007);
  FullAdder U429 (w2007, w1920, IN34[10], w2008, w2009);
  FullAdder U430 (w2009, w1922, IN35[10], w2010, w2011);
  FullAdder U431 (w2011, w1924, IN36[10], w2012, w2013);
  FullAdder U432 (w2013, w1926, IN37[10], w2014, w2015);
  FullAdder U433 (w2015, w1928, IN38[10], w2016, w2017);
  FullAdder U434 (w2017, w1930, IN39[10], w2018, w2019);
  FullAdder U435 (w2019, w1932, IN40[10], w2020, w2021);
  FullAdder U436 (w2021, w1934, IN41[10], w2022, w2023);
  FullAdder U437 (w2023, w1936, IN42[10], w2024, w2025);
  FullAdder U438 (w2025, w1938, IN43[10], w2026, w2027);
  FullAdder U439 (w2027, w1940, IN44[10], w2028, w2029);
  FullAdder U440 (w2029, w1942, IN45[10], w2030, w2031);
  FullAdder U441 (w2031, w1944, IN46[8], w2032, w2033);
  FullAdder U442 (w2033, w1946, IN47[7], w2034, w2035);
  FullAdder U443 (w2035, w1948, IN48[6], w2036, w2037);
  FullAdder U444 (w2037, w1950, IN49[5], w2038, w2039);
  FullAdder U445 (w2039, w1952, IN50[4], w2040, w2041);
  FullAdder U446 (w2041, w1954, IN51[3], w2042, w2043);
  FullAdder U447 (w2043, w1956, IN52[2], w2044, w2045);
  FullAdder U448 (w2045, w1958, IN53[1], w2046, w2047);
  FullAdder U449 (w2047, w1959, IN54[0], w2048, w2049);
  HalfAdder U450 (w1962, IN11[11], Out1[11], w2051);
  FullAdder U451 (w2051, w1964, IN12[11], w2052, w2053);
  FullAdder U452 (w2053, w1966, IN13[11], w2054, w2055);
  FullAdder U453 (w2055, w1968, IN14[11], w2056, w2057);
  FullAdder U454 (w2057, w1970, IN15[11], w2058, w2059);
  FullAdder U455 (w2059, w1972, IN16[11], w2060, w2061);
  FullAdder U456 (w2061, w1974, IN17[11], w2062, w2063);
  FullAdder U457 (w2063, w1976, IN18[11], w2064, w2065);
  FullAdder U458 (w2065, w1978, IN19[11], w2066, w2067);
  FullAdder U459 (w2067, w1980, IN20[11], w2068, w2069);
  FullAdder U460 (w2069, w1982, IN21[11], w2070, w2071);
  FullAdder U461 (w2071, w1984, IN22[11], w2072, w2073);
  FullAdder U462 (w2073, w1986, IN23[11], w2074, w2075);
  FullAdder U463 (w2075, w1988, IN24[11], w2076, w2077);
  FullAdder U464 (w2077, w1990, IN25[11], w2078, w2079);
  FullAdder U465 (w2079, w1992, IN26[11], w2080, w2081);
  FullAdder U466 (w2081, w1994, IN27[11], w2082, w2083);
  FullAdder U467 (w2083, w1996, IN28[11], w2084, w2085);
  FullAdder U468 (w2085, w1998, IN29[11], w2086, w2087);
  FullAdder U469 (w2087, w2000, IN30[11], w2088, w2089);
  FullAdder U470 (w2089, w2002, IN31[11], w2090, w2091);
  FullAdder U471 (w2091, w2004, IN32[11], w2092, w2093);
  FullAdder U472 (w2093, w2006, IN33[11], w2094, w2095);
  FullAdder U473 (w2095, w2008, IN34[11], w2096, w2097);
  FullAdder U474 (w2097, w2010, IN35[11], w2098, w2099);
  FullAdder U475 (w2099, w2012, IN36[11], w2100, w2101);
  FullAdder U476 (w2101, w2014, IN37[11], w2102, w2103);
  FullAdder U477 (w2103, w2016, IN38[11], w2104, w2105);
  FullAdder U478 (w2105, w2018, IN39[11], w2106, w2107);
  FullAdder U479 (w2107, w2020, IN40[11], w2108, w2109);
  FullAdder U480 (w2109, w2022, IN41[11], w2110, w2111);
  FullAdder U481 (w2111, w2024, IN42[11], w2112, w2113);
  FullAdder U482 (w2113, w2026, IN43[11], w2114, w2115);
  FullAdder U483 (w2115, w2028, IN44[11], w2116, w2117);
  FullAdder U484 (w2117, w2030, IN45[11], w2118, w2119);
  FullAdder U485 (w2119, w2032, IN46[9], w2120, w2121);
  FullAdder U486 (w2121, w2034, IN47[8], w2122, w2123);
  FullAdder U487 (w2123, w2036, IN48[7], w2124, w2125);
  FullAdder U488 (w2125, w2038, IN49[6], w2126, w2127);
  FullAdder U489 (w2127, w2040, IN50[5], w2128, w2129);
  FullAdder U490 (w2129, w2042, IN51[4], w2130, w2131);
  FullAdder U491 (w2131, w2044, IN52[3], w2132, w2133);
  FullAdder U492 (w2133, w2046, IN53[2], w2134, w2135);
  FullAdder U493 (w2135, w2048, IN54[1], w2136, w2137);
  FullAdder U494 (w2137, w2049, IN55[0], w2138, w2139);
  HalfAdder U495 (w2052, IN12[12], Out1[12], w2141);
  FullAdder U496 (w2141, w2054, IN13[12], w2142, w2143);
  FullAdder U497 (w2143, w2056, IN14[12], w2144, w2145);
  FullAdder U498 (w2145, w2058, IN15[12], w2146, w2147);
  FullAdder U499 (w2147, w2060, IN16[12], w2148, w2149);
  FullAdder U500 (w2149, w2062, IN17[12], w2150, w2151);
  FullAdder U501 (w2151, w2064, IN18[12], w2152, w2153);
  FullAdder U502 (w2153, w2066, IN19[12], w2154, w2155);
  FullAdder U503 (w2155, w2068, IN20[12], w2156, w2157);
  FullAdder U504 (w2157, w2070, IN21[12], w2158, w2159);
  FullAdder U505 (w2159, w2072, IN22[12], w2160, w2161);
  FullAdder U506 (w2161, w2074, IN23[12], w2162, w2163);
  FullAdder U507 (w2163, w2076, IN24[12], w2164, w2165);
  FullAdder U508 (w2165, w2078, IN25[12], w2166, w2167);
  FullAdder U509 (w2167, w2080, IN26[12], w2168, w2169);
  FullAdder U510 (w2169, w2082, IN27[12], w2170, w2171);
  FullAdder U511 (w2171, w2084, IN28[12], w2172, w2173);
  FullAdder U512 (w2173, w2086, IN29[12], w2174, w2175);
  FullAdder U513 (w2175, w2088, IN30[12], w2176, w2177);
  FullAdder U514 (w2177, w2090, IN31[12], w2178, w2179);
  FullAdder U515 (w2179, w2092, IN32[12], w2180, w2181);
  FullAdder U516 (w2181, w2094, IN33[12], w2182, w2183);
  FullAdder U517 (w2183, w2096, IN34[12], w2184, w2185);
  FullAdder U518 (w2185, w2098, IN35[12], w2186, w2187);
  FullAdder U519 (w2187, w2100, IN36[12], w2188, w2189);
  FullAdder U520 (w2189, w2102, IN37[12], w2190, w2191);
  FullAdder U521 (w2191, w2104, IN38[12], w2192, w2193);
  FullAdder U522 (w2193, w2106, IN39[12], w2194, w2195);
  FullAdder U523 (w2195, w2108, IN40[12], w2196, w2197);
  FullAdder U524 (w2197, w2110, IN41[12], w2198, w2199);
  FullAdder U525 (w2199, w2112, IN42[12], w2200, w2201);
  FullAdder U526 (w2201, w2114, IN43[12], w2202, w2203);
  FullAdder U527 (w2203, w2116, IN44[12], w2204, w2205);
  FullAdder U528 (w2205, w2118, IN45[12], w2206, w2207);
  FullAdder U529 (w2207, w2120, IN46[10], w2208, w2209);
  FullAdder U530 (w2209, w2122, IN47[9], w2210, w2211);
  FullAdder U531 (w2211, w2124, IN48[8], w2212, w2213);
  FullAdder U532 (w2213, w2126, IN49[7], w2214, w2215);
  FullAdder U533 (w2215, w2128, IN50[6], w2216, w2217);
  FullAdder U534 (w2217, w2130, IN51[5], w2218, w2219);
  FullAdder U535 (w2219, w2132, IN52[4], w2220, w2221);
  FullAdder U536 (w2221, w2134, IN53[3], w2222, w2223);
  FullAdder U537 (w2223, w2136, IN54[2], w2224, w2225);
  FullAdder U538 (w2225, w2138, IN55[1], w2226, w2227);
  FullAdder U539 (w2227, w2139, IN56[0], w2228, w2229);
  HalfAdder U540 (w2142, IN13[13], Out1[13], w2231);
  FullAdder U541 (w2231, w2144, IN14[13], w2232, w2233);
  FullAdder U542 (w2233, w2146, IN15[13], w2234, w2235);
  FullAdder U543 (w2235, w2148, IN16[13], w2236, w2237);
  FullAdder U544 (w2237, w2150, IN17[13], w2238, w2239);
  FullAdder U545 (w2239, w2152, IN18[13], w2240, w2241);
  FullAdder U546 (w2241, w2154, IN19[13], w2242, w2243);
  FullAdder U547 (w2243, w2156, IN20[13], w2244, w2245);
  FullAdder U548 (w2245, w2158, IN21[13], w2246, w2247);
  FullAdder U549 (w2247, w2160, IN22[13], w2248, w2249);
  FullAdder U550 (w2249, w2162, IN23[13], w2250, w2251);
  FullAdder U551 (w2251, w2164, IN24[13], w2252, w2253);
  FullAdder U552 (w2253, w2166, IN25[13], w2254, w2255);
  FullAdder U553 (w2255, w2168, IN26[13], w2256, w2257);
  FullAdder U554 (w2257, w2170, IN27[13], w2258, w2259);
  FullAdder U555 (w2259, w2172, IN28[13], w2260, w2261);
  FullAdder U556 (w2261, w2174, IN29[13], w2262, w2263);
  FullAdder U557 (w2263, w2176, IN30[13], w2264, w2265);
  FullAdder U558 (w2265, w2178, IN31[13], w2266, w2267);
  FullAdder U559 (w2267, w2180, IN32[13], w2268, w2269);
  FullAdder U560 (w2269, w2182, IN33[13], w2270, w2271);
  FullAdder U561 (w2271, w2184, IN34[13], w2272, w2273);
  FullAdder U562 (w2273, w2186, IN35[13], w2274, w2275);
  FullAdder U563 (w2275, w2188, IN36[13], w2276, w2277);
  FullAdder U564 (w2277, w2190, IN37[13], w2278, w2279);
  FullAdder U565 (w2279, w2192, IN38[13], w2280, w2281);
  FullAdder U566 (w2281, w2194, IN39[13], w2282, w2283);
  FullAdder U567 (w2283, w2196, IN40[13], w2284, w2285);
  FullAdder U568 (w2285, w2198, IN41[13], w2286, w2287);
  FullAdder U569 (w2287, w2200, IN42[13], w2288, w2289);
  FullAdder U570 (w2289, w2202, IN43[13], w2290, w2291);
  FullAdder U571 (w2291, w2204, IN44[13], w2292, w2293);
  FullAdder U572 (w2293, w2206, IN45[13], w2294, w2295);
  FullAdder U573 (w2295, w2208, IN46[11], w2296, w2297);
  FullAdder U574 (w2297, w2210, IN47[10], w2298, w2299);
  FullAdder U575 (w2299, w2212, IN48[9], w2300, w2301);
  FullAdder U576 (w2301, w2214, IN49[8], w2302, w2303);
  FullAdder U577 (w2303, w2216, IN50[7], w2304, w2305);
  FullAdder U578 (w2305, w2218, IN51[6], w2306, w2307);
  FullAdder U579 (w2307, w2220, IN52[5], w2308, w2309);
  FullAdder U580 (w2309, w2222, IN53[4], w2310, w2311);
  FullAdder U581 (w2311, w2224, IN54[3], w2312, w2313);
  FullAdder U582 (w2313, w2226, IN55[2], w2314, w2315);
  FullAdder U583 (w2315, w2228, IN56[1], w2316, w2317);
  FullAdder U584 (w2317, w2229, IN57[0], w2318, w2319);
  HalfAdder U585 (w2232, IN14[14], Out1[14], w2321);
  FullAdder U586 (w2321, w2234, IN15[14], w2322, w2323);
  FullAdder U587 (w2323, w2236, IN16[14], w2324, w2325);
  FullAdder U588 (w2325, w2238, IN17[14], w2326, w2327);
  FullAdder U589 (w2327, w2240, IN18[14], w2328, w2329);
  FullAdder U590 (w2329, w2242, IN19[14], w2330, w2331);
  FullAdder U591 (w2331, w2244, IN20[14], w2332, w2333);
  FullAdder U592 (w2333, w2246, IN21[14], w2334, w2335);
  FullAdder U593 (w2335, w2248, IN22[14], w2336, w2337);
  FullAdder U594 (w2337, w2250, IN23[14], w2338, w2339);
  FullAdder U595 (w2339, w2252, IN24[14], w2340, w2341);
  FullAdder U596 (w2341, w2254, IN25[14], w2342, w2343);
  FullAdder U597 (w2343, w2256, IN26[14], w2344, w2345);
  FullAdder U598 (w2345, w2258, IN27[14], w2346, w2347);
  FullAdder U599 (w2347, w2260, IN28[14], w2348, w2349);
  FullAdder U600 (w2349, w2262, IN29[14], w2350, w2351);
  FullAdder U601 (w2351, w2264, IN30[14], w2352, w2353);
  FullAdder U602 (w2353, w2266, IN31[14], w2354, w2355);
  FullAdder U603 (w2355, w2268, IN32[14], w2356, w2357);
  FullAdder U604 (w2357, w2270, IN33[14], w2358, w2359);
  FullAdder U605 (w2359, w2272, IN34[14], w2360, w2361);
  FullAdder U606 (w2361, w2274, IN35[14], w2362, w2363);
  FullAdder U607 (w2363, w2276, IN36[14], w2364, w2365);
  FullAdder U608 (w2365, w2278, IN37[14], w2366, w2367);
  FullAdder U609 (w2367, w2280, IN38[14], w2368, w2369);
  FullAdder U610 (w2369, w2282, IN39[14], w2370, w2371);
  FullAdder U611 (w2371, w2284, IN40[14], w2372, w2373);
  FullAdder U612 (w2373, w2286, IN41[14], w2374, w2375);
  FullAdder U613 (w2375, w2288, IN42[14], w2376, w2377);
  FullAdder U614 (w2377, w2290, IN43[14], w2378, w2379);
  FullAdder U615 (w2379, w2292, IN44[14], w2380, w2381);
  FullAdder U616 (w2381, w2294, IN45[14], w2382, w2383);
  FullAdder U617 (w2383, w2296, IN46[12], w2384, w2385);
  FullAdder U618 (w2385, w2298, IN47[11], w2386, w2387);
  FullAdder U619 (w2387, w2300, IN48[10], w2388, w2389);
  FullAdder U620 (w2389, w2302, IN49[9], w2390, w2391);
  FullAdder U621 (w2391, w2304, IN50[8], w2392, w2393);
  FullAdder U622 (w2393, w2306, IN51[7], w2394, w2395);
  FullAdder U623 (w2395, w2308, IN52[6], w2396, w2397);
  FullAdder U624 (w2397, w2310, IN53[5], w2398, w2399);
  FullAdder U625 (w2399, w2312, IN54[4], w2400, w2401);
  FullAdder U626 (w2401, w2314, IN55[3], w2402, w2403);
  FullAdder U627 (w2403, w2316, IN56[2], w2404, w2405);
  FullAdder U628 (w2405, w2318, IN57[1], w2406, w2407);
  FullAdder U629 (w2407, w2319, IN58[0], w2408, w2409);
  HalfAdder U630 (w2322, IN15[15], Out1[15], w2411);
  FullAdder U631 (w2411, w2324, IN16[15], w2412, w2413);
  FullAdder U632 (w2413, w2326, IN17[15], w2414, w2415);
  FullAdder U633 (w2415, w2328, IN18[15], w2416, w2417);
  FullAdder U634 (w2417, w2330, IN19[15], w2418, w2419);
  FullAdder U635 (w2419, w2332, IN20[15], w2420, w2421);
  FullAdder U636 (w2421, w2334, IN21[15], w2422, w2423);
  FullAdder U637 (w2423, w2336, IN22[15], w2424, w2425);
  FullAdder U638 (w2425, w2338, IN23[15], w2426, w2427);
  FullAdder U639 (w2427, w2340, IN24[15], w2428, w2429);
  FullAdder U640 (w2429, w2342, IN25[15], w2430, w2431);
  FullAdder U641 (w2431, w2344, IN26[15], w2432, w2433);
  FullAdder U642 (w2433, w2346, IN27[15], w2434, w2435);
  FullAdder U643 (w2435, w2348, IN28[15], w2436, w2437);
  FullAdder U644 (w2437, w2350, IN29[15], w2438, w2439);
  FullAdder U645 (w2439, w2352, IN30[15], w2440, w2441);
  FullAdder U646 (w2441, w2354, IN31[15], w2442, w2443);
  FullAdder U647 (w2443, w2356, IN32[15], w2444, w2445);
  FullAdder U648 (w2445, w2358, IN33[15], w2446, w2447);
  FullAdder U649 (w2447, w2360, IN34[15], w2448, w2449);
  FullAdder U650 (w2449, w2362, IN35[15], w2450, w2451);
  FullAdder U651 (w2451, w2364, IN36[15], w2452, w2453);
  FullAdder U652 (w2453, w2366, IN37[15], w2454, w2455);
  FullAdder U653 (w2455, w2368, IN38[15], w2456, w2457);
  FullAdder U654 (w2457, w2370, IN39[15], w2458, w2459);
  FullAdder U655 (w2459, w2372, IN40[15], w2460, w2461);
  FullAdder U656 (w2461, w2374, IN41[15], w2462, w2463);
  FullAdder U657 (w2463, w2376, IN42[15], w2464, w2465);
  FullAdder U658 (w2465, w2378, IN43[15], w2466, w2467);
  FullAdder U659 (w2467, w2380, IN44[15], w2468, w2469);
  FullAdder U660 (w2469, w2382, IN45[15], w2470, w2471);
  FullAdder U661 (w2471, w2384, IN46[13], w2472, w2473);
  FullAdder U662 (w2473, w2386, IN47[12], w2474, w2475);
  FullAdder U663 (w2475, w2388, IN48[11], w2476, w2477);
  FullAdder U664 (w2477, w2390, IN49[10], w2478, w2479);
  FullAdder U665 (w2479, w2392, IN50[9], w2480, w2481);
  FullAdder U666 (w2481, w2394, IN51[8], w2482, w2483);
  FullAdder U667 (w2483, w2396, IN52[7], w2484, w2485);
  FullAdder U668 (w2485, w2398, IN53[6], w2486, w2487);
  FullAdder U669 (w2487, w2400, IN54[5], w2488, w2489);
  FullAdder U670 (w2489, w2402, IN55[4], w2490, w2491);
  FullAdder U671 (w2491, w2404, IN56[3], w2492, w2493);
  FullAdder U672 (w2493, w2406, IN57[2], w2494, w2495);
  FullAdder U673 (w2495, w2408, IN58[1], w2496, w2497);
  FullAdder U674 (w2497, w2409, IN59[0], w2498, w2499);
  HalfAdder U675 (w2412, IN16[16], Out1[16], w2501);
  FullAdder U676 (w2501, w2414, IN17[16], w2502, w2503);
  FullAdder U677 (w2503, w2416, IN18[16], w2504, w2505);
  FullAdder U678 (w2505, w2418, IN19[16], w2506, w2507);
  FullAdder U679 (w2507, w2420, IN20[16], w2508, w2509);
  FullAdder U680 (w2509, w2422, IN21[16], w2510, w2511);
  FullAdder U681 (w2511, w2424, IN22[16], w2512, w2513);
  FullAdder U682 (w2513, w2426, IN23[16], w2514, w2515);
  FullAdder U683 (w2515, w2428, IN24[16], w2516, w2517);
  FullAdder U684 (w2517, w2430, IN25[16], w2518, w2519);
  FullAdder U685 (w2519, w2432, IN26[16], w2520, w2521);
  FullAdder U686 (w2521, w2434, IN27[16], w2522, w2523);
  FullAdder U687 (w2523, w2436, IN28[16], w2524, w2525);
  FullAdder U688 (w2525, w2438, IN29[16], w2526, w2527);
  FullAdder U689 (w2527, w2440, IN30[16], w2528, w2529);
  FullAdder U690 (w2529, w2442, IN31[16], w2530, w2531);
  FullAdder U691 (w2531, w2444, IN32[16], w2532, w2533);
  FullAdder U692 (w2533, w2446, IN33[16], w2534, w2535);
  FullAdder U693 (w2535, w2448, IN34[16], w2536, w2537);
  FullAdder U694 (w2537, w2450, IN35[16], w2538, w2539);
  FullAdder U695 (w2539, w2452, IN36[16], w2540, w2541);
  FullAdder U696 (w2541, w2454, IN37[16], w2542, w2543);
  FullAdder U697 (w2543, w2456, IN38[16], w2544, w2545);
  FullAdder U698 (w2545, w2458, IN39[16], w2546, w2547);
  FullAdder U699 (w2547, w2460, IN40[16], w2548, w2549);
  FullAdder U700 (w2549, w2462, IN41[16], w2550, w2551);
  FullAdder U701 (w2551, w2464, IN42[16], w2552, w2553);
  FullAdder U702 (w2553, w2466, IN43[16], w2554, w2555);
  FullAdder U703 (w2555, w2468, IN44[16], w2556, w2557);
  FullAdder U704 (w2557, w2470, IN45[16], w2558, w2559);
  FullAdder U705 (w2559, w2472, IN46[14], w2560, w2561);
  FullAdder U706 (w2561, w2474, IN47[13], w2562, w2563);
  FullAdder U707 (w2563, w2476, IN48[12], w2564, w2565);
  FullAdder U708 (w2565, w2478, IN49[11], w2566, w2567);
  FullAdder U709 (w2567, w2480, IN50[10], w2568, w2569);
  FullAdder U710 (w2569, w2482, IN51[9], w2570, w2571);
  FullAdder U711 (w2571, w2484, IN52[8], w2572, w2573);
  FullAdder U712 (w2573, w2486, IN53[7], w2574, w2575);
  FullAdder U713 (w2575, w2488, IN54[6], w2576, w2577);
  FullAdder U714 (w2577, w2490, IN55[5], w2578, w2579);
  FullAdder U715 (w2579, w2492, IN56[4], w2580, w2581);
  FullAdder U716 (w2581, w2494, IN57[3], w2582, w2583);
  FullAdder U717 (w2583, w2496, IN58[2], w2584, w2585);
  FullAdder U718 (w2585, w2498, IN59[1], w2586, w2587);
  FullAdder U719 (w2587, w2499, IN60[0], w2588, w2589);
  HalfAdder U720 (w2502, IN17[17], Out1[17], w2591);
  FullAdder U721 (w2591, w2504, IN18[17], w2592, w2593);
  FullAdder U722 (w2593, w2506, IN19[17], w2594, w2595);
  FullAdder U723 (w2595, w2508, IN20[17], w2596, w2597);
  FullAdder U724 (w2597, w2510, IN21[17], w2598, w2599);
  FullAdder U725 (w2599, w2512, IN22[17], w2600, w2601);
  FullAdder U726 (w2601, w2514, IN23[17], w2602, w2603);
  FullAdder U727 (w2603, w2516, IN24[17], w2604, w2605);
  FullAdder U728 (w2605, w2518, IN25[17], w2606, w2607);
  FullAdder U729 (w2607, w2520, IN26[17], w2608, w2609);
  FullAdder U730 (w2609, w2522, IN27[17], w2610, w2611);
  FullAdder U731 (w2611, w2524, IN28[17], w2612, w2613);
  FullAdder U732 (w2613, w2526, IN29[17], w2614, w2615);
  FullAdder U733 (w2615, w2528, IN30[17], w2616, w2617);
  FullAdder U734 (w2617, w2530, IN31[17], w2618, w2619);
  FullAdder U735 (w2619, w2532, IN32[17], w2620, w2621);
  FullAdder U736 (w2621, w2534, IN33[17], w2622, w2623);
  FullAdder U737 (w2623, w2536, IN34[17], w2624, w2625);
  FullAdder U738 (w2625, w2538, IN35[17], w2626, w2627);
  FullAdder U739 (w2627, w2540, IN36[17], w2628, w2629);
  FullAdder U740 (w2629, w2542, IN37[17], w2630, w2631);
  FullAdder U741 (w2631, w2544, IN38[17], w2632, w2633);
  FullAdder U742 (w2633, w2546, IN39[17], w2634, w2635);
  FullAdder U743 (w2635, w2548, IN40[17], w2636, w2637);
  FullAdder U744 (w2637, w2550, IN41[17], w2638, w2639);
  FullAdder U745 (w2639, w2552, IN42[17], w2640, w2641);
  FullAdder U746 (w2641, w2554, IN43[17], w2642, w2643);
  FullAdder U747 (w2643, w2556, IN44[17], w2644, w2645);
  FullAdder U748 (w2645, w2558, IN45[17], w2646, w2647);
  FullAdder U749 (w2647, w2560, IN46[15], w2648, w2649);
  FullAdder U750 (w2649, w2562, IN47[14], w2650, w2651);
  FullAdder U751 (w2651, w2564, IN48[13], w2652, w2653);
  FullAdder U752 (w2653, w2566, IN49[12], w2654, w2655);
  FullAdder U753 (w2655, w2568, IN50[11], w2656, w2657);
  FullAdder U754 (w2657, w2570, IN51[10], w2658, w2659);
  FullAdder U755 (w2659, w2572, IN52[9], w2660, w2661);
  FullAdder U756 (w2661, w2574, IN53[8], w2662, w2663);
  FullAdder U757 (w2663, w2576, IN54[7], w2664, w2665);
  FullAdder U758 (w2665, w2578, IN55[6], w2666, w2667);
  FullAdder U759 (w2667, w2580, IN56[5], w2668, w2669);
  FullAdder U760 (w2669, w2582, IN57[4], w2670, w2671);
  FullAdder U761 (w2671, w2584, IN58[3], w2672, w2673);
  FullAdder U762 (w2673, w2586, IN59[2], w2674, w2675);
  FullAdder U763 (w2675, w2588, IN60[1], w2676, w2677);
  FullAdder U764 (w2677, w2589, IN61[0], w2678, w2679);
  HalfAdder U765 (w2592, IN18[18], Out1[18], w2681);
  FullAdder U766 (w2681, w2594, IN19[18], w2682, w2683);
  FullAdder U767 (w2683, w2596, IN20[18], w2684, w2685);
  FullAdder U768 (w2685, w2598, IN21[18], w2686, w2687);
  FullAdder U769 (w2687, w2600, IN22[18], w2688, w2689);
  FullAdder U770 (w2689, w2602, IN23[18], w2690, w2691);
  FullAdder U771 (w2691, w2604, IN24[18], w2692, w2693);
  FullAdder U772 (w2693, w2606, IN25[18], w2694, w2695);
  FullAdder U773 (w2695, w2608, IN26[18], w2696, w2697);
  FullAdder U774 (w2697, w2610, IN27[18], w2698, w2699);
  FullAdder U775 (w2699, w2612, IN28[18], w2700, w2701);
  FullAdder U776 (w2701, w2614, IN29[18], w2702, w2703);
  FullAdder U777 (w2703, w2616, IN30[18], w2704, w2705);
  FullAdder U778 (w2705, w2618, IN31[18], w2706, w2707);
  FullAdder U779 (w2707, w2620, IN32[18], w2708, w2709);
  FullAdder U780 (w2709, w2622, IN33[18], w2710, w2711);
  FullAdder U781 (w2711, w2624, IN34[18], w2712, w2713);
  FullAdder U782 (w2713, w2626, IN35[18], w2714, w2715);
  FullAdder U783 (w2715, w2628, IN36[18], w2716, w2717);
  FullAdder U784 (w2717, w2630, IN37[18], w2718, w2719);
  FullAdder U785 (w2719, w2632, IN38[18], w2720, w2721);
  FullAdder U786 (w2721, w2634, IN39[18], w2722, w2723);
  FullAdder U787 (w2723, w2636, IN40[18], w2724, w2725);
  FullAdder U788 (w2725, w2638, IN41[18], w2726, w2727);
  FullAdder U789 (w2727, w2640, IN42[18], w2728, w2729);
  FullAdder U790 (w2729, w2642, IN43[18], w2730, w2731);
  FullAdder U791 (w2731, w2644, IN44[18], w2732, w2733);
  FullAdder U792 (w2733, w2646, IN45[18], w2734, w2735);
  FullAdder U793 (w2735, w2648, IN46[16], w2736, w2737);
  FullAdder U794 (w2737, w2650, IN47[15], w2738, w2739);
  FullAdder U795 (w2739, w2652, IN48[14], w2740, w2741);
  FullAdder U796 (w2741, w2654, IN49[13], w2742, w2743);
  FullAdder U797 (w2743, w2656, IN50[12], w2744, w2745);
  FullAdder U798 (w2745, w2658, IN51[11], w2746, w2747);
  FullAdder U799 (w2747, w2660, IN52[10], w2748, w2749);
  FullAdder U800 (w2749, w2662, IN53[9], w2750, w2751);
  FullAdder U801 (w2751, w2664, IN54[8], w2752, w2753);
  FullAdder U802 (w2753, w2666, IN55[7], w2754, w2755);
  FullAdder U803 (w2755, w2668, IN56[6], w2756, w2757);
  FullAdder U804 (w2757, w2670, IN57[5], w2758, w2759);
  FullAdder U805 (w2759, w2672, IN58[4], w2760, w2761);
  FullAdder U806 (w2761, w2674, IN59[3], w2762, w2763);
  FullAdder U807 (w2763, w2676, IN60[2], w2764, w2765);
  FullAdder U808 (w2765, w2678, IN61[1], w2766, w2767);
  FullAdder U809 (w2767, w2679, IN62[0], w2768, w2769);
  HalfAdder U810 (w2682, IN19[19], Out1[19], w2771);
  FullAdder U811 (w2771, w2684, IN20[19], w2772, w2773);
  FullAdder U812 (w2773, w2686, IN21[19], w2774, w2775);
  FullAdder U813 (w2775, w2688, IN22[19], w2776, w2777);
  FullAdder U814 (w2777, w2690, IN23[19], w2778, w2779);
  FullAdder U815 (w2779, w2692, IN24[19], w2780, w2781);
  FullAdder U816 (w2781, w2694, IN25[19], w2782, w2783);
  FullAdder U817 (w2783, w2696, IN26[19], w2784, w2785);
  FullAdder U818 (w2785, w2698, IN27[19], w2786, w2787);
  FullAdder U819 (w2787, w2700, IN28[19], w2788, w2789);
  FullAdder U820 (w2789, w2702, IN29[19], w2790, w2791);
  FullAdder U821 (w2791, w2704, IN30[19], w2792, w2793);
  FullAdder U822 (w2793, w2706, IN31[19], w2794, w2795);
  FullAdder U823 (w2795, w2708, IN32[19], w2796, w2797);
  FullAdder U824 (w2797, w2710, IN33[19], w2798, w2799);
  FullAdder U825 (w2799, w2712, IN34[19], w2800, w2801);
  FullAdder U826 (w2801, w2714, IN35[19], w2802, w2803);
  FullAdder U827 (w2803, w2716, IN36[19], w2804, w2805);
  FullAdder U828 (w2805, w2718, IN37[19], w2806, w2807);
  FullAdder U829 (w2807, w2720, IN38[19], w2808, w2809);
  FullAdder U830 (w2809, w2722, IN39[19], w2810, w2811);
  FullAdder U831 (w2811, w2724, IN40[19], w2812, w2813);
  FullAdder U832 (w2813, w2726, IN41[19], w2814, w2815);
  FullAdder U833 (w2815, w2728, IN42[19], w2816, w2817);
  FullAdder U834 (w2817, w2730, IN43[19], w2818, w2819);
  FullAdder U835 (w2819, w2732, IN44[19], w2820, w2821);
  FullAdder U836 (w2821, w2734, IN45[19], w2822, w2823);
  FullAdder U837 (w2823, w2736, IN46[17], w2824, w2825);
  FullAdder U838 (w2825, w2738, IN47[16], w2826, w2827);
  FullAdder U839 (w2827, w2740, IN48[15], w2828, w2829);
  FullAdder U840 (w2829, w2742, IN49[14], w2830, w2831);
  FullAdder U841 (w2831, w2744, IN50[13], w2832, w2833);
  FullAdder U842 (w2833, w2746, IN51[12], w2834, w2835);
  FullAdder U843 (w2835, w2748, IN52[11], w2836, w2837);
  FullAdder U844 (w2837, w2750, IN53[10], w2838, w2839);
  FullAdder U845 (w2839, w2752, IN54[9], w2840, w2841);
  FullAdder U846 (w2841, w2754, IN55[8], w2842, w2843);
  FullAdder U847 (w2843, w2756, IN56[7], w2844, w2845);
  FullAdder U848 (w2845, w2758, IN57[6], w2846, w2847);
  FullAdder U849 (w2847, w2760, IN58[5], w2848, w2849);
  FullAdder U850 (w2849, w2762, IN59[4], w2850, w2851);
  FullAdder U851 (w2851, w2764, IN60[3], w2852, w2853);
  FullAdder U852 (w2853, w2766, IN61[2], w2854, w2855);
  FullAdder U853 (w2855, w2768, IN62[1], w2856, w2857);
  FullAdder U854 (w2857, w2769, IN63[0], w2858, w2859);
  HalfAdder U855 (w2772, IN20[20], Out1[20], w2861);
  FullAdder U856 (w2861, w2774, IN21[20], w2862, w2863);
  FullAdder U857 (w2863, w2776, IN22[20], w2864, w2865);
  FullAdder U858 (w2865, w2778, IN23[20], w2866, w2867);
  FullAdder U859 (w2867, w2780, IN24[20], w2868, w2869);
  FullAdder U860 (w2869, w2782, IN25[20], w2870, w2871);
  FullAdder U861 (w2871, w2784, IN26[20], w2872, w2873);
  FullAdder U862 (w2873, w2786, IN27[20], w2874, w2875);
  FullAdder U863 (w2875, w2788, IN28[20], w2876, w2877);
  FullAdder U864 (w2877, w2790, IN29[20], w2878, w2879);
  FullAdder U865 (w2879, w2792, IN30[20], w2880, w2881);
  FullAdder U866 (w2881, w2794, IN31[20], w2882, w2883);
  FullAdder U867 (w2883, w2796, IN32[20], w2884, w2885);
  FullAdder U868 (w2885, w2798, IN33[20], w2886, w2887);
  FullAdder U869 (w2887, w2800, IN34[20], w2888, w2889);
  FullAdder U870 (w2889, w2802, IN35[20], w2890, w2891);
  FullAdder U871 (w2891, w2804, IN36[20], w2892, w2893);
  FullAdder U872 (w2893, w2806, IN37[20], w2894, w2895);
  FullAdder U873 (w2895, w2808, IN38[20], w2896, w2897);
  FullAdder U874 (w2897, w2810, IN39[20], w2898, w2899);
  FullAdder U875 (w2899, w2812, IN40[20], w2900, w2901);
  FullAdder U876 (w2901, w2814, IN41[20], w2902, w2903);
  FullAdder U877 (w2903, w2816, IN42[20], w2904, w2905);
  FullAdder U878 (w2905, w2818, IN43[20], w2906, w2907);
  FullAdder U879 (w2907, w2820, IN44[20], w2908, w2909);
  FullAdder U880 (w2909, w2822, IN45[20], w2910, w2911);
  FullAdder U881 (w2911, w2824, IN46[18], w2912, w2913);
  FullAdder U882 (w2913, w2826, IN47[17], w2914, w2915);
  FullAdder U883 (w2915, w2828, IN48[16], w2916, w2917);
  FullAdder U884 (w2917, w2830, IN49[15], w2918, w2919);
  FullAdder U885 (w2919, w2832, IN50[14], w2920, w2921);
  FullAdder U886 (w2921, w2834, IN51[13], w2922, w2923);
  FullAdder U887 (w2923, w2836, IN52[12], w2924, w2925);
  FullAdder U888 (w2925, w2838, IN53[11], w2926, w2927);
  FullAdder U889 (w2927, w2840, IN54[10], w2928, w2929);
  FullAdder U890 (w2929, w2842, IN55[9], w2930, w2931);
  FullAdder U891 (w2931, w2844, IN56[8], w2932, w2933);
  FullAdder U892 (w2933, w2846, IN57[7], w2934, w2935);
  FullAdder U893 (w2935, w2848, IN58[6], w2936, w2937);
  FullAdder U894 (w2937, w2850, IN59[5], w2938, w2939);
  FullAdder U895 (w2939, w2852, IN60[4], w2940, w2941);
  FullAdder U896 (w2941, w2854, IN61[3], w2942, w2943);
  FullAdder U897 (w2943, w2856, IN62[2], w2944, w2945);
  FullAdder U898 (w2945, w2858, IN63[1], w2946, w2947);
  FullAdder U899 (w2947, w2859, IN64[0], w2948, w2949);
  HalfAdder U900 (w2862, IN21[21], Out1[21], w2951);
  FullAdder U901 (w2951, w2864, IN22[21], w2952, w2953);
  FullAdder U902 (w2953, w2866, IN23[21], w2954, w2955);
  FullAdder U903 (w2955, w2868, IN24[21], w2956, w2957);
  FullAdder U904 (w2957, w2870, IN25[21], w2958, w2959);
  FullAdder U905 (w2959, w2872, IN26[21], w2960, w2961);
  FullAdder U906 (w2961, w2874, IN27[21], w2962, w2963);
  FullAdder U907 (w2963, w2876, IN28[21], w2964, w2965);
  FullAdder U908 (w2965, w2878, IN29[21], w2966, w2967);
  FullAdder U909 (w2967, w2880, IN30[21], w2968, w2969);
  FullAdder U910 (w2969, w2882, IN31[21], w2970, w2971);
  FullAdder U911 (w2971, w2884, IN32[21], w2972, w2973);
  FullAdder U912 (w2973, w2886, IN33[21], w2974, w2975);
  FullAdder U913 (w2975, w2888, IN34[21], w2976, w2977);
  FullAdder U914 (w2977, w2890, IN35[21], w2978, w2979);
  FullAdder U915 (w2979, w2892, IN36[21], w2980, w2981);
  FullAdder U916 (w2981, w2894, IN37[21], w2982, w2983);
  FullAdder U917 (w2983, w2896, IN38[21], w2984, w2985);
  FullAdder U918 (w2985, w2898, IN39[21], w2986, w2987);
  FullAdder U919 (w2987, w2900, IN40[21], w2988, w2989);
  FullAdder U920 (w2989, w2902, IN41[21], w2990, w2991);
  FullAdder U921 (w2991, w2904, IN42[21], w2992, w2993);
  FullAdder U922 (w2993, w2906, IN43[21], w2994, w2995);
  FullAdder U923 (w2995, w2908, IN44[21], w2996, w2997);
  FullAdder U924 (w2997, w2910, IN45[21], w2998, w2999);
  FullAdder U925 (w2999, w2912, IN46[19], w3000, w3001);
  FullAdder U926 (w3001, w2914, IN47[18], w3002, w3003);
  FullAdder U927 (w3003, w2916, IN48[17], w3004, w3005);
  FullAdder U928 (w3005, w2918, IN49[16], w3006, w3007);
  FullAdder U929 (w3007, w2920, IN50[15], w3008, w3009);
  FullAdder U930 (w3009, w2922, IN51[14], w3010, w3011);
  FullAdder U931 (w3011, w2924, IN52[13], w3012, w3013);
  FullAdder U932 (w3013, w2926, IN53[12], w3014, w3015);
  FullAdder U933 (w3015, w2928, IN54[11], w3016, w3017);
  FullAdder U934 (w3017, w2930, IN55[10], w3018, w3019);
  FullAdder U935 (w3019, w2932, IN56[9], w3020, w3021);
  FullAdder U936 (w3021, w2934, IN57[8], w3022, w3023);
  FullAdder U937 (w3023, w2936, IN58[7], w3024, w3025);
  FullAdder U938 (w3025, w2938, IN59[6], w3026, w3027);
  FullAdder U939 (w3027, w2940, IN60[5], w3028, w3029);
  FullAdder U940 (w3029, w2942, IN61[4], w3030, w3031);
  FullAdder U941 (w3031, w2944, IN62[3], w3032, w3033);
  FullAdder U942 (w3033, w2946, IN63[2], w3034, w3035);
  FullAdder U943 (w3035, w2948, IN64[1], w3036, w3037);
  FullAdder U944 (w3037, w2949, IN65[0], w3038, w3039);
  HalfAdder U945 (w2952, IN22[22], Out1[22], w3041);
  FullAdder U946 (w3041, w2954, IN23[22], w3042, w3043);
  FullAdder U947 (w3043, w2956, IN24[22], w3044, w3045);
  FullAdder U948 (w3045, w2958, IN25[22], w3046, w3047);
  FullAdder U949 (w3047, w2960, IN26[22], w3048, w3049);
  FullAdder U950 (w3049, w2962, IN27[22], w3050, w3051);
  FullAdder U951 (w3051, w2964, IN28[22], w3052, w3053);
  FullAdder U952 (w3053, w2966, IN29[22], w3054, w3055);
  FullAdder U953 (w3055, w2968, IN30[22], w3056, w3057);
  FullAdder U954 (w3057, w2970, IN31[22], w3058, w3059);
  FullAdder U955 (w3059, w2972, IN32[22], w3060, w3061);
  FullAdder U956 (w3061, w2974, IN33[22], w3062, w3063);
  FullAdder U957 (w3063, w2976, IN34[22], w3064, w3065);
  FullAdder U958 (w3065, w2978, IN35[22], w3066, w3067);
  FullAdder U959 (w3067, w2980, IN36[22], w3068, w3069);
  FullAdder U960 (w3069, w2982, IN37[22], w3070, w3071);
  FullAdder U961 (w3071, w2984, IN38[22], w3072, w3073);
  FullAdder U962 (w3073, w2986, IN39[22], w3074, w3075);
  FullAdder U963 (w3075, w2988, IN40[22], w3076, w3077);
  FullAdder U964 (w3077, w2990, IN41[22], w3078, w3079);
  FullAdder U965 (w3079, w2992, IN42[22], w3080, w3081);
  FullAdder U966 (w3081, w2994, IN43[22], w3082, w3083);
  FullAdder U967 (w3083, w2996, IN44[22], w3084, w3085);
  FullAdder U968 (w3085, w2998, IN45[22], w3086, w3087);
  FullAdder U969 (w3087, w3000, IN46[20], w3088, w3089);
  FullAdder U970 (w3089, w3002, IN47[19], w3090, w3091);
  FullAdder U971 (w3091, w3004, IN48[18], w3092, w3093);
  FullAdder U972 (w3093, w3006, IN49[17], w3094, w3095);
  FullAdder U973 (w3095, w3008, IN50[16], w3096, w3097);
  FullAdder U974 (w3097, w3010, IN51[15], w3098, w3099);
  FullAdder U975 (w3099, w3012, IN52[14], w3100, w3101);
  FullAdder U976 (w3101, w3014, IN53[13], w3102, w3103);
  FullAdder U977 (w3103, w3016, IN54[12], w3104, w3105);
  FullAdder U978 (w3105, w3018, IN55[11], w3106, w3107);
  FullAdder U979 (w3107, w3020, IN56[10], w3108, w3109);
  FullAdder U980 (w3109, w3022, IN57[9], w3110, w3111);
  FullAdder U981 (w3111, w3024, IN58[8], w3112, w3113);
  FullAdder U982 (w3113, w3026, IN59[7], w3114, w3115);
  FullAdder U983 (w3115, w3028, IN60[6], w3116, w3117);
  FullAdder U984 (w3117, w3030, IN61[5], w3118, w3119);
  FullAdder U985 (w3119, w3032, IN62[4], w3120, w3121);
  FullAdder U986 (w3121, w3034, IN63[3], w3122, w3123);
  FullAdder U987 (w3123, w3036, IN64[2], w3124, w3125);
  FullAdder U988 (w3125, w3038, IN65[1], w3126, w3127);
  FullAdder U989 (w3127, w3039, IN66[0], w3128, w3129);
  HalfAdder U990 (w3042, IN23[23], Out1[23], w3131);
  FullAdder U991 (w3131, w3044, IN24[23], w3132, w3133);
  FullAdder U992 (w3133, w3046, IN25[23], w3134, w3135);
  FullAdder U993 (w3135, w3048, IN26[23], w3136, w3137);
  FullAdder U994 (w3137, w3050, IN27[23], w3138, w3139);
  FullAdder U995 (w3139, w3052, IN28[23], w3140, w3141);
  FullAdder U996 (w3141, w3054, IN29[23], w3142, w3143);
  FullAdder U997 (w3143, w3056, IN30[23], w3144, w3145);
  FullAdder U998 (w3145, w3058, IN31[23], w3146, w3147);
  FullAdder U999 (w3147, w3060, IN32[23], w3148, w3149);
  FullAdder U1000 (w3149, w3062, IN33[23], w3150, w3151);
  FullAdder U1001 (w3151, w3064, IN34[23], w3152, w3153);
  FullAdder U1002 (w3153, w3066, IN35[23], w3154, w3155);
  FullAdder U1003 (w3155, w3068, IN36[23], w3156, w3157);
  FullAdder U1004 (w3157, w3070, IN37[23], w3158, w3159);
  FullAdder U1005 (w3159, w3072, IN38[23], w3160, w3161);
  FullAdder U1006 (w3161, w3074, IN39[23], w3162, w3163);
  FullAdder U1007 (w3163, w3076, IN40[23], w3164, w3165);
  FullAdder U1008 (w3165, w3078, IN41[23], w3166, w3167);
  FullAdder U1009 (w3167, w3080, IN42[23], w3168, w3169);
  FullAdder U1010 (w3169, w3082, IN43[23], w3170, w3171);
  FullAdder U1011 (w3171, w3084, IN44[23], w3172, w3173);
  FullAdder U1012 (w3173, w3086, IN45[23], w3174, w3175);
  FullAdder U1013 (w3175, w3088, IN46[21], w3176, w3177);
  FullAdder U1014 (w3177, w3090, IN47[20], w3178, w3179);
  FullAdder U1015 (w3179, w3092, IN48[19], w3180, w3181);
  FullAdder U1016 (w3181, w3094, IN49[18], w3182, w3183);
  FullAdder U1017 (w3183, w3096, IN50[17], w3184, w3185);
  FullAdder U1018 (w3185, w3098, IN51[16], w3186, w3187);
  FullAdder U1019 (w3187, w3100, IN52[15], w3188, w3189);
  FullAdder U1020 (w3189, w3102, IN53[14], w3190, w3191);
  FullAdder U1021 (w3191, w3104, IN54[13], w3192, w3193);
  FullAdder U1022 (w3193, w3106, IN55[12], w3194, w3195);
  FullAdder U1023 (w3195, w3108, IN56[11], w3196, w3197);
  FullAdder U1024 (w3197, w3110, IN57[10], w3198, w3199);
  FullAdder U1025 (w3199, w3112, IN58[9], w3200, w3201);
  FullAdder U1026 (w3201, w3114, IN59[8], w3202, w3203);
  FullAdder U1027 (w3203, w3116, IN60[7], w3204, w3205);
  FullAdder U1028 (w3205, w3118, IN61[6], w3206, w3207);
  FullAdder U1029 (w3207, w3120, IN62[5], w3208, w3209);
  FullAdder U1030 (w3209, w3122, IN63[4], w3210, w3211);
  FullAdder U1031 (w3211, w3124, IN64[3], w3212, w3213);
  FullAdder U1032 (w3213, w3126, IN65[2], w3214, w3215);
  FullAdder U1033 (w3215, w3128, IN66[1], w3216, w3217);
  FullAdder U1034 (w3217, w3129, IN67[0], w3218, w3219);
  HalfAdder U1035 (w3132, IN24[24], Out1[24], w3221);
  FullAdder U1036 (w3221, w3134, IN25[24], Out1[25], w3223);
  FullAdder U1037 (w3223, w3136, IN26[24], Out1[26], w3225);
  FullAdder U1038 (w3225, w3138, IN27[24], Out1[27], w3227);
  FullAdder U1039 (w3227, w3140, IN28[24], Out1[28], w3229);
  FullAdder U1040 (w3229, w3142, IN29[24], Out1[29], w3231);
  FullAdder U1041 (w3231, w3144, IN30[24], Out1[30], w3233);
  FullAdder U1042 (w3233, w3146, IN31[24], Out1[31], w3235);
  FullAdder U1043 (w3235, w3148, IN32[24], Out1[32], w3237);
  FullAdder U1044 (w3237, w3150, IN33[24], Out1[33], w3239);
  FullAdder U1045 (w3239, w3152, IN34[24], Out1[34], w3241);
  FullAdder U1046 (w3241, w3154, IN35[24], Out1[35], w3243);
  FullAdder U1047 (w3243, w3156, IN36[24], Out1[36], w3245);
  FullAdder U1048 (w3245, w3158, IN37[24], Out1[37], w3247);
  FullAdder U1049 (w3247, w3160, IN38[24], Out1[38], w3249);
  FullAdder U1050 (w3249, w3162, IN39[24], Out1[39], w3251);
  FullAdder U1051 (w3251, w3164, IN40[24], Out1[40], w3253);
  FullAdder U1052 (w3253, w3166, IN41[24], Out1[41], w3255);
  FullAdder U1053 (w3255, w3168, IN42[24], Out1[42], w3257);
  FullAdder U1054 (w3257, w3170, IN43[24], Out1[43], w3259);
  FullAdder U1055 (w3259, w3172, IN44[24], Out1[44], w3261);
  FullAdder U1056 (w3261, w3174, IN45[24], Out1[45], w3263);
  FullAdder U1057 (w3263, w3176, IN46[22], Out1[46], w3265);
  FullAdder U1058 (w3265, w3178, IN47[21], Out1[47], w3267);
  FullAdder U1059 (w3267, w3180, IN48[20], Out1[48], w3269);
  FullAdder U1060 (w3269, w3182, IN49[19], Out1[49], w3271);
  FullAdder U1061 (w3271, w3184, IN50[18], Out1[50], w3273);
  FullAdder U1062 (w3273, w3186, IN51[17], Out1[51], w3275);
  FullAdder U1063 (w3275, w3188, IN52[16], Out1[52], w3277);
  FullAdder U1064 (w3277, w3190, IN53[15], Out1[53], w3279);
  FullAdder U1065 (w3279, w3192, IN54[14], Out1[54], w3281);
  FullAdder U1066 (w3281, w3194, IN55[13], Out1[55], w3283);
  FullAdder U1067 (w3283, w3196, IN56[12], Out1[56], w3285);
  FullAdder U1068 (w3285, w3198, IN57[11], Out1[57], w3287);
  FullAdder U1069 (w3287, w3200, IN58[10], Out1[58], w3289);
  FullAdder U1070 (w3289, w3202, IN59[9], Out1[59], w3291);
  FullAdder U1071 (w3291, w3204, IN60[8], Out1[60], w3293);
  FullAdder U1072 (w3293, w3206, IN61[7], Out1[61], w3295);
  FullAdder U1073 (w3295, w3208, IN62[6], Out1[62], w3297);
  FullAdder U1074 (w3297, w3210, IN63[5], Out1[63], w3299);
  FullAdder U1075 (w3299, w3212, IN64[4], Out1[64], w3301);
  FullAdder U1076 (w3301, w3214, IN65[3], Out1[65], w3303);
  FullAdder U1077 (w3303, w3216, IN66[2], Out1[66], w3305);
  FullAdder U1078 (w3305, w3218, IN67[1], Out1[67], w3307);
  FullAdder U1079 (w3307, w3219, IN68[0], Out1[68], Out1[69]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN46[23];
  assign Out2[1] = IN47[22];
  assign Out2[2] = IN48[21];
  assign Out2[3] = IN49[20];
  assign Out2[4] = IN50[19];
  assign Out2[5] = IN51[18];
  assign Out2[6] = IN52[17];
  assign Out2[7] = IN53[16];
  assign Out2[8] = IN54[15];
  assign Out2[9] = IN55[14];
  assign Out2[10] = IN56[13];
  assign Out2[11] = IN57[12];
  assign Out2[12] = IN58[11];
  assign Out2[13] = IN59[10];
  assign Out2[14] = IN60[9];
  assign Out2[15] = IN61[8];
  assign Out2[16] = IN62[7];
  assign Out2[17] = IN63[6];
  assign Out2[18] = IN64[5];
  assign Out2[19] = IN65[4];
  assign Out2[20] = IN66[3];
  assign Out2[21] = IN67[2];
  assign Out2[22] = IN68[1];
  assign Out2[23] = IN69[0];

endmodule
module RC_24_24(IN1, IN2, Out);
  input [23:0] IN1;
  input [23:0] IN2;
  output [24:0] Out;
  wire w49;
  wire w51;
  wire w53;
  wire w55;
  wire w57;
  wire w59;
  wire w61;
  wire w63;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w49);
  FullAdder U1 (IN1[1], IN2[1], w49, Out[1], w51);
  FullAdder U2 (IN1[2], IN2[2], w51, Out[2], w53);
  FullAdder U3 (IN1[3], IN2[3], w53, Out[3], w55);
  FullAdder U4 (IN1[4], IN2[4], w55, Out[4], w57);
  FullAdder U5 (IN1[5], IN2[5], w57, Out[5], w59);
  FullAdder U6 (IN1[6], IN2[6], w59, Out[6], w61);
  FullAdder U7 (IN1[7], IN2[7], w61, Out[7], w63);
  FullAdder U8 (IN1[8], IN2[8], w63, Out[8], w65);
  FullAdder U9 (IN1[9], IN2[9], w65, Out[9], w67);
  FullAdder U10 (IN1[10], IN2[10], w67, Out[10], w69);
  FullAdder U11 (IN1[11], IN2[11], w69, Out[11], w71);
  FullAdder U12 (IN1[12], IN2[12], w71, Out[12], w73);
  FullAdder U13 (IN1[13], IN2[13], w73, Out[13], w75);
  FullAdder U14 (IN1[14], IN2[14], w75, Out[14], w77);
  FullAdder U15 (IN1[15], IN2[15], w77, Out[15], w79);
  FullAdder U16 (IN1[16], IN2[16], w79, Out[16], w81);
  FullAdder U17 (IN1[17], IN2[17], w81, Out[17], w83);
  FullAdder U18 (IN1[18], IN2[18], w83, Out[18], w85);
  FullAdder U19 (IN1[19], IN2[19], w85, Out[19], w87);
  FullAdder U20 (IN1[20], IN2[20], w87, Out[20], w89);
  FullAdder U21 (IN1[21], IN2[21], w89, Out[21], w91);
  FullAdder U22 (IN1[22], IN2[22], w91, Out[22], w93);
  FullAdder U23 (IN1[23], IN2[23], w93, Out[23], Out[24]);

endmodule
module NR_46_25(IN1, IN2, Out);
  input [45:0] IN1;
  input [24:0] IN2;
  output [70:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [24:0] P25;
  wire [24:0] P26;
  wire [24:0] P27;
  wire [24:0] P28;
  wire [24:0] P29;
  wire [24:0] P30;
  wire [24:0] P31;
  wire [24:0] P32;
  wire [24:0] P33;
  wire [24:0] P34;
  wire [24:0] P35;
  wire [24:0] P36;
  wire [24:0] P37;
  wire [24:0] P38;
  wire [24:0] P39;
  wire [24:0] P40;
  wire [24:0] P41;
  wire [24:0] P42;
  wire [24:0] P43;
  wire [24:0] P44;
  wire [24:0] P45;
  wire [23:0] P46;
  wire [22:0] P47;
  wire [21:0] P48;
  wire [20:0] P49;
  wire [19:0] P50;
  wire [18:0] P51;
  wire [17:0] P52;
  wire [16:0] P53;
  wire [15:0] P54;
  wire [14:0] P55;
  wire [13:0] P56;
  wire [12:0] P57;
  wire [11:0] P58;
  wire [10:0] P59;
  wire [9:0] P60;
  wire [8:0] P61;
  wire [7:0] P62;
  wire [6:0] P63;
  wire [5:0] P64;
  wire [4:0] P65;
  wire [3:0] P66;
  wire [2:0] P67;
  wire [1:0] P68;
  wire [0:0] P69;
  wire [69:0] R1;
  wire [23:0] R2;
  wire [70:0] aOut;
  U_SP_46_25 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, R1, R2);
  RC_24_24 S2 (R1[69:46], R2, aOut[70:46]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign Out = aOut[70:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
