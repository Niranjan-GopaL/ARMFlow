
module NR_1_62(
    input [0:0]IN1,
    input [61:0]IN2,
    output [61:0]Out
);
    assign Out = IN2;
endmodule
