
module NR_1_33(
    input [0:0]IN1,
    input [32:0]IN2,
    output [32:0]Out
);
    assign Out = IN2;
endmodule
