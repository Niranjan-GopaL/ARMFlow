//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 35
  second input length: 8
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_35_8(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41);
  input [34:0] IN1;
  input [7:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [7:0] P8;
  output [7:0] P9;
  output [7:0] P10;
  output [7:0] P11;
  output [7:0] P12;
  output [7:0] P13;
  output [7:0] P14;
  output [7:0] P15;
  output [7:0] P16;
  output [7:0] P17;
  output [7:0] P18;
  output [7:0] P19;
  output [7:0] P20;
  output [7:0] P21;
  output [7:0] P22;
  output [7:0] P23;
  output [7:0] P24;
  output [7:0] P25;
  output [7:0] P26;
  output [7:0] P27;
  output [7:0] P28;
  output [7:0] P29;
  output [7:0] P30;
  output [7:0] P31;
  output [7:0] P32;
  output [7:0] P33;
  output [7:0] P34;
  output [6:0] P35;
  output [5:0] P36;
  output [4:0] P37;
  output [3:0] P38;
  output [2:0] P39;
  output [1:0] P40;
  output [0:0] P41;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[0] = IN1[1]&IN2[7];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[1] = IN1[2]&IN2[6];
  assign P9[0] = IN1[2]&IN2[7];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[2] = IN1[3]&IN2[5];
  assign P9[1] = IN1[3]&IN2[6];
  assign P10[0] = IN1[3]&IN2[7];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[3] = IN1[4]&IN2[4];
  assign P9[2] = IN1[4]&IN2[5];
  assign P10[1] = IN1[4]&IN2[6];
  assign P11[0] = IN1[4]&IN2[7];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[4] = IN1[5]&IN2[3];
  assign P9[3] = IN1[5]&IN2[4];
  assign P10[2] = IN1[5]&IN2[5];
  assign P11[1] = IN1[5]&IN2[6];
  assign P12[0] = IN1[5]&IN2[7];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[5] = IN1[6]&IN2[2];
  assign P9[4] = IN1[6]&IN2[3];
  assign P10[3] = IN1[6]&IN2[4];
  assign P11[2] = IN1[6]&IN2[5];
  assign P12[1] = IN1[6]&IN2[6];
  assign P13[0] = IN1[6]&IN2[7];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[6] = IN1[7]&IN2[1];
  assign P9[5] = IN1[7]&IN2[2];
  assign P10[4] = IN1[7]&IN2[3];
  assign P11[3] = IN1[7]&IN2[4];
  assign P12[2] = IN1[7]&IN2[5];
  assign P13[1] = IN1[7]&IN2[6];
  assign P14[0] = IN1[7]&IN2[7];
  assign P8[7] = IN1[8]&IN2[0];
  assign P9[6] = IN1[8]&IN2[1];
  assign P10[5] = IN1[8]&IN2[2];
  assign P11[4] = IN1[8]&IN2[3];
  assign P12[3] = IN1[8]&IN2[4];
  assign P13[2] = IN1[8]&IN2[5];
  assign P14[1] = IN1[8]&IN2[6];
  assign P15[0] = IN1[8]&IN2[7];
  assign P9[7] = IN1[9]&IN2[0];
  assign P10[6] = IN1[9]&IN2[1];
  assign P11[5] = IN1[9]&IN2[2];
  assign P12[4] = IN1[9]&IN2[3];
  assign P13[3] = IN1[9]&IN2[4];
  assign P14[2] = IN1[9]&IN2[5];
  assign P15[1] = IN1[9]&IN2[6];
  assign P16[0] = IN1[9]&IN2[7];
  assign P10[7] = IN1[10]&IN2[0];
  assign P11[6] = IN1[10]&IN2[1];
  assign P12[5] = IN1[10]&IN2[2];
  assign P13[4] = IN1[10]&IN2[3];
  assign P14[3] = IN1[10]&IN2[4];
  assign P15[2] = IN1[10]&IN2[5];
  assign P16[1] = IN1[10]&IN2[6];
  assign P17[0] = IN1[10]&IN2[7];
  assign P11[7] = IN1[11]&IN2[0];
  assign P12[6] = IN1[11]&IN2[1];
  assign P13[5] = IN1[11]&IN2[2];
  assign P14[4] = IN1[11]&IN2[3];
  assign P15[3] = IN1[11]&IN2[4];
  assign P16[2] = IN1[11]&IN2[5];
  assign P17[1] = IN1[11]&IN2[6];
  assign P18[0] = IN1[11]&IN2[7];
  assign P12[7] = IN1[12]&IN2[0];
  assign P13[6] = IN1[12]&IN2[1];
  assign P14[5] = IN1[12]&IN2[2];
  assign P15[4] = IN1[12]&IN2[3];
  assign P16[3] = IN1[12]&IN2[4];
  assign P17[2] = IN1[12]&IN2[5];
  assign P18[1] = IN1[12]&IN2[6];
  assign P19[0] = IN1[12]&IN2[7];
  assign P13[7] = IN1[13]&IN2[0];
  assign P14[6] = IN1[13]&IN2[1];
  assign P15[5] = IN1[13]&IN2[2];
  assign P16[4] = IN1[13]&IN2[3];
  assign P17[3] = IN1[13]&IN2[4];
  assign P18[2] = IN1[13]&IN2[5];
  assign P19[1] = IN1[13]&IN2[6];
  assign P20[0] = IN1[13]&IN2[7];
  assign P14[7] = IN1[14]&IN2[0];
  assign P15[6] = IN1[14]&IN2[1];
  assign P16[5] = IN1[14]&IN2[2];
  assign P17[4] = IN1[14]&IN2[3];
  assign P18[3] = IN1[14]&IN2[4];
  assign P19[2] = IN1[14]&IN2[5];
  assign P20[1] = IN1[14]&IN2[6];
  assign P21[0] = IN1[14]&IN2[7];
  assign P15[7] = IN1[15]&IN2[0];
  assign P16[6] = IN1[15]&IN2[1];
  assign P17[5] = IN1[15]&IN2[2];
  assign P18[4] = IN1[15]&IN2[3];
  assign P19[3] = IN1[15]&IN2[4];
  assign P20[2] = IN1[15]&IN2[5];
  assign P21[1] = IN1[15]&IN2[6];
  assign P22[0] = IN1[15]&IN2[7];
  assign P16[7] = IN1[16]&IN2[0];
  assign P17[6] = IN1[16]&IN2[1];
  assign P18[5] = IN1[16]&IN2[2];
  assign P19[4] = IN1[16]&IN2[3];
  assign P20[3] = IN1[16]&IN2[4];
  assign P21[2] = IN1[16]&IN2[5];
  assign P22[1] = IN1[16]&IN2[6];
  assign P23[0] = IN1[16]&IN2[7];
  assign P17[7] = IN1[17]&IN2[0];
  assign P18[6] = IN1[17]&IN2[1];
  assign P19[5] = IN1[17]&IN2[2];
  assign P20[4] = IN1[17]&IN2[3];
  assign P21[3] = IN1[17]&IN2[4];
  assign P22[2] = IN1[17]&IN2[5];
  assign P23[1] = IN1[17]&IN2[6];
  assign P24[0] = IN1[17]&IN2[7];
  assign P18[7] = IN1[18]&IN2[0];
  assign P19[6] = IN1[18]&IN2[1];
  assign P20[5] = IN1[18]&IN2[2];
  assign P21[4] = IN1[18]&IN2[3];
  assign P22[3] = IN1[18]&IN2[4];
  assign P23[2] = IN1[18]&IN2[5];
  assign P24[1] = IN1[18]&IN2[6];
  assign P25[0] = IN1[18]&IN2[7];
  assign P19[7] = IN1[19]&IN2[0];
  assign P20[6] = IN1[19]&IN2[1];
  assign P21[5] = IN1[19]&IN2[2];
  assign P22[4] = IN1[19]&IN2[3];
  assign P23[3] = IN1[19]&IN2[4];
  assign P24[2] = IN1[19]&IN2[5];
  assign P25[1] = IN1[19]&IN2[6];
  assign P26[0] = IN1[19]&IN2[7];
  assign P20[7] = IN1[20]&IN2[0];
  assign P21[6] = IN1[20]&IN2[1];
  assign P22[5] = IN1[20]&IN2[2];
  assign P23[4] = IN1[20]&IN2[3];
  assign P24[3] = IN1[20]&IN2[4];
  assign P25[2] = IN1[20]&IN2[5];
  assign P26[1] = IN1[20]&IN2[6];
  assign P27[0] = IN1[20]&IN2[7];
  assign P21[7] = IN1[21]&IN2[0];
  assign P22[6] = IN1[21]&IN2[1];
  assign P23[5] = IN1[21]&IN2[2];
  assign P24[4] = IN1[21]&IN2[3];
  assign P25[3] = IN1[21]&IN2[4];
  assign P26[2] = IN1[21]&IN2[5];
  assign P27[1] = IN1[21]&IN2[6];
  assign P28[0] = IN1[21]&IN2[7];
  assign P22[7] = IN1[22]&IN2[0];
  assign P23[6] = IN1[22]&IN2[1];
  assign P24[5] = IN1[22]&IN2[2];
  assign P25[4] = IN1[22]&IN2[3];
  assign P26[3] = IN1[22]&IN2[4];
  assign P27[2] = IN1[22]&IN2[5];
  assign P28[1] = IN1[22]&IN2[6];
  assign P29[0] = IN1[22]&IN2[7];
  assign P23[7] = IN1[23]&IN2[0];
  assign P24[6] = IN1[23]&IN2[1];
  assign P25[5] = IN1[23]&IN2[2];
  assign P26[4] = IN1[23]&IN2[3];
  assign P27[3] = IN1[23]&IN2[4];
  assign P28[2] = IN1[23]&IN2[5];
  assign P29[1] = IN1[23]&IN2[6];
  assign P30[0] = IN1[23]&IN2[7];
  assign P24[7] = IN1[24]&IN2[0];
  assign P25[6] = IN1[24]&IN2[1];
  assign P26[5] = IN1[24]&IN2[2];
  assign P27[4] = IN1[24]&IN2[3];
  assign P28[3] = IN1[24]&IN2[4];
  assign P29[2] = IN1[24]&IN2[5];
  assign P30[1] = IN1[24]&IN2[6];
  assign P31[0] = IN1[24]&IN2[7];
  assign P25[7] = IN1[25]&IN2[0];
  assign P26[6] = IN1[25]&IN2[1];
  assign P27[5] = IN1[25]&IN2[2];
  assign P28[4] = IN1[25]&IN2[3];
  assign P29[3] = IN1[25]&IN2[4];
  assign P30[2] = IN1[25]&IN2[5];
  assign P31[1] = IN1[25]&IN2[6];
  assign P32[0] = IN1[25]&IN2[7];
  assign P26[7] = IN1[26]&IN2[0];
  assign P27[6] = IN1[26]&IN2[1];
  assign P28[5] = IN1[26]&IN2[2];
  assign P29[4] = IN1[26]&IN2[3];
  assign P30[3] = IN1[26]&IN2[4];
  assign P31[2] = IN1[26]&IN2[5];
  assign P32[1] = IN1[26]&IN2[6];
  assign P33[0] = IN1[26]&IN2[7];
  assign P27[7] = IN1[27]&IN2[0];
  assign P28[6] = IN1[27]&IN2[1];
  assign P29[5] = IN1[27]&IN2[2];
  assign P30[4] = IN1[27]&IN2[3];
  assign P31[3] = IN1[27]&IN2[4];
  assign P32[2] = IN1[27]&IN2[5];
  assign P33[1] = IN1[27]&IN2[6];
  assign P34[0] = IN1[27]&IN2[7];
  assign P28[7] = IN1[28]&IN2[0];
  assign P29[6] = IN1[28]&IN2[1];
  assign P30[5] = IN1[28]&IN2[2];
  assign P31[4] = IN1[28]&IN2[3];
  assign P32[3] = IN1[28]&IN2[4];
  assign P33[2] = IN1[28]&IN2[5];
  assign P34[1] = IN1[28]&IN2[6];
  assign P35[0] = IN1[28]&IN2[7];
  assign P29[7] = IN1[29]&IN2[0];
  assign P30[6] = IN1[29]&IN2[1];
  assign P31[5] = IN1[29]&IN2[2];
  assign P32[4] = IN1[29]&IN2[3];
  assign P33[3] = IN1[29]&IN2[4];
  assign P34[2] = IN1[29]&IN2[5];
  assign P35[1] = IN1[29]&IN2[6];
  assign P36[0] = IN1[29]&IN2[7];
  assign P30[7] = IN1[30]&IN2[0];
  assign P31[6] = IN1[30]&IN2[1];
  assign P32[5] = IN1[30]&IN2[2];
  assign P33[4] = IN1[30]&IN2[3];
  assign P34[3] = IN1[30]&IN2[4];
  assign P35[2] = IN1[30]&IN2[5];
  assign P36[1] = IN1[30]&IN2[6];
  assign P37[0] = IN1[30]&IN2[7];
  assign P31[7] = IN1[31]&IN2[0];
  assign P32[6] = IN1[31]&IN2[1];
  assign P33[5] = IN1[31]&IN2[2];
  assign P34[4] = IN1[31]&IN2[3];
  assign P35[3] = IN1[31]&IN2[4];
  assign P36[2] = IN1[31]&IN2[5];
  assign P37[1] = IN1[31]&IN2[6];
  assign P38[0] = IN1[31]&IN2[7];
  assign P32[7] = IN1[32]&IN2[0];
  assign P33[6] = IN1[32]&IN2[1];
  assign P34[5] = IN1[32]&IN2[2];
  assign P35[4] = IN1[32]&IN2[3];
  assign P36[3] = IN1[32]&IN2[4];
  assign P37[2] = IN1[32]&IN2[5];
  assign P38[1] = IN1[32]&IN2[6];
  assign P39[0] = IN1[32]&IN2[7];
  assign P33[7] = IN1[33]&IN2[0];
  assign P34[6] = IN1[33]&IN2[1];
  assign P35[5] = IN1[33]&IN2[2];
  assign P36[4] = IN1[33]&IN2[3];
  assign P37[3] = IN1[33]&IN2[4];
  assign P38[2] = IN1[33]&IN2[5];
  assign P39[1] = IN1[33]&IN2[6];
  assign P40[0] = IN1[33]&IN2[7];
  assign P34[7] = IN1[34]&IN2[0];
  assign P35[6] = IN1[34]&IN2[1];
  assign P36[5] = IN1[34]&IN2[2];
  assign P37[4] = IN1[34]&IN2[3];
  assign P38[3] = IN1[34]&IN2[4];
  assign P39[2] = IN1[34]&IN2[5];
  assign P40[1] = IN1[34]&IN2[6];
  assign P41[0] = IN1[34]&IN2[7];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [7:0] IN8;
  input [7:0] IN9;
  input [7:0] IN10;
  input [7:0] IN11;
  input [7:0] IN12;
  input [7:0] IN13;
  input [7:0] IN14;
  input [7:0] IN15;
  input [7:0] IN16;
  input [7:0] IN17;
  input [7:0] IN18;
  input [7:0] IN19;
  input [7:0] IN20;
  input [7:0] IN21;
  input [7:0] IN22;
  input [7:0] IN23;
  input [7:0] IN24;
  input [7:0] IN25;
  input [7:0] IN26;
  input [7:0] IN27;
  input [7:0] IN28;
  input [7:0] IN29;
  input [7:0] IN30;
  input [7:0] IN31;
  input [7:0] IN32;
  input [7:0] IN33;
  input [7:0] IN34;
  input [6:0] IN35;
  input [5:0] IN36;
  input [4:0] IN37;
  input [3:0] IN38;
  input [2:0] IN39;
  input [1:0] IN40;
  input [0:0] IN41;
  output [41:0] Out1;
  output [6:0] Out2;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w689;
  wire w691;
  wire w693;
  wire w695;
  wire w697;
  wire w699;
  wire w701;
  wire w703;
  wire w705;
  wire w707;
  wire w709;
  wire w711;
  wire w713;
  wire w715;
  wire w717;
  wire w719;
  wire w721;
  wire w723;
  wire w725;
  wire w727;
  wire w729;
  wire w731;
  wire w733;
  wire w735;
  wire w737;
  wire w739;
  wire w741;
  wire w743;
  wire w745;
  wire w747;
  wire w749;
  wire w751;
  wire w753;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w281);
  FullAdder U1 (w281, IN2[0], IN2[1], w282, w283);
  FullAdder U2 (w283, IN3[0], IN3[1], w284, w285);
  FullAdder U3 (w285, IN4[0], IN4[1], w286, w287);
  FullAdder U4 (w287, IN5[0], IN5[1], w288, w289);
  FullAdder U5 (w289, IN6[0], IN6[1], w290, w291);
  FullAdder U6 (w291, IN7[0], IN7[1], w292, w293);
  FullAdder U7 (w293, IN8[0], IN8[1], w294, w295);
  FullAdder U8 (w295, IN9[0], IN9[1], w296, w297);
  FullAdder U9 (w297, IN10[0], IN10[1], w298, w299);
  FullAdder U10 (w299, IN11[0], IN11[1], w300, w301);
  FullAdder U11 (w301, IN12[0], IN12[1], w302, w303);
  FullAdder U12 (w303, IN13[0], IN13[1], w304, w305);
  FullAdder U13 (w305, IN14[0], IN14[1], w306, w307);
  FullAdder U14 (w307, IN15[0], IN15[1], w308, w309);
  FullAdder U15 (w309, IN16[0], IN16[1], w310, w311);
  FullAdder U16 (w311, IN17[0], IN17[1], w312, w313);
  FullAdder U17 (w313, IN18[0], IN18[1], w314, w315);
  FullAdder U18 (w315, IN19[0], IN19[1], w316, w317);
  FullAdder U19 (w317, IN20[0], IN20[1], w318, w319);
  FullAdder U20 (w319, IN21[0], IN21[1], w320, w321);
  FullAdder U21 (w321, IN22[0], IN22[1], w322, w323);
  FullAdder U22 (w323, IN23[0], IN23[1], w324, w325);
  FullAdder U23 (w325, IN24[0], IN24[1], w326, w327);
  FullAdder U24 (w327, IN25[0], IN25[1], w328, w329);
  FullAdder U25 (w329, IN26[0], IN26[1], w330, w331);
  FullAdder U26 (w331, IN27[0], IN27[1], w332, w333);
  FullAdder U27 (w333, IN28[0], IN28[1], w334, w335);
  FullAdder U28 (w335, IN29[0], IN29[1], w336, w337);
  FullAdder U29 (w337, IN30[0], IN30[1], w338, w339);
  FullAdder U30 (w339, IN31[0], IN31[1], w340, w341);
  FullAdder U31 (w341, IN32[0], IN32[1], w342, w343);
  FullAdder U32 (w343, IN33[0], IN33[1], w344, w345);
  FullAdder U33 (w345, IN34[0], IN34[1], w346, w347);
  HalfAdder U34 (w282, IN2[2], Out1[2], w349);
  FullAdder U35 (w349, w284, IN3[2], w350, w351);
  FullAdder U36 (w351, w286, IN4[2], w352, w353);
  FullAdder U37 (w353, w288, IN5[2], w354, w355);
  FullAdder U38 (w355, w290, IN6[2], w356, w357);
  FullAdder U39 (w357, w292, IN7[2], w358, w359);
  FullAdder U40 (w359, w294, IN8[2], w360, w361);
  FullAdder U41 (w361, w296, IN9[2], w362, w363);
  FullAdder U42 (w363, w298, IN10[2], w364, w365);
  FullAdder U43 (w365, w300, IN11[2], w366, w367);
  FullAdder U44 (w367, w302, IN12[2], w368, w369);
  FullAdder U45 (w369, w304, IN13[2], w370, w371);
  FullAdder U46 (w371, w306, IN14[2], w372, w373);
  FullAdder U47 (w373, w308, IN15[2], w374, w375);
  FullAdder U48 (w375, w310, IN16[2], w376, w377);
  FullAdder U49 (w377, w312, IN17[2], w378, w379);
  FullAdder U50 (w379, w314, IN18[2], w380, w381);
  FullAdder U51 (w381, w316, IN19[2], w382, w383);
  FullAdder U52 (w383, w318, IN20[2], w384, w385);
  FullAdder U53 (w385, w320, IN21[2], w386, w387);
  FullAdder U54 (w387, w322, IN22[2], w388, w389);
  FullAdder U55 (w389, w324, IN23[2], w390, w391);
  FullAdder U56 (w391, w326, IN24[2], w392, w393);
  FullAdder U57 (w393, w328, IN25[2], w394, w395);
  FullAdder U58 (w395, w330, IN26[2], w396, w397);
  FullAdder U59 (w397, w332, IN27[2], w398, w399);
  FullAdder U60 (w399, w334, IN28[2], w400, w401);
  FullAdder U61 (w401, w336, IN29[2], w402, w403);
  FullAdder U62 (w403, w338, IN30[2], w404, w405);
  FullAdder U63 (w405, w340, IN31[2], w406, w407);
  FullAdder U64 (w407, w342, IN32[2], w408, w409);
  FullAdder U65 (w409, w344, IN33[2], w410, w411);
  FullAdder U66 (w411, w346, IN34[2], w412, w413);
  FullAdder U67 (w413, w347, IN35[0], w414, w415);
  HalfAdder U68 (w350, IN3[3], Out1[3], w417);
  FullAdder U69 (w417, w352, IN4[3], w418, w419);
  FullAdder U70 (w419, w354, IN5[3], w420, w421);
  FullAdder U71 (w421, w356, IN6[3], w422, w423);
  FullAdder U72 (w423, w358, IN7[3], w424, w425);
  FullAdder U73 (w425, w360, IN8[3], w426, w427);
  FullAdder U74 (w427, w362, IN9[3], w428, w429);
  FullAdder U75 (w429, w364, IN10[3], w430, w431);
  FullAdder U76 (w431, w366, IN11[3], w432, w433);
  FullAdder U77 (w433, w368, IN12[3], w434, w435);
  FullAdder U78 (w435, w370, IN13[3], w436, w437);
  FullAdder U79 (w437, w372, IN14[3], w438, w439);
  FullAdder U80 (w439, w374, IN15[3], w440, w441);
  FullAdder U81 (w441, w376, IN16[3], w442, w443);
  FullAdder U82 (w443, w378, IN17[3], w444, w445);
  FullAdder U83 (w445, w380, IN18[3], w446, w447);
  FullAdder U84 (w447, w382, IN19[3], w448, w449);
  FullAdder U85 (w449, w384, IN20[3], w450, w451);
  FullAdder U86 (w451, w386, IN21[3], w452, w453);
  FullAdder U87 (w453, w388, IN22[3], w454, w455);
  FullAdder U88 (w455, w390, IN23[3], w456, w457);
  FullAdder U89 (w457, w392, IN24[3], w458, w459);
  FullAdder U90 (w459, w394, IN25[3], w460, w461);
  FullAdder U91 (w461, w396, IN26[3], w462, w463);
  FullAdder U92 (w463, w398, IN27[3], w464, w465);
  FullAdder U93 (w465, w400, IN28[3], w466, w467);
  FullAdder U94 (w467, w402, IN29[3], w468, w469);
  FullAdder U95 (w469, w404, IN30[3], w470, w471);
  FullAdder U96 (w471, w406, IN31[3], w472, w473);
  FullAdder U97 (w473, w408, IN32[3], w474, w475);
  FullAdder U98 (w475, w410, IN33[3], w476, w477);
  FullAdder U99 (w477, w412, IN34[3], w478, w479);
  FullAdder U100 (w479, w414, IN35[1], w480, w481);
  FullAdder U101 (w481, w415, IN36[0], w482, w483);
  HalfAdder U102 (w418, IN4[4], Out1[4], w485);
  FullAdder U103 (w485, w420, IN5[4], w486, w487);
  FullAdder U104 (w487, w422, IN6[4], w488, w489);
  FullAdder U105 (w489, w424, IN7[4], w490, w491);
  FullAdder U106 (w491, w426, IN8[4], w492, w493);
  FullAdder U107 (w493, w428, IN9[4], w494, w495);
  FullAdder U108 (w495, w430, IN10[4], w496, w497);
  FullAdder U109 (w497, w432, IN11[4], w498, w499);
  FullAdder U110 (w499, w434, IN12[4], w500, w501);
  FullAdder U111 (w501, w436, IN13[4], w502, w503);
  FullAdder U112 (w503, w438, IN14[4], w504, w505);
  FullAdder U113 (w505, w440, IN15[4], w506, w507);
  FullAdder U114 (w507, w442, IN16[4], w508, w509);
  FullAdder U115 (w509, w444, IN17[4], w510, w511);
  FullAdder U116 (w511, w446, IN18[4], w512, w513);
  FullAdder U117 (w513, w448, IN19[4], w514, w515);
  FullAdder U118 (w515, w450, IN20[4], w516, w517);
  FullAdder U119 (w517, w452, IN21[4], w518, w519);
  FullAdder U120 (w519, w454, IN22[4], w520, w521);
  FullAdder U121 (w521, w456, IN23[4], w522, w523);
  FullAdder U122 (w523, w458, IN24[4], w524, w525);
  FullAdder U123 (w525, w460, IN25[4], w526, w527);
  FullAdder U124 (w527, w462, IN26[4], w528, w529);
  FullAdder U125 (w529, w464, IN27[4], w530, w531);
  FullAdder U126 (w531, w466, IN28[4], w532, w533);
  FullAdder U127 (w533, w468, IN29[4], w534, w535);
  FullAdder U128 (w535, w470, IN30[4], w536, w537);
  FullAdder U129 (w537, w472, IN31[4], w538, w539);
  FullAdder U130 (w539, w474, IN32[4], w540, w541);
  FullAdder U131 (w541, w476, IN33[4], w542, w543);
  FullAdder U132 (w543, w478, IN34[4], w544, w545);
  FullAdder U133 (w545, w480, IN35[2], w546, w547);
  FullAdder U134 (w547, w482, IN36[1], w548, w549);
  FullAdder U135 (w549, w483, IN37[0], w550, w551);
  HalfAdder U136 (w486, IN5[5], Out1[5], w553);
  FullAdder U137 (w553, w488, IN6[5], w554, w555);
  FullAdder U138 (w555, w490, IN7[5], w556, w557);
  FullAdder U139 (w557, w492, IN8[5], w558, w559);
  FullAdder U140 (w559, w494, IN9[5], w560, w561);
  FullAdder U141 (w561, w496, IN10[5], w562, w563);
  FullAdder U142 (w563, w498, IN11[5], w564, w565);
  FullAdder U143 (w565, w500, IN12[5], w566, w567);
  FullAdder U144 (w567, w502, IN13[5], w568, w569);
  FullAdder U145 (w569, w504, IN14[5], w570, w571);
  FullAdder U146 (w571, w506, IN15[5], w572, w573);
  FullAdder U147 (w573, w508, IN16[5], w574, w575);
  FullAdder U148 (w575, w510, IN17[5], w576, w577);
  FullAdder U149 (w577, w512, IN18[5], w578, w579);
  FullAdder U150 (w579, w514, IN19[5], w580, w581);
  FullAdder U151 (w581, w516, IN20[5], w582, w583);
  FullAdder U152 (w583, w518, IN21[5], w584, w585);
  FullAdder U153 (w585, w520, IN22[5], w586, w587);
  FullAdder U154 (w587, w522, IN23[5], w588, w589);
  FullAdder U155 (w589, w524, IN24[5], w590, w591);
  FullAdder U156 (w591, w526, IN25[5], w592, w593);
  FullAdder U157 (w593, w528, IN26[5], w594, w595);
  FullAdder U158 (w595, w530, IN27[5], w596, w597);
  FullAdder U159 (w597, w532, IN28[5], w598, w599);
  FullAdder U160 (w599, w534, IN29[5], w600, w601);
  FullAdder U161 (w601, w536, IN30[5], w602, w603);
  FullAdder U162 (w603, w538, IN31[5], w604, w605);
  FullAdder U163 (w605, w540, IN32[5], w606, w607);
  FullAdder U164 (w607, w542, IN33[5], w608, w609);
  FullAdder U165 (w609, w544, IN34[5], w610, w611);
  FullAdder U166 (w611, w546, IN35[3], w612, w613);
  FullAdder U167 (w613, w548, IN36[2], w614, w615);
  FullAdder U168 (w615, w550, IN37[1], w616, w617);
  FullAdder U169 (w617, w551, IN38[0], w618, w619);
  HalfAdder U170 (w554, IN6[6], Out1[6], w621);
  FullAdder U171 (w621, w556, IN7[6], w622, w623);
  FullAdder U172 (w623, w558, IN8[6], w624, w625);
  FullAdder U173 (w625, w560, IN9[6], w626, w627);
  FullAdder U174 (w627, w562, IN10[6], w628, w629);
  FullAdder U175 (w629, w564, IN11[6], w630, w631);
  FullAdder U176 (w631, w566, IN12[6], w632, w633);
  FullAdder U177 (w633, w568, IN13[6], w634, w635);
  FullAdder U178 (w635, w570, IN14[6], w636, w637);
  FullAdder U179 (w637, w572, IN15[6], w638, w639);
  FullAdder U180 (w639, w574, IN16[6], w640, w641);
  FullAdder U181 (w641, w576, IN17[6], w642, w643);
  FullAdder U182 (w643, w578, IN18[6], w644, w645);
  FullAdder U183 (w645, w580, IN19[6], w646, w647);
  FullAdder U184 (w647, w582, IN20[6], w648, w649);
  FullAdder U185 (w649, w584, IN21[6], w650, w651);
  FullAdder U186 (w651, w586, IN22[6], w652, w653);
  FullAdder U187 (w653, w588, IN23[6], w654, w655);
  FullAdder U188 (w655, w590, IN24[6], w656, w657);
  FullAdder U189 (w657, w592, IN25[6], w658, w659);
  FullAdder U190 (w659, w594, IN26[6], w660, w661);
  FullAdder U191 (w661, w596, IN27[6], w662, w663);
  FullAdder U192 (w663, w598, IN28[6], w664, w665);
  FullAdder U193 (w665, w600, IN29[6], w666, w667);
  FullAdder U194 (w667, w602, IN30[6], w668, w669);
  FullAdder U195 (w669, w604, IN31[6], w670, w671);
  FullAdder U196 (w671, w606, IN32[6], w672, w673);
  FullAdder U197 (w673, w608, IN33[6], w674, w675);
  FullAdder U198 (w675, w610, IN34[6], w676, w677);
  FullAdder U199 (w677, w612, IN35[4], w678, w679);
  FullAdder U200 (w679, w614, IN36[3], w680, w681);
  FullAdder U201 (w681, w616, IN37[2], w682, w683);
  FullAdder U202 (w683, w618, IN38[1], w684, w685);
  FullAdder U203 (w685, w619, IN39[0], w686, w687);
  HalfAdder U204 (w622, IN7[7], Out1[7], w689);
  FullAdder U205 (w689, w624, IN8[7], Out1[8], w691);
  FullAdder U206 (w691, w626, IN9[7], Out1[9], w693);
  FullAdder U207 (w693, w628, IN10[7], Out1[10], w695);
  FullAdder U208 (w695, w630, IN11[7], Out1[11], w697);
  FullAdder U209 (w697, w632, IN12[7], Out1[12], w699);
  FullAdder U210 (w699, w634, IN13[7], Out1[13], w701);
  FullAdder U211 (w701, w636, IN14[7], Out1[14], w703);
  FullAdder U212 (w703, w638, IN15[7], Out1[15], w705);
  FullAdder U213 (w705, w640, IN16[7], Out1[16], w707);
  FullAdder U214 (w707, w642, IN17[7], Out1[17], w709);
  FullAdder U215 (w709, w644, IN18[7], Out1[18], w711);
  FullAdder U216 (w711, w646, IN19[7], Out1[19], w713);
  FullAdder U217 (w713, w648, IN20[7], Out1[20], w715);
  FullAdder U218 (w715, w650, IN21[7], Out1[21], w717);
  FullAdder U219 (w717, w652, IN22[7], Out1[22], w719);
  FullAdder U220 (w719, w654, IN23[7], Out1[23], w721);
  FullAdder U221 (w721, w656, IN24[7], Out1[24], w723);
  FullAdder U222 (w723, w658, IN25[7], Out1[25], w725);
  FullAdder U223 (w725, w660, IN26[7], Out1[26], w727);
  FullAdder U224 (w727, w662, IN27[7], Out1[27], w729);
  FullAdder U225 (w729, w664, IN28[7], Out1[28], w731);
  FullAdder U226 (w731, w666, IN29[7], Out1[29], w733);
  FullAdder U227 (w733, w668, IN30[7], Out1[30], w735);
  FullAdder U228 (w735, w670, IN31[7], Out1[31], w737);
  FullAdder U229 (w737, w672, IN32[7], Out1[32], w739);
  FullAdder U230 (w739, w674, IN33[7], Out1[33], w741);
  FullAdder U231 (w741, w676, IN34[7], Out1[34], w743);
  FullAdder U232 (w743, w678, IN35[5], Out1[35], w745);
  FullAdder U233 (w745, w680, IN36[4], Out1[36], w747);
  FullAdder U234 (w747, w682, IN37[3], Out1[37], w749);
  FullAdder U235 (w749, w684, IN38[2], Out1[38], w751);
  FullAdder U236 (w751, w686, IN39[1], Out1[39], w753);
  FullAdder U237 (w753, w687, IN40[0], Out1[40], Out1[41]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN35[6];
  assign Out2[1] = IN36[5];
  assign Out2[2] = IN37[4];
  assign Out2[3] = IN38[3];
  assign Out2[4] = IN39[2];
  assign Out2[5] = IN40[1];
  assign Out2[6] = IN41[0];

endmodule
module RC_7_7(IN1, IN2, Out);
  input [6:0] IN1;
  input [6:0] IN2;
  output [7:0] Out;
  wire w15;
  wire w17;
  wire w19;
  wire w21;
  wire w23;
  wire w25;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w15);
  FullAdder U1 (IN1[1], IN2[1], w15, Out[1], w17);
  FullAdder U2 (IN1[2], IN2[2], w17, Out[2], w19);
  FullAdder U3 (IN1[3], IN2[3], w19, Out[3], w21);
  FullAdder U4 (IN1[4], IN2[4], w21, Out[4], w23);
  FullAdder U5 (IN1[5], IN2[5], w23, Out[5], w25);
  FullAdder U6 (IN1[6], IN2[6], w25, Out[6], Out[7]);

endmodule
module NR_35_8(IN1, IN2, Out);
  input [34:0] IN1;
  input [7:0] IN2;
  output [42:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [7:0] P8;
  wire [7:0] P9;
  wire [7:0] P10;
  wire [7:0] P11;
  wire [7:0] P12;
  wire [7:0] P13;
  wire [7:0] P14;
  wire [7:0] P15;
  wire [7:0] P16;
  wire [7:0] P17;
  wire [7:0] P18;
  wire [7:0] P19;
  wire [7:0] P20;
  wire [7:0] P21;
  wire [7:0] P22;
  wire [7:0] P23;
  wire [7:0] P24;
  wire [7:0] P25;
  wire [7:0] P26;
  wire [7:0] P27;
  wire [7:0] P28;
  wire [7:0] P29;
  wire [7:0] P30;
  wire [7:0] P31;
  wire [7:0] P32;
  wire [7:0] P33;
  wire [7:0] P34;
  wire [6:0] P35;
  wire [5:0] P36;
  wire [4:0] P37;
  wire [3:0] P38;
  wire [2:0] P39;
  wire [1:0] P40;
  wire [0:0] P41;
  wire [41:0] R1;
  wire [6:0] R2;
  wire [42:0] aOut;
  U_SP_35_8 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, R1, R2);
  RC_7_7 S2 (R1[41:35], R2, aOut[42:35]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign Out = aOut[42:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
