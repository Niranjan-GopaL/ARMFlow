
module customAdder40_0(
    input [39 : 0] A,
    input [39 : 0] B,
    output [40 : 0] Sum
);

    assign Sum = A+B;

endmodule
