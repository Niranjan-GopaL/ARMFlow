
module NR_1_49(
    input [0:0]IN1,
    input [48:0]IN2,
    output [48:0]Out
);
    assign Out = IN2;
endmodule
