
module NR_46_1(
    input [45:0]IN1,
    input [0:0]IN2,
    output [45:0]Out
);
    assign Out = IN2;
endmodule
