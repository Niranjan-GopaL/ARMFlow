
module customAdder49_0(
    input [48 : 0] A,
    input [48 : 0] B,
    output [49 : 0] Sum
);

    assign Sum = A+B;

endmodule
