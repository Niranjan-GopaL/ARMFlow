
module customAdder61_0(
    input [60 : 0] A,
    input [60 : 0] B,
    output [61 : 0] Sum
);

    assign Sum = A+B;

endmodule
