
module multiplier32bit_7(
    input [31:0] A, 
    input [31:0] B, 
    output [63:0] P
);
    
    wire [26:0] A_H, B_H;
    wire [4:0] A_L, B_L;
    
    assign A_H = A[31:5];
    assign B_H = B[31:5];
    assign A_L = A[4:0];
    assign B_L = B[4:0];
    
    
    wire [53:0] P1;
    wire [31:0] P2, P3;
    wire [9:0] P4;
    
    NR_27_27 M1(A_H, B_H, P1);
    NR_27_5 M2(A_H, B_L, P2);
    NR_5_27 M3(A_L, B_H, P3);
    NR_5_5 M4(A_L, B_L, P4);
    
    wire[4:0] P4_L;
    wire[4:0] P4_H;

    wire[58:0] operand1;
    wire[32:0] operand2;
    wire[59:0] out;
    
    assign P4_L = P4[4:0];
    assign P4_H = P4[9:5];
    assign operand1 = {P1,P4_H};

    customAdder32_0 adder1(
        P2,
        P3,
        operand2
    );

    customAdder59_26 adder2(
        operand1,
        operand2,
        out
    );
    assign P = {out[58:0],P4_L};
endmodule
        