//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 6
  second input length: 54
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_6_54(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58);
  input [5:0] IN1;
  input [53:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [5:0] P6;
  output [5:0] P7;
  output [5:0] P8;
  output [5:0] P9;
  output [5:0] P10;
  output [5:0] P11;
  output [5:0] P12;
  output [5:0] P13;
  output [5:0] P14;
  output [5:0] P15;
  output [5:0] P16;
  output [5:0] P17;
  output [5:0] P18;
  output [5:0] P19;
  output [5:0] P20;
  output [5:0] P21;
  output [5:0] P22;
  output [5:0] P23;
  output [5:0] P24;
  output [5:0] P25;
  output [5:0] P26;
  output [5:0] P27;
  output [5:0] P28;
  output [5:0] P29;
  output [5:0] P30;
  output [5:0] P31;
  output [5:0] P32;
  output [5:0] P33;
  output [5:0] P34;
  output [5:0] P35;
  output [5:0] P36;
  output [5:0] P37;
  output [5:0] P38;
  output [5:0] P39;
  output [5:0] P40;
  output [5:0] P41;
  output [5:0] P42;
  output [5:0] P43;
  output [5:0] P44;
  output [5:0] P45;
  output [5:0] P46;
  output [5:0] P47;
  output [5:0] P48;
  output [5:0] P49;
  output [5:0] P50;
  output [5:0] P51;
  output [5:0] P52;
  output [5:0] P53;
  output [4:0] P54;
  output [3:0] P55;
  output [2:0] P56;
  output [1:0] P57;
  output [0:0] P58;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[0] = IN1[1]&IN2[53];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[1] = IN1[2]&IN2[52];
  assign P55[0] = IN1[2]&IN2[53];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[2] = IN1[3]&IN2[51];
  assign P55[1] = IN1[3]&IN2[52];
  assign P56[0] = IN1[3]&IN2[53];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[3] = IN1[4]&IN2[50];
  assign P55[2] = IN1[4]&IN2[51];
  assign P56[1] = IN1[4]&IN2[52];
  assign P57[0] = IN1[4]&IN2[53];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[4] = IN1[5]&IN2[49];
  assign P55[3] = IN1[5]&IN2[50];
  assign P56[2] = IN1[5]&IN2[51];
  assign P57[1] = IN1[5]&IN2[52];
  assign P58[0] = IN1[5]&IN2[53];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [5:0] IN6;
  input [5:0] IN7;
  input [5:0] IN8;
  input [5:0] IN9;
  input [5:0] IN10;
  input [5:0] IN11;
  input [5:0] IN12;
  input [5:0] IN13;
  input [5:0] IN14;
  input [5:0] IN15;
  input [5:0] IN16;
  input [5:0] IN17;
  input [5:0] IN18;
  input [5:0] IN19;
  input [5:0] IN20;
  input [5:0] IN21;
  input [5:0] IN22;
  input [5:0] IN23;
  input [5:0] IN24;
  input [5:0] IN25;
  input [5:0] IN26;
  input [5:0] IN27;
  input [5:0] IN28;
  input [5:0] IN29;
  input [5:0] IN30;
  input [5:0] IN31;
  input [5:0] IN32;
  input [5:0] IN33;
  input [5:0] IN34;
  input [5:0] IN35;
  input [5:0] IN36;
  input [5:0] IN37;
  input [5:0] IN38;
  input [5:0] IN39;
  input [5:0] IN40;
  input [5:0] IN41;
  input [5:0] IN42;
  input [5:0] IN43;
  input [5:0] IN44;
  input [5:0] IN45;
  input [5:0] IN46;
  input [5:0] IN47;
  input [5:0] IN48;
  input [5:0] IN49;
  input [5:0] IN50;
  input [5:0] IN51;
  input [5:0] IN52;
  input [5:0] IN53;
  input [4:0] IN54;
  input [3:0] IN55;
  input [2:0] IN56;
  input [1:0] IN57;
  input [0:0] IN58;
  output [58:0] Out1;
  output [52:0] Out2;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w845;
  wire w847;
  wire w849;
  wire w851;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w325);
  FullAdder U1 (w325, IN2[0], IN2[1], w326, w327);
  FullAdder U2 (w327, IN3[0], IN3[1], w328, w329);
  FullAdder U3 (w329, IN4[0], IN4[1], w330, w331);
  FullAdder U4 (w331, IN5[0], IN5[1], w332, w333);
  HalfAdder U5 (w326, IN2[2], Out1[2], w335);
  FullAdder U6 (w335, w328, IN3[2], w336, w337);
  FullAdder U7 (w337, w330, IN4[2], w338, w339);
  FullAdder U8 (w339, w332, IN5[2], w340, w341);
  FullAdder U9 (w341, w333, IN6[0], w342, w343);
  HalfAdder U10 (w336, IN3[3], Out1[3], w345);
  FullAdder U11 (w345, w338, IN4[3], w346, w347);
  FullAdder U12 (w347, w340, IN5[3], w348, w349);
  FullAdder U13 (w349, w342, IN6[1], w350, w351);
  FullAdder U14 (w351, w343, IN7[0], w352, w353);
  HalfAdder U15 (w346, IN4[4], Out1[4], w355);
  FullAdder U16 (w355, w348, IN5[4], w356, w357);
  FullAdder U17 (w357, w350, IN6[2], w358, w359);
  FullAdder U18 (w359, w352, IN7[1], w360, w361);
  FullAdder U19 (w361, w353, IN8[0], w362, w363);
  HalfAdder U20 (w356, IN5[5], Out1[5], w365);
  FullAdder U21 (w365, w358, IN6[3], w366, w367);
  FullAdder U22 (w367, w360, IN7[2], w368, w369);
  FullAdder U23 (w369, w362, IN8[1], w370, w371);
  FullAdder U24 (w371, w363, IN9[0], w372, w373);
  HalfAdder U25 (w366, IN6[4], Out1[6], w375);
  FullAdder U26 (w375, w368, IN7[3], w376, w377);
  FullAdder U27 (w377, w370, IN8[2], w378, w379);
  FullAdder U28 (w379, w372, IN9[1], w380, w381);
  FullAdder U29 (w381, w373, IN10[0], w382, w383);
  HalfAdder U30 (w376, IN7[4], Out1[7], w385);
  FullAdder U31 (w385, w378, IN8[3], w386, w387);
  FullAdder U32 (w387, w380, IN9[2], w388, w389);
  FullAdder U33 (w389, w382, IN10[1], w390, w391);
  FullAdder U34 (w391, w383, IN11[0], w392, w393);
  HalfAdder U35 (w386, IN8[4], Out1[8], w395);
  FullAdder U36 (w395, w388, IN9[3], w396, w397);
  FullAdder U37 (w397, w390, IN10[2], w398, w399);
  FullAdder U38 (w399, w392, IN11[1], w400, w401);
  FullAdder U39 (w401, w393, IN12[0], w402, w403);
  HalfAdder U40 (w396, IN9[4], Out1[9], w405);
  FullAdder U41 (w405, w398, IN10[3], w406, w407);
  FullAdder U42 (w407, w400, IN11[2], w408, w409);
  FullAdder U43 (w409, w402, IN12[1], w410, w411);
  FullAdder U44 (w411, w403, IN13[0], w412, w413);
  HalfAdder U45 (w406, IN10[4], Out1[10], w415);
  FullAdder U46 (w415, w408, IN11[3], w416, w417);
  FullAdder U47 (w417, w410, IN12[2], w418, w419);
  FullAdder U48 (w419, w412, IN13[1], w420, w421);
  FullAdder U49 (w421, w413, IN14[0], w422, w423);
  HalfAdder U50 (w416, IN11[4], Out1[11], w425);
  FullAdder U51 (w425, w418, IN12[3], w426, w427);
  FullAdder U52 (w427, w420, IN13[2], w428, w429);
  FullAdder U53 (w429, w422, IN14[1], w430, w431);
  FullAdder U54 (w431, w423, IN15[0], w432, w433);
  HalfAdder U55 (w426, IN12[4], Out1[12], w435);
  FullAdder U56 (w435, w428, IN13[3], w436, w437);
  FullAdder U57 (w437, w430, IN14[2], w438, w439);
  FullAdder U58 (w439, w432, IN15[1], w440, w441);
  FullAdder U59 (w441, w433, IN16[0], w442, w443);
  HalfAdder U60 (w436, IN13[4], Out1[13], w445);
  FullAdder U61 (w445, w438, IN14[3], w446, w447);
  FullAdder U62 (w447, w440, IN15[2], w448, w449);
  FullAdder U63 (w449, w442, IN16[1], w450, w451);
  FullAdder U64 (w451, w443, IN17[0], w452, w453);
  HalfAdder U65 (w446, IN14[4], Out1[14], w455);
  FullAdder U66 (w455, w448, IN15[3], w456, w457);
  FullAdder U67 (w457, w450, IN16[2], w458, w459);
  FullAdder U68 (w459, w452, IN17[1], w460, w461);
  FullAdder U69 (w461, w453, IN18[0], w462, w463);
  HalfAdder U70 (w456, IN15[4], Out1[15], w465);
  FullAdder U71 (w465, w458, IN16[3], w466, w467);
  FullAdder U72 (w467, w460, IN17[2], w468, w469);
  FullAdder U73 (w469, w462, IN18[1], w470, w471);
  FullAdder U74 (w471, w463, IN19[0], w472, w473);
  HalfAdder U75 (w466, IN16[4], Out1[16], w475);
  FullAdder U76 (w475, w468, IN17[3], w476, w477);
  FullAdder U77 (w477, w470, IN18[2], w478, w479);
  FullAdder U78 (w479, w472, IN19[1], w480, w481);
  FullAdder U79 (w481, w473, IN20[0], w482, w483);
  HalfAdder U80 (w476, IN17[4], Out1[17], w485);
  FullAdder U81 (w485, w478, IN18[3], w486, w487);
  FullAdder U82 (w487, w480, IN19[2], w488, w489);
  FullAdder U83 (w489, w482, IN20[1], w490, w491);
  FullAdder U84 (w491, w483, IN21[0], w492, w493);
  HalfAdder U85 (w486, IN18[4], Out1[18], w495);
  FullAdder U86 (w495, w488, IN19[3], w496, w497);
  FullAdder U87 (w497, w490, IN20[2], w498, w499);
  FullAdder U88 (w499, w492, IN21[1], w500, w501);
  FullAdder U89 (w501, w493, IN22[0], w502, w503);
  HalfAdder U90 (w496, IN19[4], Out1[19], w505);
  FullAdder U91 (w505, w498, IN20[3], w506, w507);
  FullAdder U92 (w507, w500, IN21[2], w508, w509);
  FullAdder U93 (w509, w502, IN22[1], w510, w511);
  FullAdder U94 (w511, w503, IN23[0], w512, w513);
  HalfAdder U95 (w506, IN20[4], Out1[20], w515);
  FullAdder U96 (w515, w508, IN21[3], w516, w517);
  FullAdder U97 (w517, w510, IN22[2], w518, w519);
  FullAdder U98 (w519, w512, IN23[1], w520, w521);
  FullAdder U99 (w521, w513, IN24[0], w522, w523);
  HalfAdder U100 (w516, IN21[4], Out1[21], w525);
  FullAdder U101 (w525, w518, IN22[3], w526, w527);
  FullAdder U102 (w527, w520, IN23[2], w528, w529);
  FullAdder U103 (w529, w522, IN24[1], w530, w531);
  FullAdder U104 (w531, w523, IN25[0], w532, w533);
  HalfAdder U105 (w526, IN22[4], Out1[22], w535);
  FullAdder U106 (w535, w528, IN23[3], w536, w537);
  FullAdder U107 (w537, w530, IN24[2], w538, w539);
  FullAdder U108 (w539, w532, IN25[1], w540, w541);
  FullAdder U109 (w541, w533, IN26[0], w542, w543);
  HalfAdder U110 (w536, IN23[4], Out1[23], w545);
  FullAdder U111 (w545, w538, IN24[3], w546, w547);
  FullAdder U112 (w547, w540, IN25[2], w548, w549);
  FullAdder U113 (w549, w542, IN26[1], w550, w551);
  FullAdder U114 (w551, w543, IN27[0], w552, w553);
  HalfAdder U115 (w546, IN24[4], Out1[24], w555);
  FullAdder U116 (w555, w548, IN25[3], w556, w557);
  FullAdder U117 (w557, w550, IN26[2], w558, w559);
  FullAdder U118 (w559, w552, IN27[1], w560, w561);
  FullAdder U119 (w561, w553, IN28[0], w562, w563);
  HalfAdder U120 (w556, IN25[4], Out1[25], w565);
  FullAdder U121 (w565, w558, IN26[3], w566, w567);
  FullAdder U122 (w567, w560, IN27[2], w568, w569);
  FullAdder U123 (w569, w562, IN28[1], w570, w571);
  FullAdder U124 (w571, w563, IN29[0], w572, w573);
  HalfAdder U125 (w566, IN26[4], Out1[26], w575);
  FullAdder U126 (w575, w568, IN27[3], w576, w577);
  FullAdder U127 (w577, w570, IN28[2], w578, w579);
  FullAdder U128 (w579, w572, IN29[1], w580, w581);
  FullAdder U129 (w581, w573, IN30[0], w582, w583);
  HalfAdder U130 (w576, IN27[4], Out1[27], w585);
  FullAdder U131 (w585, w578, IN28[3], w586, w587);
  FullAdder U132 (w587, w580, IN29[2], w588, w589);
  FullAdder U133 (w589, w582, IN30[1], w590, w591);
  FullAdder U134 (w591, w583, IN31[0], w592, w593);
  HalfAdder U135 (w586, IN28[4], Out1[28], w595);
  FullAdder U136 (w595, w588, IN29[3], w596, w597);
  FullAdder U137 (w597, w590, IN30[2], w598, w599);
  FullAdder U138 (w599, w592, IN31[1], w600, w601);
  FullAdder U139 (w601, w593, IN32[0], w602, w603);
  HalfAdder U140 (w596, IN29[4], Out1[29], w605);
  FullAdder U141 (w605, w598, IN30[3], w606, w607);
  FullAdder U142 (w607, w600, IN31[2], w608, w609);
  FullAdder U143 (w609, w602, IN32[1], w610, w611);
  FullAdder U144 (w611, w603, IN33[0], w612, w613);
  HalfAdder U145 (w606, IN30[4], Out1[30], w615);
  FullAdder U146 (w615, w608, IN31[3], w616, w617);
  FullAdder U147 (w617, w610, IN32[2], w618, w619);
  FullAdder U148 (w619, w612, IN33[1], w620, w621);
  FullAdder U149 (w621, w613, IN34[0], w622, w623);
  HalfAdder U150 (w616, IN31[4], Out1[31], w625);
  FullAdder U151 (w625, w618, IN32[3], w626, w627);
  FullAdder U152 (w627, w620, IN33[2], w628, w629);
  FullAdder U153 (w629, w622, IN34[1], w630, w631);
  FullAdder U154 (w631, w623, IN35[0], w632, w633);
  HalfAdder U155 (w626, IN32[4], Out1[32], w635);
  FullAdder U156 (w635, w628, IN33[3], w636, w637);
  FullAdder U157 (w637, w630, IN34[2], w638, w639);
  FullAdder U158 (w639, w632, IN35[1], w640, w641);
  FullAdder U159 (w641, w633, IN36[0], w642, w643);
  HalfAdder U160 (w636, IN33[4], Out1[33], w645);
  FullAdder U161 (w645, w638, IN34[3], w646, w647);
  FullAdder U162 (w647, w640, IN35[2], w648, w649);
  FullAdder U163 (w649, w642, IN36[1], w650, w651);
  FullAdder U164 (w651, w643, IN37[0], w652, w653);
  HalfAdder U165 (w646, IN34[4], Out1[34], w655);
  FullAdder U166 (w655, w648, IN35[3], w656, w657);
  FullAdder U167 (w657, w650, IN36[2], w658, w659);
  FullAdder U168 (w659, w652, IN37[1], w660, w661);
  FullAdder U169 (w661, w653, IN38[0], w662, w663);
  HalfAdder U170 (w656, IN35[4], Out1[35], w665);
  FullAdder U171 (w665, w658, IN36[3], w666, w667);
  FullAdder U172 (w667, w660, IN37[2], w668, w669);
  FullAdder U173 (w669, w662, IN38[1], w670, w671);
  FullAdder U174 (w671, w663, IN39[0], w672, w673);
  HalfAdder U175 (w666, IN36[4], Out1[36], w675);
  FullAdder U176 (w675, w668, IN37[3], w676, w677);
  FullAdder U177 (w677, w670, IN38[2], w678, w679);
  FullAdder U178 (w679, w672, IN39[1], w680, w681);
  FullAdder U179 (w681, w673, IN40[0], w682, w683);
  HalfAdder U180 (w676, IN37[4], Out1[37], w685);
  FullAdder U181 (w685, w678, IN38[3], w686, w687);
  FullAdder U182 (w687, w680, IN39[2], w688, w689);
  FullAdder U183 (w689, w682, IN40[1], w690, w691);
  FullAdder U184 (w691, w683, IN41[0], w692, w693);
  HalfAdder U185 (w686, IN38[4], Out1[38], w695);
  FullAdder U186 (w695, w688, IN39[3], w696, w697);
  FullAdder U187 (w697, w690, IN40[2], w698, w699);
  FullAdder U188 (w699, w692, IN41[1], w700, w701);
  FullAdder U189 (w701, w693, IN42[0], w702, w703);
  HalfAdder U190 (w696, IN39[4], Out1[39], w705);
  FullAdder U191 (w705, w698, IN40[3], w706, w707);
  FullAdder U192 (w707, w700, IN41[2], w708, w709);
  FullAdder U193 (w709, w702, IN42[1], w710, w711);
  FullAdder U194 (w711, w703, IN43[0], w712, w713);
  HalfAdder U195 (w706, IN40[4], Out1[40], w715);
  FullAdder U196 (w715, w708, IN41[3], w716, w717);
  FullAdder U197 (w717, w710, IN42[2], w718, w719);
  FullAdder U198 (w719, w712, IN43[1], w720, w721);
  FullAdder U199 (w721, w713, IN44[0], w722, w723);
  HalfAdder U200 (w716, IN41[4], Out1[41], w725);
  FullAdder U201 (w725, w718, IN42[3], w726, w727);
  FullAdder U202 (w727, w720, IN43[2], w728, w729);
  FullAdder U203 (w729, w722, IN44[1], w730, w731);
  FullAdder U204 (w731, w723, IN45[0], w732, w733);
  HalfAdder U205 (w726, IN42[4], Out1[42], w735);
  FullAdder U206 (w735, w728, IN43[3], w736, w737);
  FullAdder U207 (w737, w730, IN44[2], w738, w739);
  FullAdder U208 (w739, w732, IN45[1], w740, w741);
  FullAdder U209 (w741, w733, IN46[0], w742, w743);
  HalfAdder U210 (w736, IN43[4], Out1[43], w745);
  FullAdder U211 (w745, w738, IN44[3], w746, w747);
  FullAdder U212 (w747, w740, IN45[2], w748, w749);
  FullAdder U213 (w749, w742, IN46[1], w750, w751);
  FullAdder U214 (w751, w743, IN47[0], w752, w753);
  HalfAdder U215 (w746, IN44[4], Out1[44], w755);
  FullAdder U216 (w755, w748, IN45[3], w756, w757);
  FullAdder U217 (w757, w750, IN46[2], w758, w759);
  FullAdder U218 (w759, w752, IN47[1], w760, w761);
  FullAdder U219 (w761, w753, IN48[0], w762, w763);
  HalfAdder U220 (w756, IN45[4], Out1[45], w765);
  FullAdder U221 (w765, w758, IN46[3], w766, w767);
  FullAdder U222 (w767, w760, IN47[2], w768, w769);
  FullAdder U223 (w769, w762, IN48[1], w770, w771);
  FullAdder U224 (w771, w763, IN49[0], w772, w773);
  HalfAdder U225 (w766, IN46[4], Out1[46], w775);
  FullAdder U226 (w775, w768, IN47[3], w776, w777);
  FullAdder U227 (w777, w770, IN48[2], w778, w779);
  FullAdder U228 (w779, w772, IN49[1], w780, w781);
  FullAdder U229 (w781, w773, IN50[0], w782, w783);
  HalfAdder U230 (w776, IN47[4], Out1[47], w785);
  FullAdder U231 (w785, w778, IN48[3], w786, w787);
  FullAdder U232 (w787, w780, IN49[2], w788, w789);
  FullAdder U233 (w789, w782, IN50[1], w790, w791);
  FullAdder U234 (w791, w783, IN51[0], w792, w793);
  HalfAdder U235 (w786, IN48[4], Out1[48], w795);
  FullAdder U236 (w795, w788, IN49[3], w796, w797);
  FullAdder U237 (w797, w790, IN50[2], w798, w799);
  FullAdder U238 (w799, w792, IN51[1], w800, w801);
  FullAdder U239 (w801, w793, IN52[0], w802, w803);
  HalfAdder U240 (w796, IN49[4], Out1[49], w805);
  FullAdder U241 (w805, w798, IN50[3], w806, w807);
  FullAdder U242 (w807, w800, IN51[2], w808, w809);
  FullAdder U243 (w809, w802, IN52[1], w810, w811);
  FullAdder U244 (w811, w803, IN53[0], w812, w813);
  HalfAdder U245 (w806, IN50[4], Out1[50], w815);
  FullAdder U246 (w815, w808, IN51[3], w816, w817);
  FullAdder U247 (w817, w810, IN52[2], w818, w819);
  FullAdder U248 (w819, w812, IN53[1], w820, w821);
  FullAdder U249 (w821, w813, IN54[0], w822, w823);
  HalfAdder U250 (w816, IN51[4], Out1[51], w825);
  FullAdder U251 (w825, w818, IN52[3], w826, w827);
  FullAdder U252 (w827, w820, IN53[2], w828, w829);
  FullAdder U253 (w829, w822, IN54[1], w830, w831);
  FullAdder U254 (w831, w823, IN55[0], w832, w833);
  HalfAdder U255 (w826, IN52[4], Out1[52], w835);
  FullAdder U256 (w835, w828, IN53[3], w836, w837);
  FullAdder U257 (w837, w830, IN54[2], w838, w839);
  FullAdder U258 (w839, w832, IN55[1], w840, w841);
  FullAdder U259 (w841, w833, IN56[0], w842, w843);
  HalfAdder U260 (w836, IN53[4], Out1[53], w845);
  FullAdder U261 (w845, w838, IN54[3], Out1[54], w847);
  FullAdder U262 (w847, w840, IN55[2], Out1[55], w849);
  FullAdder U263 (w849, w842, IN56[1], Out1[56], w851);
  FullAdder U264 (w851, w843, IN57[0], Out1[57], Out1[58]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN6[5];
  assign Out2[1] = IN7[5];
  assign Out2[2] = IN8[5];
  assign Out2[3] = IN9[5];
  assign Out2[4] = IN10[5];
  assign Out2[5] = IN11[5];
  assign Out2[6] = IN12[5];
  assign Out2[7] = IN13[5];
  assign Out2[8] = IN14[5];
  assign Out2[9] = IN15[5];
  assign Out2[10] = IN16[5];
  assign Out2[11] = IN17[5];
  assign Out2[12] = IN18[5];
  assign Out2[13] = IN19[5];
  assign Out2[14] = IN20[5];
  assign Out2[15] = IN21[5];
  assign Out2[16] = IN22[5];
  assign Out2[17] = IN23[5];
  assign Out2[18] = IN24[5];
  assign Out2[19] = IN25[5];
  assign Out2[20] = IN26[5];
  assign Out2[21] = IN27[5];
  assign Out2[22] = IN28[5];
  assign Out2[23] = IN29[5];
  assign Out2[24] = IN30[5];
  assign Out2[25] = IN31[5];
  assign Out2[26] = IN32[5];
  assign Out2[27] = IN33[5];
  assign Out2[28] = IN34[5];
  assign Out2[29] = IN35[5];
  assign Out2[30] = IN36[5];
  assign Out2[31] = IN37[5];
  assign Out2[32] = IN38[5];
  assign Out2[33] = IN39[5];
  assign Out2[34] = IN40[5];
  assign Out2[35] = IN41[5];
  assign Out2[36] = IN42[5];
  assign Out2[37] = IN43[5];
  assign Out2[38] = IN44[5];
  assign Out2[39] = IN45[5];
  assign Out2[40] = IN46[5];
  assign Out2[41] = IN47[5];
  assign Out2[42] = IN48[5];
  assign Out2[43] = IN49[5];
  assign Out2[44] = IN50[5];
  assign Out2[45] = IN51[5];
  assign Out2[46] = IN52[5];
  assign Out2[47] = IN53[5];
  assign Out2[48] = IN54[4];
  assign Out2[49] = IN55[3];
  assign Out2[50] = IN56[2];
  assign Out2[51] = IN57[1];
  assign Out2[52] = IN58[0];

endmodule
module RC_53_53(IN1, IN2, Out);
  input [52:0] IN1;
  input [52:0] IN2;
  output [53:0] Out;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w107);
  FullAdder U1 (IN1[1], IN2[1], w107, Out[1], w109);
  FullAdder U2 (IN1[2], IN2[2], w109, Out[2], w111);
  FullAdder U3 (IN1[3], IN2[3], w111, Out[3], w113);
  FullAdder U4 (IN1[4], IN2[4], w113, Out[4], w115);
  FullAdder U5 (IN1[5], IN2[5], w115, Out[5], w117);
  FullAdder U6 (IN1[6], IN2[6], w117, Out[6], w119);
  FullAdder U7 (IN1[7], IN2[7], w119, Out[7], w121);
  FullAdder U8 (IN1[8], IN2[8], w121, Out[8], w123);
  FullAdder U9 (IN1[9], IN2[9], w123, Out[9], w125);
  FullAdder U10 (IN1[10], IN2[10], w125, Out[10], w127);
  FullAdder U11 (IN1[11], IN2[11], w127, Out[11], w129);
  FullAdder U12 (IN1[12], IN2[12], w129, Out[12], w131);
  FullAdder U13 (IN1[13], IN2[13], w131, Out[13], w133);
  FullAdder U14 (IN1[14], IN2[14], w133, Out[14], w135);
  FullAdder U15 (IN1[15], IN2[15], w135, Out[15], w137);
  FullAdder U16 (IN1[16], IN2[16], w137, Out[16], w139);
  FullAdder U17 (IN1[17], IN2[17], w139, Out[17], w141);
  FullAdder U18 (IN1[18], IN2[18], w141, Out[18], w143);
  FullAdder U19 (IN1[19], IN2[19], w143, Out[19], w145);
  FullAdder U20 (IN1[20], IN2[20], w145, Out[20], w147);
  FullAdder U21 (IN1[21], IN2[21], w147, Out[21], w149);
  FullAdder U22 (IN1[22], IN2[22], w149, Out[22], w151);
  FullAdder U23 (IN1[23], IN2[23], w151, Out[23], w153);
  FullAdder U24 (IN1[24], IN2[24], w153, Out[24], w155);
  FullAdder U25 (IN1[25], IN2[25], w155, Out[25], w157);
  FullAdder U26 (IN1[26], IN2[26], w157, Out[26], w159);
  FullAdder U27 (IN1[27], IN2[27], w159, Out[27], w161);
  FullAdder U28 (IN1[28], IN2[28], w161, Out[28], w163);
  FullAdder U29 (IN1[29], IN2[29], w163, Out[29], w165);
  FullAdder U30 (IN1[30], IN2[30], w165, Out[30], w167);
  FullAdder U31 (IN1[31], IN2[31], w167, Out[31], w169);
  FullAdder U32 (IN1[32], IN2[32], w169, Out[32], w171);
  FullAdder U33 (IN1[33], IN2[33], w171, Out[33], w173);
  FullAdder U34 (IN1[34], IN2[34], w173, Out[34], w175);
  FullAdder U35 (IN1[35], IN2[35], w175, Out[35], w177);
  FullAdder U36 (IN1[36], IN2[36], w177, Out[36], w179);
  FullAdder U37 (IN1[37], IN2[37], w179, Out[37], w181);
  FullAdder U38 (IN1[38], IN2[38], w181, Out[38], w183);
  FullAdder U39 (IN1[39], IN2[39], w183, Out[39], w185);
  FullAdder U40 (IN1[40], IN2[40], w185, Out[40], w187);
  FullAdder U41 (IN1[41], IN2[41], w187, Out[41], w189);
  FullAdder U42 (IN1[42], IN2[42], w189, Out[42], w191);
  FullAdder U43 (IN1[43], IN2[43], w191, Out[43], w193);
  FullAdder U44 (IN1[44], IN2[44], w193, Out[44], w195);
  FullAdder U45 (IN1[45], IN2[45], w195, Out[45], w197);
  FullAdder U46 (IN1[46], IN2[46], w197, Out[46], w199);
  FullAdder U47 (IN1[47], IN2[47], w199, Out[47], w201);
  FullAdder U48 (IN1[48], IN2[48], w201, Out[48], w203);
  FullAdder U49 (IN1[49], IN2[49], w203, Out[49], w205);
  FullAdder U50 (IN1[50], IN2[50], w205, Out[50], w207);
  FullAdder U51 (IN1[51], IN2[51], w207, Out[51], w209);
  FullAdder U52 (IN1[52], IN2[52], w209, Out[52], Out[53]);

endmodule
module NR_6_54(IN1, IN2, Out);
  input [5:0] IN1;
  input [53:0] IN2;
  output [59:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [5:0] P6;
  wire [5:0] P7;
  wire [5:0] P8;
  wire [5:0] P9;
  wire [5:0] P10;
  wire [5:0] P11;
  wire [5:0] P12;
  wire [5:0] P13;
  wire [5:0] P14;
  wire [5:0] P15;
  wire [5:0] P16;
  wire [5:0] P17;
  wire [5:0] P18;
  wire [5:0] P19;
  wire [5:0] P20;
  wire [5:0] P21;
  wire [5:0] P22;
  wire [5:0] P23;
  wire [5:0] P24;
  wire [5:0] P25;
  wire [5:0] P26;
  wire [5:0] P27;
  wire [5:0] P28;
  wire [5:0] P29;
  wire [5:0] P30;
  wire [5:0] P31;
  wire [5:0] P32;
  wire [5:0] P33;
  wire [5:0] P34;
  wire [5:0] P35;
  wire [5:0] P36;
  wire [5:0] P37;
  wire [5:0] P38;
  wire [5:0] P39;
  wire [5:0] P40;
  wire [5:0] P41;
  wire [5:0] P42;
  wire [5:0] P43;
  wire [5:0] P44;
  wire [5:0] P45;
  wire [5:0] P46;
  wire [5:0] P47;
  wire [5:0] P48;
  wire [5:0] P49;
  wire [5:0] P50;
  wire [5:0] P51;
  wire [5:0] P52;
  wire [5:0] P53;
  wire [4:0] P54;
  wire [3:0] P55;
  wire [2:0] P56;
  wire [1:0] P57;
  wire [0:0] P58;
  wire [58:0] R1;
  wire [52:0] R2;
  wire [59:0] aOut;
  U_SP_6_54 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, R1, R2);
  RC_53_53 S2 (R1[58:6], R2, aOut[59:6]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign Out = aOut[59:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
