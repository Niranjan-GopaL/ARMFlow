//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 48
  second input length: 29
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_48_29(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75);
  input [47:0] IN1;
  input [28:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [28:0] P29;
  output [28:0] P30;
  output [28:0] P31;
  output [28:0] P32;
  output [28:0] P33;
  output [28:0] P34;
  output [28:0] P35;
  output [28:0] P36;
  output [28:0] P37;
  output [28:0] P38;
  output [28:0] P39;
  output [28:0] P40;
  output [28:0] P41;
  output [28:0] P42;
  output [28:0] P43;
  output [28:0] P44;
  output [28:0] P45;
  output [28:0] P46;
  output [28:0] P47;
  output [27:0] P48;
  output [26:0] P49;
  output [25:0] P50;
  output [24:0] P51;
  output [23:0] P52;
  output [22:0] P53;
  output [21:0] P54;
  output [20:0] P55;
  output [19:0] P56;
  output [18:0] P57;
  output [17:0] P58;
  output [16:0] P59;
  output [15:0] P60;
  output [14:0] P61;
  output [13:0] P62;
  output [12:0] P63;
  output [11:0] P64;
  output [10:0] P65;
  output [9:0] P66;
  output [8:0] P67;
  output [7:0] P68;
  output [6:0] P69;
  output [5:0] P70;
  output [4:0] P71;
  output [3:0] P72;
  output [2:0] P73;
  output [1:0] P74;
  output [0:0] P75;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[0] = IN1[1]&IN2[28];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[1] = IN1[2]&IN2[27];
  assign P30[0] = IN1[2]&IN2[28];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[2] = IN1[3]&IN2[26];
  assign P30[1] = IN1[3]&IN2[27];
  assign P31[0] = IN1[3]&IN2[28];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[3] = IN1[4]&IN2[25];
  assign P30[2] = IN1[4]&IN2[26];
  assign P31[1] = IN1[4]&IN2[27];
  assign P32[0] = IN1[4]&IN2[28];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[4] = IN1[5]&IN2[24];
  assign P30[3] = IN1[5]&IN2[25];
  assign P31[2] = IN1[5]&IN2[26];
  assign P32[1] = IN1[5]&IN2[27];
  assign P33[0] = IN1[5]&IN2[28];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[5] = IN1[6]&IN2[23];
  assign P30[4] = IN1[6]&IN2[24];
  assign P31[3] = IN1[6]&IN2[25];
  assign P32[2] = IN1[6]&IN2[26];
  assign P33[1] = IN1[6]&IN2[27];
  assign P34[0] = IN1[6]&IN2[28];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[6] = IN1[7]&IN2[22];
  assign P30[5] = IN1[7]&IN2[23];
  assign P31[4] = IN1[7]&IN2[24];
  assign P32[3] = IN1[7]&IN2[25];
  assign P33[2] = IN1[7]&IN2[26];
  assign P34[1] = IN1[7]&IN2[27];
  assign P35[0] = IN1[7]&IN2[28];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[7] = IN1[8]&IN2[21];
  assign P30[6] = IN1[8]&IN2[22];
  assign P31[5] = IN1[8]&IN2[23];
  assign P32[4] = IN1[8]&IN2[24];
  assign P33[3] = IN1[8]&IN2[25];
  assign P34[2] = IN1[8]&IN2[26];
  assign P35[1] = IN1[8]&IN2[27];
  assign P36[0] = IN1[8]&IN2[28];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[8] = IN1[9]&IN2[20];
  assign P30[7] = IN1[9]&IN2[21];
  assign P31[6] = IN1[9]&IN2[22];
  assign P32[5] = IN1[9]&IN2[23];
  assign P33[4] = IN1[9]&IN2[24];
  assign P34[3] = IN1[9]&IN2[25];
  assign P35[2] = IN1[9]&IN2[26];
  assign P36[1] = IN1[9]&IN2[27];
  assign P37[0] = IN1[9]&IN2[28];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[9] = IN1[10]&IN2[19];
  assign P30[8] = IN1[10]&IN2[20];
  assign P31[7] = IN1[10]&IN2[21];
  assign P32[6] = IN1[10]&IN2[22];
  assign P33[5] = IN1[10]&IN2[23];
  assign P34[4] = IN1[10]&IN2[24];
  assign P35[3] = IN1[10]&IN2[25];
  assign P36[2] = IN1[10]&IN2[26];
  assign P37[1] = IN1[10]&IN2[27];
  assign P38[0] = IN1[10]&IN2[28];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[10] = IN1[11]&IN2[18];
  assign P30[9] = IN1[11]&IN2[19];
  assign P31[8] = IN1[11]&IN2[20];
  assign P32[7] = IN1[11]&IN2[21];
  assign P33[6] = IN1[11]&IN2[22];
  assign P34[5] = IN1[11]&IN2[23];
  assign P35[4] = IN1[11]&IN2[24];
  assign P36[3] = IN1[11]&IN2[25];
  assign P37[2] = IN1[11]&IN2[26];
  assign P38[1] = IN1[11]&IN2[27];
  assign P39[0] = IN1[11]&IN2[28];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[11] = IN1[12]&IN2[17];
  assign P30[10] = IN1[12]&IN2[18];
  assign P31[9] = IN1[12]&IN2[19];
  assign P32[8] = IN1[12]&IN2[20];
  assign P33[7] = IN1[12]&IN2[21];
  assign P34[6] = IN1[12]&IN2[22];
  assign P35[5] = IN1[12]&IN2[23];
  assign P36[4] = IN1[12]&IN2[24];
  assign P37[3] = IN1[12]&IN2[25];
  assign P38[2] = IN1[12]&IN2[26];
  assign P39[1] = IN1[12]&IN2[27];
  assign P40[0] = IN1[12]&IN2[28];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[12] = IN1[13]&IN2[16];
  assign P30[11] = IN1[13]&IN2[17];
  assign P31[10] = IN1[13]&IN2[18];
  assign P32[9] = IN1[13]&IN2[19];
  assign P33[8] = IN1[13]&IN2[20];
  assign P34[7] = IN1[13]&IN2[21];
  assign P35[6] = IN1[13]&IN2[22];
  assign P36[5] = IN1[13]&IN2[23];
  assign P37[4] = IN1[13]&IN2[24];
  assign P38[3] = IN1[13]&IN2[25];
  assign P39[2] = IN1[13]&IN2[26];
  assign P40[1] = IN1[13]&IN2[27];
  assign P41[0] = IN1[13]&IN2[28];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[13] = IN1[14]&IN2[15];
  assign P30[12] = IN1[14]&IN2[16];
  assign P31[11] = IN1[14]&IN2[17];
  assign P32[10] = IN1[14]&IN2[18];
  assign P33[9] = IN1[14]&IN2[19];
  assign P34[8] = IN1[14]&IN2[20];
  assign P35[7] = IN1[14]&IN2[21];
  assign P36[6] = IN1[14]&IN2[22];
  assign P37[5] = IN1[14]&IN2[23];
  assign P38[4] = IN1[14]&IN2[24];
  assign P39[3] = IN1[14]&IN2[25];
  assign P40[2] = IN1[14]&IN2[26];
  assign P41[1] = IN1[14]&IN2[27];
  assign P42[0] = IN1[14]&IN2[28];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[14] = IN1[15]&IN2[14];
  assign P30[13] = IN1[15]&IN2[15];
  assign P31[12] = IN1[15]&IN2[16];
  assign P32[11] = IN1[15]&IN2[17];
  assign P33[10] = IN1[15]&IN2[18];
  assign P34[9] = IN1[15]&IN2[19];
  assign P35[8] = IN1[15]&IN2[20];
  assign P36[7] = IN1[15]&IN2[21];
  assign P37[6] = IN1[15]&IN2[22];
  assign P38[5] = IN1[15]&IN2[23];
  assign P39[4] = IN1[15]&IN2[24];
  assign P40[3] = IN1[15]&IN2[25];
  assign P41[2] = IN1[15]&IN2[26];
  assign P42[1] = IN1[15]&IN2[27];
  assign P43[0] = IN1[15]&IN2[28];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[15] = IN1[16]&IN2[13];
  assign P30[14] = IN1[16]&IN2[14];
  assign P31[13] = IN1[16]&IN2[15];
  assign P32[12] = IN1[16]&IN2[16];
  assign P33[11] = IN1[16]&IN2[17];
  assign P34[10] = IN1[16]&IN2[18];
  assign P35[9] = IN1[16]&IN2[19];
  assign P36[8] = IN1[16]&IN2[20];
  assign P37[7] = IN1[16]&IN2[21];
  assign P38[6] = IN1[16]&IN2[22];
  assign P39[5] = IN1[16]&IN2[23];
  assign P40[4] = IN1[16]&IN2[24];
  assign P41[3] = IN1[16]&IN2[25];
  assign P42[2] = IN1[16]&IN2[26];
  assign P43[1] = IN1[16]&IN2[27];
  assign P44[0] = IN1[16]&IN2[28];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[16] = IN1[17]&IN2[12];
  assign P30[15] = IN1[17]&IN2[13];
  assign P31[14] = IN1[17]&IN2[14];
  assign P32[13] = IN1[17]&IN2[15];
  assign P33[12] = IN1[17]&IN2[16];
  assign P34[11] = IN1[17]&IN2[17];
  assign P35[10] = IN1[17]&IN2[18];
  assign P36[9] = IN1[17]&IN2[19];
  assign P37[8] = IN1[17]&IN2[20];
  assign P38[7] = IN1[17]&IN2[21];
  assign P39[6] = IN1[17]&IN2[22];
  assign P40[5] = IN1[17]&IN2[23];
  assign P41[4] = IN1[17]&IN2[24];
  assign P42[3] = IN1[17]&IN2[25];
  assign P43[2] = IN1[17]&IN2[26];
  assign P44[1] = IN1[17]&IN2[27];
  assign P45[0] = IN1[17]&IN2[28];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[17] = IN1[18]&IN2[11];
  assign P30[16] = IN1[18]&IN2[12];
  assign P31[15] = IN1[18]&IN2[13];
  assign P32[14] = IN1[18]&IN2[14];
  assign P33[13] = IN1[18]&IN2[15];
  assign P34[12] = IN1[18]&IN2[16];
  assign P35[11] = IN1[18]&IN2[17];
  assign P36[10] = IN1[18]&IN2[18];
  assign P37[9] = IN1[18]&IN2[19];
  assign P38[8] = IN1[18]&IN2[20];
  assign P39[7] = IN1[18]&IN2[21];
  assign P40[6] = IN1[18]&IN2[22];
  assign P41[5] = IN1[18]&IN2[23];
  assign P42[4] = IN1[18]&IN2[24];
  assign P43[3] = IN1[18]&IN2[25];
  assign P44[2] = IN1[18]&IN2[26];
  assign P45[1] = IN1[18]&IN2[27];
  assign P46[0] = IN1[18]&IN2[28];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[18] = IN1[19]&IN2[10];
  assign P30[17] = IN1[19]&IN2[11];
  assign P31[16] = IN1[19]&IN2[12];
  assign P32[15] = IN1[19]&IN2[13];
  assign P33[14] = IN1[19]&IN2[14];
  assign P34[13] = IN1[19]&IN2[15];
  assign P35[12] = IN1[19]&IN2[16];
  assign P36[11] = IN1[19]&IN2[17];
  assign P37[10] = IN1[19]&IN2[18];
  assign P38[9] = IN1[19]&IN2[19];
  assign P39[8] = IN1[19]&IN2[20];
  assign P40[7] = IN1[19]&IN2[21];
  assign P41[6] = IN1[19]&IN2[22];
  assign P42[5] = IN1[19]&IN2[23];
  assign P43[4] = IN1[19]&IN2[24];
  assign P44[3] = IN1[19]&IN2[25];
  assign P45[2] = IN1[19]&IN2[26];
  assign P46[1] = IN1[19]&IN2[27];
  assign P47[0] = IN1[19]&IN2[28];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[19] = IN1[20]&IN2[9];
  assign P30[18] = IN1[20]&IN2[10];
  assign P31[17] = IN1[20]&IN2[11];
  assign P32[16] = IN1[20]&IN2[12];
  assign P33[15] = IN1[20]&IN2[13];
  assign P34[14] = IN1[20]&IN2[14];
  assign P35[13] = IN1[20]&IN2[15];
  assign P36[12] = IN1[20]&IN2[16];
  assign P37[11] = IN1[20]&IN2[17];
  assign P38[10] = IN1[20]&IN2[18];
  assign P39[9] = IN1[20]&IN2[19];
  assign P40[8] = IN1[20]&IN2[20];
  assign P41[7] = IN1[20]&IN2[21];
  assign P42[6] = IN1[20]&IN2[22];
  assign P43[5] = IN1[20]&IN2[23];
  assign P44[4] = IN1[20]&IN2[24];
  assign P45[3] = IN1[20]&IN2[25];
  assign P46[2] = IN1[20]&IN2[26];
  assign P47[1] = IN1[20]&IN2[27];
  assign P48[0] = IN1[20]&IN2[28];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[20] = IN1[21]&IN2[8];
  assign P30[19] = IN1[21]&IN2[9];
  assign P31[18] = IN1[21]&IN2[10];
  assign P32[17] = IN1[21]&IN2[11];
  assign P33[16] = IN1[21]&IN2[12];
  assign P34[15] = IN1[21]&IN2[13];
  assign P35[14] = IN1[21]&IN2[14];
  assign P36[13] = IN1[21]&IN2[15];
  assign P37[12] = IN1[21]&IN2[16];
  assign P38[11] = IN1[21]&IN2[17];
  assign P39[10] = IN1[21]&IN2[18];
  assign P40[9] = IN1[21]&IN2[19];
  assign P41[8] = IN1[21]&IN2[20];
  assign P42[7] = IN1[21]&IN2[21];
  assign P43[6] = IN1[21]&IN2[22];
  assign P44[5] = IN1[21]&IN2[23];
  assign P45[4] = IN1[21]&IN2[24];
  assign P46[3] = IN1[21]&IN2[25];
  assign P47[2] = IN1[21]&IN2[26];
  assign P48[1] = IN1[21]&IN2[27];
  assign P49[0] = IN1[21]&IN2[28];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[21] = IN1[22]&IN2[7];
  assign P30[20] = IN1[22]&IN2[8];
  assign P31[19] = IN1[22]&IN2[9];
  assign P32[18] = IN1[22]&IN2[10];
  assign P33[17] = IN1[22]&IN2[11];
  assign P34[16] = IN1[22]&IN2[12];
  assign P35[15] = IN1[22]&IN2[13];
  assign P36[14] = IN1[22]&IN2[14];
  assign P37[13] = IN1[22]&IN2[15];
  assign P38[12] = IN1[22]&IN2[16];
  assign P39[11] = IN1[22]&IN2[17];
  assign P40[10] = IN1[22]&IN2[18];
  assign P41[9] = IN1[22]&IN2[19];
  assign P42[8] = IN1[22]&IN2[20];
  assign P43[7] = IN1[22]&IN2[21];
  assign P44[6] = IN1[22]&IN2[22];
  assign P45[5] = IN1[22]&IN2[23];
  assign P46[4] = IN1[22]&IN2[24];
  assign P47[3] = IN1[22]&IN2[25];
  assign P48[2] = IN1[22]&IN2[26];
  assign P49[1] = IN1[22]&IN2[27];
  assign P50[0] = IN1[22]&IN2[28];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[22] = IN1[23]&IN2[6];
  assign P30[21] = IN1[23]&IN2[7];
  assign P31[20] = IN1[23]&IN2[8];
  assign P32[19] = IN1[23]&IN2[9];
  assign P33[18] = IN1[23]&IN2[10];
  assign P34[17] = IN1[23]&IN2[11];
  assign P35[16] = IN1[23]&IN2[12];
  assign P36[15] = IN1[23]&IN2[13];
  assign P37[14] = IN1[23]&IN2[14];
  assign P38[13] = IN1[23]&IN2[15];
  assign P39[12] = IN1[23]&IN2[16];
  assign P40[11] = IN1[23]&IN2[17];
  assign P41[10] = IN1[23]&IN2[18];
  assign P42[9] = IN1[23]&IN2[19];
  assign P43[8] = IN1[23]&IN2[20];
  assign P44[7] = IN1[23]&IN2[21];
  assign P45[6] = IN1[23]&IN2[22];
  assign P46[5] = IN1[23]&IN2[23];
  assign P47[4] = IN1[23]&IN2[24];
  assign P48[3] = IN1[23]&IN2[25];
  assign P49[2] = IN1[23]&IN2[26];
  assign P50[1] = IN1[23]&IN2[27];
  assign P51[0] = IN1[23]&IN2[28];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[23] = IN1[24]&IN2[5];
  assign P30[22] = IN1[24]&IN2[6];
  assign P31[21] = IN1[24]&IN2[7];
  assign P32[20] = IN1[24]&IN2[8];
  assign P33[19] = IN1[24]&IN2[9];
  assign P34[18] = IN1[24]&IN2[10];
  assign P35[17] = IN1[24]&IN2[11];
  assign P36[16] = IN1[24]&IN2[12];
  assign P37[15] = IN1[24]&IN2[13];
  assign P38[14] = IN1[24]&IN2[14];
  assign P39[13] = IN1[24]&IN2[15];
  assign P40[12] = IN1[24]&IN2[16];
  assign P41[11] = IN1[24]&IN2[17];
  assign P42[10] = IN1[24]&IN2[18];
  assign P43[9] = IN1[24]&IN2[19];
  assign P44[8] = IN1[24]&IN2[20];
  assign P45[7] = IN1[24]&IN2[21];
  assign P46[6] = IN1[24]&IN2[22];
  assign P47[5] = IN1[24]&IN2[23];
  assign P48[4] = IN1[24]&IN2[24];
  assign P49[3] = IN1[24]&IN2[25];
  assign P50[2] = IN1[24]&IN2[26];
  assign P51[1] = IN1[24]&IN2[27];
  assign P52[0] = IN1[24]&IN2[28];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[24] = IN1[25]&IN2[4];
  assign P30[23] = IN1[25]&IN2[5];
  assign P31[22] = IN1[25]&IN2[6];
  assign P32[21] = IN1[25]&IN2[7];
  assign P33[20] = IN1[25]&IN2[8];
  assign P34[19] = IN1[25]&IN2[9];
  assign P35[18] = IN1[25]&IN2[10];
  assign P36[17] = IN1[25]&IN2[11];
  assign P37[16] = IN1[25]&IN2[12];
  assign P38[15] = IN1[25]&IN2[13];
  assign P39[14] = IN1[25]&IN2[14];
  assign P40[13] = IN1[25]&IN2[15];
  assign P41[12] = IN1[25]&IN2[16];
  assign P42[11] = IN1[25]&IN2[17];
  assign P43[10] = IN1[25]&IN2[18];
  assign P44[9] = IN1[25]&IN2[19];
  assign P45[8] = IN1[25]&IN2[20];
  assign P46[7] = IN1[25]&IN2[21];
  assign P47[6] = IN1[25]&IN2[22];
  assign P48[5] = IN1[25]&IN2[23];
  assign P49[4] = IN1[25]&IN2[24];
  assign P50[3] = IN1[25]&IN2[25];
  assign P51[2] = IN1[25]&IN2[26];
  assign P52[1] = IN1[25]&IN2[27];
  assign P53[0] = IN1[25]&IN2[28];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[25] = IN1[26]&IN2[3];
  assign P30[24] = IN1[26]&IN2[4];
  assign P31[23] = IN1[26]&IN2[5];
  assign P32[22] = IN1[26]&IN2[6];
  assign P33[21] = IN1[26]&IN2[7];
  assign P34[20] = IN1[26]&IN2[8];
  assign P35[19] = IN1[26]&IN2[9];
  assign P36[18] = IN1[26]&IN2[10];
  assign P37[17] = IN1[26]&IN2[11];
  assign P38[16] = IN1[26]&IN2[12];
  assign P39[15] = IN1[26]&IN2[13];
  assign P40[14] = IN1[26]&IN2[14];
  assign P41[13] = IN1[26]&IN2[15];
  assign P42[12] = IN1[26]&IN2[16];
  assign P43[11] = IN1[26]&IN2[17];
  assign P44[10] = IN1[26]&IN2[18];
  assign P45[9] = IN1[26]&IN2[19];
  assign P46[8] = IN1[26]&IN2[20];
  assign P47[7] = IN1[26]&IN2[21];
  assign P48[6] = IN1[26]&IN2[22];
  assign P49[5] = IN1[26]&IN2[23];
  assign P50[4] = IN1[26]&IN2[24];
  assign P51[3] = IN1[26]&IN2[25];
  assign P52[2] = IN1[26]&IN2[26];
  assign P53[1] = IN1[26]&IN2[27];
  assign P54[0] = IN1[26]&IN2[28];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[26] = IN1[27]&IN2[2];
  assign P30[25] = IN1[27]&IN2[3];
  assign P31[24] = IN1[27]&IN2[4];
  assign P32[23] = IN1[27]&IN2[5];
  assign P33[22] = IN1[27]&IN2[6];
  assign P34[21] = IN1[27]&IN2[7];
  assign P35[20] = IN1[27]&IN2[8];
  assign P36[19] = IN1[27]&IN2[9];
  assign P37[18] = IN1[27]&IN2[10];
  assign P38[17] = IN1[27]&IN2[11];
  assign P39[16] = IN1[27]&IN2[12];
  assign P40[15] = IN1[27]&IN2[13];
  assign P41[14] = IN1[27]&IN2[14];
  assign P42[13] = IN1[27]&IN2[15];
  assign P43[12] = IN1[27]&IN2[16];
  assign P44[11] = IN1[27]&IN2[17];
  assign P45[10] = IN1[27]&IN2[18];
  assign P46[9] = IN1[27]&IN2[19];
  assign P47[8] = IN1[27]&IN2[20];
  assign P48[7] = IN1[27]&IN2[21];
  assign P49[6] = IN1[27]&IN2[22];
  assign P50[5] = IN1[27]&IN2[23];
  assign P51[4] = IN1[27]&IN2[24];
  assign P52[3] = IN1[27]&IN2[25];
  assign P53[2] = IN1[27]&IN2[26];
  assign P54[1] = IN1[27]&IN2[27];
  assign P55[0] = IN1[27]&IN2[28];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[27] = IN1[28]&IN2[1];
  assign P30[26] = IN1[28]&IN2[2];
  assign P31[25] = IN1[28]&IN2[3];
  assign P32[24] = IN1[28]&IN2[4];
  assign P33[23] = IN1[28]&IN2[5];
  assign P34[22] = IN1[28]&IN2[6];
  assign P35[21] = IN1[28]&IN2[7];
  assign P36[20] = IN1[28]&IN2[8];
  assign P37[19] = IN1[28]&IN2[9];
  assign P38[18] = IN1[28]&IN2[10];
  assign P39[17] = IN1[28]&IN2[11];
  assign P40[16] = IN1[28]&IN2[12];
  assign P41[15] = IN1[28]&IN2[13];
  assign P42[14] = IN1[28]&IN2[14];
  assign P43[13] = IN1[28]&IN2[15];
  assign P44[12] = IN1[28]&IN2[16];
  assign P45[11] = IN1[28]&IN2[17];
  assign P46[10] = IN1[28]&IN2[18];
  assign P47[9] = IN1[28]&IN2[19];
  assign P48[8] = IN1[28]&IN2[20];
  assign P49[7] = IN1[28]&IN2[21];
  assign P50[6] = IN1[28]&IN2[22];
  assign P51[5] = IN1[28]&IN2[23];
  assign P52[4] = IN1[28]&IN2[24];
  assign P53[3] = IN1[28]&IN2[25];
  assign P54[2] = IN1[28]&IN2[26];
  assign P55[1] = IN1[28]&IN2[27];
  assign P56[0] = IN1[28]&IN2[28];
  assign P29[28] = IN1[29]&IN2[0];
  assign P30[27] = IN1[29]&IN2[1];
  assign P31[26] = IN1[29]&IN2[2];
  assign P32[25] = IN1[29]&IN2[3];
  assign P33[24] = IN1[29]&IN2[4];
  assign P34[23] = IN1[29]&IN2[5];
  assign P35[22] = IN1[29]&IN2[6];
  assign P36[21] = IN1[29]&IN2[7];
  assign P37[20] = IN1[29]&IN2[8];
  assign P38[19] = IN1[29]&IN2[9];
  assign P39[18] = IN1[29]&IN2[10];
  assign P40[17] = IN1[29]&IN2[11];
  assign P41[16] = IN1[29]&IN2[12];
  assign P42[15] = IN1[29]&IN2[13];
  assign P43[14] = IN1[29]&IN2[14];
  assign P44[13] = IN1[29]&IN2[15];
  assign P45[12] = IN1[29]&IN2[16];
  assign P46[11] = IN1[29]&IN2[17];
  assign P47[10] = IN1[29]&IN2[18];
  assign P48[9] = IN1[29]&IN2[19];
  assign P49[8] = IN1[29]&IN2[20];
  assign P50[7] = IN1[29]&IN2[21];
  assign P51[6] = IN1[29]&IN2[22];
  assign P52[5] = IN1[29]&IN2[23];
  assign P53[4] = IN1[29]&IN2[24];
  assign P54[3] = IN1[29]&IN2[25];
  assign P55[2] = IN1[29]&IN2[26];
  assign P56[1] = IN1[29]&IN2[27];
  assign P57[0] = IN1[29]&IN2[28];
  assign P30[28] = IN1[30]&IN2[0];
  assign P31[27] = IN1[30]&IN2[1];
  assign P32[26] = IN1[30]&IN2[2];
  assign P33[25] = IN1[30]&IN2[3];
  assign P34[24] = IN1[30]&IN2[4];
  assign P35[23] = IN1[30]&IN2[5];
  assign P36[22] = IN1[30]&IN2[6];
  assign P37[21] = IN1[30]&IN2[7];
  assign P38[20] = IN1[30]&IN2[8];
  assign P39[19] = IN1[30]&IN2[9];
  assign P40[18] = IN1[30]&IN2[10];
  assign P41[17] = IN1[30]&IN2[11];
  assign P42[16] = IN1[30]&IN2[12];
  assign P43[15] = IN1[30]&IN2[13];
  assign P44[14] = IN1[30]&IN2[14];
  assign P45[13] = IN1[30]&IN2[15];
  assign P46[12] = IN1[30]&IN2[16];
  assign P47[11] = IN1[30]&IN2[17];
  assign P48[10] = IN1[30]&IN2[18];
  assign P49[9] = IN1[30]&IN2[19];
  assign P50[8] = IN1[30]&IN2[20];
  assign P51[7] = IN1[30]&IN2[21];
  assign P52[6] = IN1[30]&IN2[22];
  assign P53[5] = IN1[30]&IN2[23];
  assign P54[4] = IN1[30]&IN2[24];
  assign P55[3] = IN1[30]&IN2[25];
  assign P56[2] = IN1[30]&IN2[26];
  assign P57[1] = IN1[30]&IN2[27];
  assign P58[0] = IN1[30]&IN2[28];
  assign P31[28] = IN1[31]&IN2[0];
  assign P32[27] = IN1[31]&IN2[1];
  assign P33[26] = IN1[31]&IN2[2];
  assign P34[25] = IN1[31]&IN2[3];
  assign P35[24] = IN1[31]&IN2[4];
  assign P36[23] = IN1[31]&IN2[5];
  assign P37[22] = IN1[31]&IN2[6];
  assign P38[21] = IN1[31]&IN2[7];
  assign P39[20] = IN1[31]&IN2[8];
  assign P40[19] = IN1[31]&IN2[9];
  assign P41[18] = IN1[31]&IN2[10];
  assign P42[17] = IN1[31]&IN2[11];
  assign P43[16] = IN1[31]&IN2[12];
  assign P44[15] = IN1[31]&IN2[13];
  assign P45[14] = IN1[31]&IN2[14];
  assign P46[13] = IN1[31]&IN2[15];
  assign P47[12] = IN1[31]&IN2[16];
  assign P48[11] = IN1[31]&IN2[17];
  assign P49[10] = IN1[31]&IN2[18];
  assign P50[9] = IN1[31]&IN2[19];
  assign P51[8] = IN1[31]&IN2[20];
  assign P52[7] = IN1[31]&IN2[21];
  assign P53[6] = IN1[31]&IN2[22];
  assign P54[5] = IN1[31]&IN2[23];
  assign P55[4] = IN1[31]&IN2[24];
  assign P56[3] = IN1[31]&IN2[25];
  assign P57[2] = IN1[31]&IN2[26];
  assign P58[1] = IN1[31]&IN2[27];
  assign P59[0] = IN1[31]&IN2[28];
  assign P32[28] = IN1[32]&IN2[0];
  assign P33[27] = IN1[32]&IN2[1];
  assign P34[26] = IN1[32]&IN2[2];
  assign P35[25] = IN1[32]&IN2[3];
  assign P36[24] = IN1[32]&IN2[4];
  assign P37[23] = IN1[32]&IN2[5];
  assign P38[22] = IN1[32]&IN2[6];
  assign P39[21] = IN1[32]&IN2[7];
  assign P40[20] = IN1[32]&IN2[8];
  assign P41[19] = IN1[32]&IN2[9];
  assign P42[18] = IN1[32]&IN2[10];
  assign P43[17] = IN1[32]&IN2[11];
  assign P44[16] = IN1[32]&IN2[12];
  assign P45[15] = IN1[32]&IN2[13];
  assign P46[14] = IN1[32]&IN2[14];
  assign P47[13] = IN1[32]&IN2[15];
  assign P48[12] = IN1[32]&IN2[16];
  assign P49[11] = IN1[32]&IN2[17];
  assign P50[10] = IN1[32]&IN2[18];
  assign P51[9] = IN1[32]&IN2[19];
  assign P52[8] = IN1[32]&IN2[20];
  assign P53[7] = IN1[32]&IN2[21];
  assign P54[6] = IN1[32]&IN2[22];
  assign P55[5] = IN1[32]&IN2[23];
  assign P56[4] = IN1[32]&IN2[24];
  assign P57[3] = IN1[32]&IN2[25];
  assign P58[2] = IN1[32]&IN2[26];
  assign P59[1] = IN1[32]&IN2[27];
  assign P60[0] = IN1[32]&IN2[28];
  assign P33[28] = IN1[33]&IN2[0];
  assign P34[27] = IN1[33]&IN2[1];
  assign P35[26] = IN1[33]&IN2[2];
  assign P36[25] = IN1[33]&IN2[3];
  assign P37[24] = IN1[33]&IN2[4];
  assign P38[23] = IN1[33]&IN2[5];
  assign P39[22] = IN1[33]&IN2[6];
  assign P40[21] = IN1[33]&IN2[7];
  assign P41[20] = IN1[33]&IN2[8];
  assign P42[19] = IN1[33]&IN2[9];
  assign P43[18] = IN1[33]&IN2[10];
  assign P44[17] = IN1[33]&IN2[11];
  assign P45[16] = IN1[33]&IN2[12];
  assign P46[15] = IN1[33]&IN2[13];
  assign P47[14] = IN1[33]&IN2[14];
  assign P48[13] = IN1[33]&IN2[15];
  assign P49[12] = IN1[33]&IN2[16];
  assign P50[11] = IN1[33]&IN2[17];
  assign P51[10] = IN1[33]&IN2[18];
  assign P52[9] = IN1[33]&IN2[19];
  assign P53[8] = IN1[33]&IN2[20];
  assign P54[7] = IN1[33]&IN2[21];
  assign P55[6] = IN1[33]&IN2[22];
  assign P56[5] = IN1[33]&IN2[23];
  assign P57[4] = IN1[33]&IN2[24];
  assign P58[3] = IN1[33]&IN2[25];
  assign P59[2] = IN1[33]&IN2[26];
  assign P60[1] = IN1[33]&IN2[27];
  assign P61[0] = IN1[33]&IN2[28];
  assign P34[28] = IN1[34]&IN2[0];
  assign P35[27] = IN1[34]&IN2[1];
  assign P36[26] = IN1[34]&IN2[2];
  assign P37[25] = IN1[34]&IN2[3];
  assign P38[24] = IN1[34]&IN2[4];
  assign P39[23] = IN1[34]&IN2[5];
  assign P40[22] = IN1[34]&IN2[6];
  assign P41[21] = IN1[34]&IN2[7];
  assign P42[20] = IN1[34]&IN2[8];
  assign P43[19] = IN1[34]&IN2[9];
  assign P44[18] = IN1[34]&IN2[10];
  assign P45[17] = IN1[34]&IN2[11];
  assign P46[16] = IN1[34]&IN2[12];
  assign P47[15] = IN1[34]&IN2[13];
  assign P48[14] = IN1[34]&IN2[14];
  assign P49[13] = IN1[34]&IN2[15];
  assign P50[12] = IN1[34]&IN2[16];
  assign P51[11] = IN1[34]&IN2[17];
  assign P52[10] = IN1[34]&IN2[18];
  assign P53[9] = IN1[34]&IN2[19];
  assign P54[8] = IN1[34]&IN2[20];
  assign P55[7] = IN1[34]&IN2[21];
  assign P56[6] = IN1[34]&IN2[22];
  assign P57[5] = IN1[34]&IN2[23];
  assign P58[4] = IN1[34]&IN2[24];
  assign P59[3] = IN1[34]&IN2[25];
  assign P60[2] = IN1[34]&IN2[26];
  assign P61[1] = IN1[34]&IN2[27];
  assign P62[0] = IN1[34]&IN2[28];
  assign P35[28] = IN1[35]&IN2[0];
  assign P36[27] = IN1[35]&IN2[1];
  assign P37[26] = IN1[35]&IN2[2];
  assign P38[25] = IN1[35]&IN2[3];
  assign P39[24] = IN1[35]&IN2[4];
  assign P40[23] = IN1[35]&IN2[5];
  assign P41[22] = IN1[35]&IN2[6];
  assign P42[21] = IN1[35]&IN2[7];
  assign P43[20] = IN1[35]&IN2[8];
  assign P44[19] = IN1[35]&IN2[9];
  assign P45[18] = IN1[35]&IN2[10];
  assign P46[17] = IN1[35]&IN2[11];
  assign P47[16] = IN1[35]&IN2[12];
  assign P48[15] = IN1[35]&IN2[13];
  assign P49[14] = IN1[35]&IN2[14];
  assign P50[13] = IN1[35]&IN2[15];
  assign P51[12] = IN1[35]&IN2[16];
  assign P52[11] = IN1[35]&IN2[17];
  assign P53[10] = IN1[35]&IN2[18];
  assign P54[9] = IN1[35]&IN2[19];
  assign P55[8] = IN1[35]&IN2[20];
  assign P56[7] = IN1[35]&IN2[21];
  assign P57[6] = IN1[35]&IN2[22];
  assign P58[5] = IN1[35]&IN2[23];
  assign P59[4] = IN1[35]&IN2[24];
  assign P60[3] = IN1[35]&IN2[25];
  assign P61[2] = IN1[35]&IN2[26];
  assign P62[1] = IN1[35]&IN2[27];
  assign P63[0] = IN1[35]&IN2[28];
  assign P36[28] = IN1[36]&IN2[0];
  assign P37[27] = IN1[36]&IN2[1];
  assign P38[26] = IN1[36]&IN2[2];
  assign P39[25] = IN1[36]&IN2[3];
  assign P40[24] = IN1[36]&IN2[4];
  assign P41[23] = IN1[36]&IN2[5];
  assign P42[22] = IN1[36]&IN2[6];
  assign P43[21] = IN1[36]&IN2[7];
  assign P44[20] = IN1[36]&IN2[8];
  assign P45[19] = IN1[36]&IN2[9];
  assign P46[18] = IN1[36]&IN2[10];
  assign P47[17] = IN1[36]&IN2[11];
  assign P48[16] = IN1[36]&IN2[12];
  assign P49[15] = IN1[36]&IN2[13];
  assign P50[14] = IN1[36]&IN2[14];
  assign P51[13] = IN1[36]&IN2[15];
  assign P52[12] = IN1[36]&IN2[16];
  assign P53[11] = IN1[36]&IN2[17];
  assign P54[10] = IN1[36]&IN2[18];
  assign P55[9] = IN1[36]&IN2[19];
  assign P56[8] = IN1[36]&IN2[20];
  assign P57[7] = IN1[36]&IN2[21];
  assign P58[6] = IN1[36]&IN2[22];
  assign P59[5] = IN1[36]&IN2[23];
  assign P60[4] = IN1[36]&IN2[24];
  assign P61[3] = IN1[36]&IN2[25];
  assign P62[2] = IN1[36]&IN2[26];
  assign P63[1] = IN1[36]&IN2[27];
  assign P64[0] = IN1[36]&IN2[28];
  assign P37[28] = IN1[37]&IN2[0];
  assign P38[27] = IN1[37]&IN2[1];
  assign P39[26] = IN1[37]&IN2[2];
  assign P40[25] = IN1[37]&IN2[3];
  assign P41[24] = IN1[37]&IN2[4];
  assign P42[23] = IN1[37]&IN2[5];
  assign P43[22] = IN1[37]&IN2[6];
  assign P44[21] = IN1[37]&IN2[7];
  assign P45[20] = IN1[37]&IN2[8];
  assign P46[19] = IN1[37]&IN2[9];
  assign P47[18] = IN1[37]&IN2[10];
  assign P48[17] = IN1[37]&IN2[11];
  assign P49[16] = IN1[37]&IN2[12];
  assign P50[15] = IN1[37]&IN2[13];
  assign P51[14] = IN1[37]&IN2[14];
  assign P52[13] = IN1[37]&IN2[15];
  assign P53[12] = IN1[37]&IN2[16];
  assign P54[11] = IN1[37]&IN2[17];
  assign P55[10] = IN1[37]&IN2[18];
  assign P56[9] = IN1[37]&IN2[19];
  assign P57[8] = IN1[37]&IN2[20];
  assign P58[7] = IN1[37]&IN2[21];
  assign P59[6] = IN1[37]&IN2[22];
  assign P60[5] = IN1[37]&IN2[23];
  assign P61[4] = IN1[37]&IN2[24];
  assign P62[3] = IN1[37]&IN2[25];
  assign P63[2] = IN1[37]&IN2[26];
  assign P64[1] = IN1[37]&IN2[27];
  assign P65[0] = IN1[37]&IN2[28];
  assign P38[28] = IN1[38]&IN2[0];
  assign P39[27] = IN1[38]&IN2[1];
  assign P40[26] = IN1[38]&IN2[2];
  assign P41[25] = IN1[38]&IN2[3];
  assign P42[24] = IN1[38]&IN2[4];
  assign P43[23] = IN1[38]&IN2[5];
  assign P44[22] = IN1[38]&IN2[6];
  assign P45[21] = IN1[38]&IN2[7];
  assign P46[20] = IN1[38]&IN2[8];
  assign P47[19] = IN1[38]&IN2[9];
  assign P48[18] = IN1[38]&IN2[10];
  assign P49[17] = IN1[38]&IN2[11];
  assign P50[16] = IN1[38]&IN2[12];
  assign P51[15] = IN1[38]&IN2[13];
  assign P52[14] = IN1[38]&IN2[14];
  assign P53[13] = IN1[38]&IN2[15];
  assign P54[12] = IN1[38]&IN2[16];
  assign P55[11] = IN1[38]&IN2[17];
  assign P56[10] = IN1[38]&IN2[18];
  assign P57[9] = IN1[38]&IN2[19];
  assign P58[8] = IN1[38]&IN2[20];
  assign P59[7] = IN1[38]&IN2[21];
  assign P60[6] = IN1[38]&IN2[22];
  assign P61[5] = IN1[38]&IN2[23];
  assign P62[4] = IN1[38]&IN2[24];
  assign P63[3] = IN1[38]&IN2[25];
  assign P64[2] = IN1[38]&IN2[26];
  assign P65[1] = IN1[38]&IN2[27];
  assign P66[0] = IN1[38]&IN2[28];
  assign P39[28] = IN1[39]&IN2[0];
  assign P40[27] = IN1[39]&IN2[1];
  assign P41[26] = IN1[39]&IN2[2];
  assign P42[25] = IN1[39]&IN2[3];
  assign P43[24] = IN1[39]&IN2[4];
  assign P44[23] = IN1[39]&IN2[5];
  assign P45[22] = IN1[39]&IN2[6];
  assign P46[21] = IN1[39]&IN2[7];
  assign P47[20] = IN1[39]&IN2[8];
  assign P48[19] = IN1[39]&IN2[9];
  assign P49[18] = IN1[39]&IN2[10];
  assign P50[17] = IN1[39]&IN2[11];
  assign P51[16] = IN1[39]&IN2[12];
  assign P52[15] = IN1[39]&IN2[13];
  assign P53[14] = IN1[39]&IN2[14];
  assign P54[13] = IN1[39]&IN2[15];
  assign P55[12] = IN1[39]&IN2[16];
  assign P56[11] = IN1[39]&IN2[17];
  assign P57[10] = IN1[39]&IN2[18];
  assign P58[9] = IN1[39]&IN2[19];
  assign P59[8] = IN1[39]&IN2[20];
  assign P60[7] = IN1[39]&IN2[21];
  assign P61[6] = IN1[39]&IN2[22];
  assign P62[5] = IN1[39]&IN2[23];
  assign P63[4] = IN1[39]&IN2[24];
  assign P64[3] = IN1[39]&IN2[25];
  assign P65[2] = IN1[39]&IN2[26];
  assign P66[1] = IN1[39]&IN2[27];
  assign P67[0] = IN1[39]&IN2[28];
  assign P40[28] = IN1[40]&IN2[0];
  assign P41[27] = IN1[40]&IN2[1];
  assign P42[26] = IN1[40]&IN2[2];
  assign P43[25] = IN1[40]&IN2[3];
  assign P44[24] = IN1[40]&IN2[4];
  assign P45[23] = IN1[40]&IN2[5];
  assign P46[22] = IN1[40]&IN2[6];
  assign P47[21] = IN1[40]&IN2[7];
  assign P48[20] = IN1[40]&IN2[8];
  assign P49[19] = IN1[40]&IN2[9];
  assign P50[18] = IN1[40]&IN2[10];
  assign P51[17] = IN1[40]&IN2[11];
  assign P52[16] = IN1[40]&IN2[12];
  assign P53[15] = IN1[40]&IN2[13];
  assign P54[14] = IN1[40]&IN2[14];
  assign P55[13] = IN1[40]&IN2[15];
  assign P56[12] = IN1[40]&IN2[16];
  assign P57[11] = IN1[40]&IN2[17];
  assign P58[10] = IN1[40]&IN2[18];
  assign P59[9] = IN1[40]&IN2[19];
  assign P60[8] = IN1[40]&IN2[20];
  assign P61[7] = IN1[40]&IN2[21];
  assign P62[6] = IN1[40]&IN2[22];
  assign P63[5] = IN1[40]&IN2[23];
  assign P64[4] = IN1[40]&IN2[24];
  assign P65[3] = IN1[40]&IN2[25];
  assign P66[2] = IN1[40]&IN2[26];
  assign P67[1] = IN1[40]&IN2[27];
  assign P68[0] = IN1[40]&IN2[28];
  assign P41[28] = IN1[41]&IN2[0];
  assign P42[27] = IN1[41]&IN2[1];
  assign P43[26] = IN1[41]&IN2[2];
  assign P44[25] = IN1[41]&IN2[3];
  assign P45[24] = IN1[41]&IN2[4];
  assign P46[23] = IN1[41]&IN2[5];
  assign P47[22] = IN1[41]&IN2[6];
  assign P48[21] = IN1[41]&IN2[7];
  assign P49[20] = IN1[41]&IN2[8];
  assign P50[19] = IN1[41]&IN2[9];
  assign P51[18] = IN1[41]&IN2[10];
  assign P52[17] = IN1[41]&IN2[11];
  assign P53[16] = IN1[41]&IN2[12];
  assign P54[15] = IN1[41]&IN2[13];
  assign P55[14] = IN1[41]&IN2[14];
  assign P56[13] = IN1[41]&IN2[15];
  assign P57[12] = IN1[41]&IN2[16];
  assign P58[11] = IN1[41]&IN2[17];
  assign P59[10] = IN1[41]&IN2[18];
  assign P60[9] = IN1[41]&IN2[19];
  assign P61[8] = IN1[41]&IN2[20];
  assign P62[7] = IN1[41]&IN2[21];
  assign P63[6] = IN1[41]&IN2[22];
  assign P64[5] = IN1[41]&IN2[23];
  assign P65[4] = IN1[41]&IN2[24];
  assign P66[3] = IN1[41]&IN2[25];
  assign P67[2] = IN1[41]&IN2[26];
  assign P68[1] = IN1[41]&IN2[27];
  assign P69[0] = IN1[41]&IN2[28];
  assign P42[28] = IN1[42]&IN2[0];
  assign P43[27] = IN1[42]&IN2[1];
  assign P44[26] = IN1[42]&IN2[2];
  assign P45[25] = IN1[42]&IN2[3];
  assign P46[24] = IN1[42]&IN2[4];
  assign P47[23] = IN1[42]&IN2[5];
  assign P48[22] = IN1[42]&IN2[6];
  assign P49[21] = IN1[42]&IN2[7];
  assign P50[20] = IN1[42]&IN2[8];
  assign P51[19] = IN1[42]&IN2[9];
  assign P52[18] = IN1[42]&IN2[10];
  assign P53[17] = IN1[42]&IN2[11];
  assign P54[16] = IN1[42]&IN2[12];
  assign P55[15] = IN1[42]&IN2[13];
  assign P56[14] = IN1[42]&IN2[14];
  assign P57[13] = IN1[42]&IN2[15];
  assign P58[12] = IN1[42]&IN2[16];
  assign P59[11] = IN1[42]&IN2[17];
  assign P60[10] = IN1[42]&IN2[18];
  assign P61[9] = IN1[42]&IN2[19];
  assign P62[8] = IN1[42]&IN2[20];
  assign P63[7] = IN1[42]&IN2[21];
  assign P64[6] = IN1[42]&IN2[22];
  assign P65[5] = IN1[42]&IN2[23];
  assign P66[4] = IN1[42]&IN2[24];
  assign P67[3] = IN1[42]&IN2[25];
  assign P68[2] = IN1[42]&IN2[26];
  assign P69[1] = IN1[42]&IN2[27];
  assign P70[0] = IN1[42]&IN2[28];
  assign P43[28] = IN1[43]&IN2[0];
  assign P44[27] = IN1[43]&IN2[1];
  assign P45[26] = IN1[43]&IN2[2];
  assign P46[25] = IN1[43]&IN2[3];
  assign P47[24] = IN1[43]&IN2[4];
  assign P48[23] = IN1[43]&IN2[5];
  assign P49[22] = IN1[43]&IN2[6];
  assign P50[21] = IN1[43]&IN2[7];
  assign P51[20] = IN1[43]&IN2[8];
  assign P52[19] = IN1[43]&IN2[9];
  assign P53[18] = IN1[43]&IN2[10];
  assign P54[17] = IN1[43]&IN2[11];
  assign P55[16] = IN1[43]&IN2[12];
  assign P56[15] = IN1[43]&IN2[13];
  assign P57[14] = IN1[43]&IN2[14];
  assign P58[13] = IN1[43]&IN2[15];
  assign P59[12] = IN1[43]&IN2[16];
  assign P60[11] = IN1[43]&IN2[17];
  assign P61[10] = IN1[43]&IN2[18];
  assign P62[9] = IN1[43]&IN2[19];
  assign P63[8] = IN1[43]&IN2[20];
  assign P64[7] = IN1[43]&IN2[21];
  assign P65[6] = IN1[43]&IN2[22];
  assign P66[5] = IN1[43]&IN2[23];
  assign P67[4] = IN1[43]&IN2[24];
  assign P68[3] = IN1[43]&IN2[25];
  assign P69[2] = IN1[43]&IN2[26];
  assign P70[1] = IN1[43]&IN2[27];
  assign P71[0] = IN1[43]&IN2[28];
  assign P44[28] = IN1[44]&IN2[0];
  assign P45[27] = IN1[44]&IN2[1];
  assign P46[26] = IN1[44]&IN2[2];
  assign P47[25] = IN1[44]&IN2[3];
  assign P48[24] = IN1[44]&IN2[4];
  assign P49[23] = IN1[44]&IN2[5];
  assign P50[22] = IN1[44]&IN2[6];
  assign P51[21] = IN1[44]&IN2[7];
  assign P52[20] = IN1[44]&IN2[8];
  assign P53[19] = IN1[44]&IN2[9];
  assign P54[18] = IN1[44]&IN2[10];
  assign P55[17] = IN1[44]&IN2[11];
  assign P56[16] = IN1[44]&IN2[12];
  assign P57[15] = IN1[44]&IN2[13];
  assign P58[14] = IN1[44]&IN2[14];
  assign P59[13] = IN1[44]&IN2[15];
  assign P60[12] = IN1[44]&IN2[16];
  assign P61[11] = IN1[44]&IN2[17];
  assign P62[10] = IN1[44]&IN2[18];
  assign P63[9] = IN1[44]&IN2[19];
  assign P64[8] = IN1[44]&IN2[20];
  assign P65[7] = IN1[44]&IN2[21];
  assign P66[6] = IN1[44]&IN2[22];
  assign P67[5] = IN1[44]&IN2[23];
  assign P68[4] = IN1[44]&IN2[24];
  assign P69[3] = IN1[44]&IN2[25];
  assign P70[2] = IN1[44]&IN2[26];
  assign P71[1] = IN1[44]&IN2[27];
  assign P72[0] = IN1[44]&IN2[28];
  assign P45[28] = IN1[45]&IN2[0];
  assign P46[27] = IN1[45]&IN2[1];
  assign P47[26] = IN1[45]&IN2[2];
  assign P48[25] = IN1[45]&IN2[3];
  assign P49[24] = IN1[45]&IN2[4];
  assign P50[23] = IN1[45]&IN2[5];
  assign P51[22] = IN1[45]&IN2[6];
  assign P52[21] = IN1[45]&IN2[7];
  assign P53[20] = IN1[45]&IN2[8];
  assign P54[19] = IN1[45]&IN2[9];
  assign P55[18] = IN1[45]&IN2[10];
  assign P56[17] = IN1[45]&IN2[11];
  assign P57[16] = IN1[45]&IN2[12];
  assign P58[15] = IN1[45]&IN2[13];
  assign P59[14] = IN1[45]&IN2[14];
  assign P60[13] = IN1[45]&IN2[15];
  assign P61[12] = IN1[45]&IN2[16];
  assign P62[11] = IN1[45]&IN2[17];
  assign P63[10] = IN1[45]&IN2[18];
  assign P64[9] = IN1[45]&IN2[19];
  assign P65[8] = IN1[45]&IN2[20];
  assign P66[7] = IN1[45]&IN2[21];
  assign P67[6] = IN1[45]&IN2[22];
  assign P68[5] = IN1[45]&IN2[23];
  assign P69[4] = IN1[45]&IN2[24];
  assign P70[3] = IN1[45]&IN2[25];
  assign P71[2] = IN1[45]&IN2[26];
  assign P72[1] = IN1[45]&IN2[27];
  assign P73[0] = IN1[45]&IN2[28];
  assign P46[28] = IN1[46]&IN2[0];
  assign P47[27] = IN1[46]&IN2[1];
  assign P48[26] = IN1[46]&IN2[2];
  assign P49[25] = IN1[46]&IN2[3];
  assign P50[24] = IN1[46]&IN2[4];
  assign P51[23] = IN1[46]&IN2[5];
  assign P52[22] = IN1[46]&IN2[6];
  assign P53[21] = IN1[46]&IN2[7];
  assign P54[20] = IN1[46]&IN2[8];
  assign P55[19] = IN1[46]&IN2[9];
  assign P56[18] = IN1[46]&IN2[10];
  assign P57[17] = IN1[46]&IN2[11];
  assign P58[16] = IN1[46]&IN2[12];
  assign P59[15] = IN1[46]&IN2[13];
  assign P60[14] = IN1[46]&IN2[14];
  assign P61[13] = IN1[46]&IN2[15];
  assign P62[12] = IN1[46]&IN2[16];
  assign P63[11] = IN1[46]&IN2[17];
  assign P64[10] = IN1[46]&IN2[18];
  assign P65[9] = IN1[46]&IN2[19];
  assign P66[8] = IN1[46]&IN2[20];
  assign P67[7] = IN1[46]&IN2[21];
  assign P68[6] = IN1[46]&IN2[22];
  assign P69[5] = IN1[46]&IN2[23];
  assign P70[4] = IN1[46]&IN2[24];
  assign P71[3] = IN1[46]&IN2[25];
  assign P72[2] = IN1[46]&IN2[26];
  assign P73[1] = IN1[46]&IN2[27];
  assign P74[0] = IN1[46]&IN2[28];
  assign P47[28] = IN1[47]&IN2[0];
  assign P48[27] = IN1[47]&IN2[1];
  assign P49[26] = IN1[47]&IN2[2];
  assign P50[25] = IN1[47]&IN2[3];
  assign P51[24] = IN1[47]&IN2[4];
  assign P52[23] = IN1[47]&IN2[5];
  assign P53[22] = IN1[47]&IN2[6];
  assign P54[21] = IN1[47]&IN2[7];
  assign P55[20] = IN1[47]&IN2[8];
  assign P56[19] = IN1[47]&IN2[9];
  assign P57[18] = IN1[47]&IN2[10];
  assign P58[17] = IN1[47]&IN2[11];
  assign P59[16] = IN1[47]&IN2[12];
  assign P60[15] = IN1[47]&IN2[13];
  assign P61[14] = IN1[47]&IN2[14];
  assign P62[13] = IN1[47]&IN2[15];
  assign P63[12] = IN1[47]&IN2[16];
  assign P64[11] = IN1[47]&IN2[17];
  assign P65[10] = IN1[47]&IN2[18];
  assign P66[9] = IN1[47]&IN2[19];
  assign P67[8] = IN1[47]&IN2[20];
  assign P68[7] = IN1[47]&IN2[21];
  assign P69[6] = IN1[47]&IN2[22];
  assign P70[5] = IN1[47]&IN2[23];
  assign P71[4] = IN1[47]&IN2[24];
  assign P72[3] = IN1[47]&IN2[25];
  assign P73[2] = IN1[47]&IN2[26];
  assign P74[1] = IN1[47]&IN2[27];
  assign P75[0] = IN1[47]&IN2[28];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [28:0] IN29;
  input [28:0] IN30;
  input [28:0] IN31;
  input [28:0] IN32;
  input [28:0] IN33;
  input [28:0] IN34;
  input [28:0] IN35;
  input [28:0] IN36;
  input [28:0] IN37;
  input [28:0] IN38;
  input [28:0] IN39;
  input [28:0] IN40;
  input [28:0] IN41;
  input [28:0] IN42;
  input [28:0] IN43;
  input [28:0] IN44;
  input [28:0] IN45;
  input [28:0] IN46;
  input [28:0] IN47;
  input [27:0] IN48;
  input [26:0] IN49;
  input [25:0] IN50;
  input [24:0] IN51;
  input [23:0] IN52;
  input [22:0] IN53;
  input [21:0] IN54;
  input [20:0] IN55;
  input [19:0] IN56;
  input [18:0] IN57;
  input [17:0] IN58;
  input [16:0] IN59;
  input [15:0] IN60;
  input [14:0] IN61;
  input [13:0] IN62;
  input [12:0] IN63;
  input [11:0] IN64;
  input [10:0] IN65;
  input [9:0] IN66;
  input [8:0] IN67;
  input [7:0] IN68;
  input [6:0] IN69;
  input [5:0] IN70;
  input [4:0] IN71;
  input [3:0] IN72;
  input [2:0] IN73;
  input [1:0] IN74;
  input [0:0] IN75;
  output [75:0] Out1;
  output [27:0] Out2;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1984;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2088;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2140;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2585;
  wire w2586;
  wire w2587;
  wire w2588;
  wire w2589;
  wire w2590;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2631;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2638;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2680;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2685;
  wire w2686;
  wire w2687;
  wire w2688;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2694;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2738;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2747;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2770;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2774;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2785;
  wire w2786;
  wire w2787;
  wire w2788;
  wire w2789;
  wire w2790;
  wire w2791;
  wire w2792;
  wire w2793;
  wire w2794;
  wire w2795;
  wire w2796;
  wire w2797;
  wire w2798;
  wire w2799;
  wire w2800;
  wire w2801;
  wire w2803;
  wire w2804;
  wire w2805;
  wire w2806;
  wire w2807;
  wire w2808;
  wire w2809;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2854;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2860;
  wire w2861;
  wire w2862;
  wire w2863;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2885;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2913;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2934;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2950;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2979;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2985;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3014;
  wire w3015;
  wire w3016;
  wire w3017;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3040;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3085;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3094;
  wire w3095;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3121;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3130;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3225;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3254;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3262;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3285;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3327;
  wire w3328;
  wire w3329;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3334;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3362;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3385;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3414;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3433;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3443;
  wire w3444;
  wire w3445;
  wire w3446;
  wire w3447;
  wire w3448;
  wire w3449;
  wire w3450;
  wire w3451;
  wire w3452;
  wire w3453;
  wire w3454;
  wire w3455;
  wire w3456;
  wire w3457;
  wire w3458;
  wire w3459;
  wire w3461;
  wire w3462;
  wire w3463;
  wire w3464;
  wire w3465;
  wire w3466;
  wire w3467;
  wire w3468;
  wire w3469;
  wire w3470;
  wire w3471;
  wire w3472;
  wire w3473;
  wire w3474;
  wire w3475;
  wire w3476;
  wire w3477;
  wire w3478;
  wire w3479;
  wire w3480;
  wire w3481;
  wire w3482;
  wire w3483;
  wire w3484;
  wire w3485;
  wire w3486;
  wire w3487;
  wire w3488;
  wire w3489;
  wire w3490;
  wire w3491;
  wire w3492;
  wire w3493;
  wire w3494;
  wire w3495;
  wire w3496;
  wire w3497;
  wire w3498;
  wire w3499;
  wire w3500;
  wire w3501;
  wire w3502;
  wire w3503;
  wire w3504;
  wire w3505;
  wire w3506;
  wire w3507;
  wire w3508;
  wire w3509;
  wire w3510;
  wire w3511;
  wire w3512;
  wire w3513;
  wire w3514;
  wire w3515;
  wire w3516;
  wire w3517;
  wire w3518;
  wire w3519;
  wire w3520;
  wire w3521;
  wire w3522;
  wire w3523;
  wire w3524;
  wire w3525;
  wire w3526;
  wire w3527;
  wire w3528;
  wire w3529;
  wire w3530;
  wire w3531;
  wire w3532;
  wire w3533;
  wire w3534;
  wire w3535;
  wire w3536;
  wire w3537;
  wire w3538;
  wire w3539;
  wire w3540;
  wire w3541;
  wire w3542;
  wire w3543;
  wire w3544;
  wire w3545;
  wire w3546;
  wire w3547;
  wire w3548;
  wire w3549;
  wire w3550;
  wire w3551;
  wire w3552;
  wire w3553;
  wire w3555;
  wire w3556;
  wire w3557;
  wire w3558;
  wire w3559;
  wire w3560;
  wire w3561;
  wire w3562;
  wire w3563;
  wire w3564;
  wire w3565;
  wire w3566;
  wire w3567;
  wire w3568;
  wire w3569;
  wire w3570;
  wire w3571;
  wire w3572;
  wire w3573;
  wire w3574;
  wire w3575;
  wire w3576;
  wire w3577;
  wire w3578;
  wire w3579;
  wire w3580;
  wire w3581;
  wire w3582;
  wire w3583;
  wire w3584;
  wire w3585;
  wire w3586;
  wire w3587;
  wire w3588;
  wire w3589;
  wire w3590;
  wire w3591;
  wire w3592;
  wire w3593;
  wire w3594;
  wire w3595;
  wire w3596;
  wire w3597;
  wire w3598;
  wire w3599;
  wire w3600;
  wire w3601;
  wire w3602;
  wire w3603;
  wire w3604;
  wire w3605;
  wire w3606;
  wire w3607;
  wire w3608;
  wire w3609;
  wire w3610;
  wire w3611;
  wire w3612;
  wire w3613;
  wire w3614;
  wire w3615;
  wire w3616;
  wire w3617;
  wire w3618;
  wire w3619;
  wire w3620;
  wire w3621;
  wire w3622;
  wire w3623;
  wire w3624;
  wire w3625;
  wire w3626;
  wire w3627;
  wire w3628;
  wire w3629;
  wire w3630;
  wire w3631;
  wire w3632;
  wire w3633;
  wire w3634;
  wire w3635;
  wire w3636;
  wire w3637;
  wire w3638;
  wire w3639;
  wire w3640;
  wire w3641;
  wire w3642;
  wire w3643;
  wire w3644;
  wire w3645;
  wire w3646;
  wire w3647;
  wire w3649;
  wire w3650;
  wire w3651;
  wire w3652;
  wire w3653;
  wire w3654;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3662;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3685;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3734;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3743;
  wire w3744;
  wire w3745;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3762;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3768;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3785;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3814;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3849;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3862;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3882;
  wire w3883;
  wire w3884;
  wire w3885;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3894;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3931;
  wire w3933;
  wire w3935;
  wire w3937;
  wire w3939;
  wire w3941;
  wire w3943;
  wire w3945;
  wire w3947;
  wire w3949;
  wire w3951;
  wire w3953;
  wire w3955;
  wire w3957;
  wire w3959;
  wire w3961;
  wire w3963;
  wire w3965;
  wire w3967;
  wire w3969;
  wire w3971;
  wire w3973;
  wire w3975;
  wire w3977;
  wire w3979;
  wire w3981;
  wire w3983;
  wire w3985;
  wire w3987;
  wire w3989;
  wire w3991;
  wire w3993;
  wire w3995;
  wire w3997;
  wire w3999;
  wire w4001;
  wire w4003;
  wire w4005;
  wire w4007;
  wire w4009;
  wire w4011;
  wire w4013;
  wire w4015;
  wire w4017;
  wire w4019;
  wire w4021;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w1393);
  FullAdder U1 (w1393, IN2[0], IN2[1], w1394, w1395);
  FullAdder U2 (w1395, IN3[0], IN3[1], w1396, w1397);
  FullAdder U3 (w1397, IN4[0], IN4[1], w1398, w1399);
  FullAdder U4 (w1399, IN5[0], IN5[1], w1400, w1401);
  FullAdder U5 (w1401, IN6[0], IN6[1], w1402, w1403);
  FullAdder U6 (w1403, IN7[0], IN7[1], w1404, w1405);
  FullAdder U7 (w1405, IN8[0], IN8[1], w1406, w1407);
  FullAdder U8 (w1407, IN9[0], IN9[1], w1408, w1409);
  FullAdder U9 (w1409, IN10[0], IN10[1], w1410, w1411);
  FullAdder U10 (w1411, IN11[0], IN11[1], w1412, w1413);
  FullAdder U11 (w1413, IN12[0], IN12[1], w1414, w1415);
  FullAdder U12 (w1415, IN13[0], IN13[1], w1416, w1417);
  FullAdder U13 (w1417, IN14[0], IN14[1], w1418, w1419);
  FullAdder U14 (w1419, IN15[0], IN15[1], w1420, w1421);
  FullAdder U15 (w1421, IN16[0], IN16[1], w1422, w1423);
  FullAdder U16 (w1423, IN17[0], IN17[1], w1424, w1425);
  FullAdder U17 (w1425, IN18[0], IN18[1], w1426, w1427);
  FullAdder U18 (w1427, IN19[0], IN19[1], w1428, w1429);
  FullAdder U19 (w1429, IN20[0], IN20[1], w1430, w1431);
  FullAdder U20 (w1431, IN21[0], IN21[1], w1432, w1433);
  FullAdder U21 (w1433, IN22[0], IN22[1], w1434, w1435);
  FullAdder U22 (w1435, IN23[0], IN23[1], w1436, w1437);
  FullAdder U23 (w1437, IN24[0], IN24[1], w1438, w1439);
  FullAdder U24 (w1439, IN25[0], IN25[1], w1440, w1441);
  FullAdder U25 (w1441, IN26[0], IN26[1], w1442, w1443);
  FullAdder U26 (w1443, IN27[0], IN27[1], w1444, w1445);
  FullAdder U27 (w1445, IN28[0], IN28[1], w1446, w1447);
  FullAdder U28 (w1447, IN29[0], IN29[1], w1448, w1449);
  FullAdder U29 (w1449, IN30[0], IN30[1], w1450, w1451);
  FullAdder U30 (w1451, IN31[0], IN31[1], w1452, w1453);
  FullAdder U31 (w1453, IN32[0], IN32[1], w1454, w1455);
  FullAdder U32 (w1455, IN33[0], IN33[1], w1456, w1457);
  FullAdder U33 (w1457, IN34[0], IN34[1], w1458, w1459);
  FullAdder U34 (w1459, IN35[0], IN35[1], w1460, w1461);
  FullAdder U35 (w1461, IN36[0], IN36[1], w1462, w1463);
  FullAdder U36 (w1463, IN37[0], IN37[1], w1464, w1465);
  FullAdder U37 (w1465, IN38[0], IN38[1], w1466, w1467);
  FullAdder U38 (w1467, IN39[0], IN39[1], w1468, w1469);
  FullAdder U39 (w1469, IN40[0], IN40[1], w1470, w1471);
  FullAdder U40 (w1471, IN41[0], IN41[1], w1472, w1473);
  FullAdder U41 (w1473, IN42[0], IN42[1], w1474, w1475);
  FullAdder U42 (w1475, IN43[0], IN43[1], w1476, w1477);
  FullAdder U43 (w1477, IN44[0], IN44[1], w1478, w1479);
  FullAdder U44 (w1479, IN45[0], IN45[1], w1480, w1481);
  FullAdder U45 (w1481, IN46[0], IN46[1], w1482, w1483);
  FullAdder U46 (w1483, IN47[0], IN47[1], w1484, w1485);
  HalfAdder U47 (w1394, IN2[2], Out1[2], w1487);
  FullAdder U48 (w1487, w1396, IN3[2], w1488, w1489);
  FullAdder U49 (w1489, w1398, IN4[2], w1490, w1491);
  FullAdder U50 (w1491, w1400, IN5[2], w1492, w1493);
  FullAdder U51 (w1493, w1402, IN6[2], w1494, w1495);
  FullAdder U52 (w1495, w1404, IN7[2], w1496, w1497);
  FullAdder U53 (w1497, w1406, IN8[2], w1498, w1499);
  FullAdder U54 (w1499, w1408, IN9[2], w1500, w1501);
  FullAdder U55 (w1501, w1410, IN10[2], w1502, w1503);
  FullAdder U56 (w1503, w1412, IN11[2], w1504, w1505);
  FullAdder U57 (w1505, w1414, IN12[2], w1506, w1507);
  FullAdder U58 (w1507, w1416, IN13[2], w1508, w1509);
  FullAdder U59 (w1509, w1418, IN14[2], w1510, w1511);
  FullAdder U60 (w1511, w1420, IN15[2], w1512, w1513);
  FullAdder U61 (w1513, w1422, IN16[2], w1514, w1515);
  FullAdder U62 (w1515, w1424, IN17[2], w1516, w1517);
  FullAdder U63 (w1517, w1426, IN18[2], w1518, w1519);
  FullAdder U64 (w1519, w1428, IN19[2], w1520, w1521);
  FullAdder U65 (w1521, w1430, IN20[2], w1522, w1523);
  FullAdder U66 (w1523, w1432, IN21[2], w1524, w1525);
  FullAdder U67 (w1525, w1434, IN22[2], w1526, w1527);
  FullAdder U68 (w1527, w1436, IN23[2], w1528, w1529);
  FullAdder U69 (w1529, w1438, IN24[2], w1530, w1531);
  FullAdder U70 (w1531, w1440, IN25[2], w1532, w1533);
  FullAdder U71 (w1533, w1442, IN26[2], w1534, w1535);
  FullAdder U72 (w1535, w1444, IN27[2], w1536, w1537);
  FullAdder U73 (w1537, w1446, IN28[2], w1538, w1539);
  FullAdder U74 (w1539, w1448, IN29[2], w1540, w1541);
  FullAdder U75 (w1541, w1450, IN30[2], w1542, w1543);
  FullAdder U76 (w1543, w1452, IN31[2], w1544, w1545);
  FullAdder U77 (w1545, w1454, IN32[2], w1546, w1547);
  FullAdder U78 (w1547, w1456, IN33[2], w1548, w1549);
  FullAdder U79 (w1549, w1458, IN34[2], w1550, w1551);
  FullAdder U80 (w1551, w1460, IN35[2], w1552, w1553);
  FullAdder U81 (w1553, w1462, IN36[2], w1554, w1555);
  FullAdder U82 (w1555, w1464, IN37[2], w1556, w1557);
  FullAdder U83 (w1557, w1466, IN38[2], w1558, w1559);
  FullAdder U84 (w1559, w1468, IN39[2], w1560, w1561);
  FullAdder U85 (w1561, w1470, IN40[2], w1562, w1563);
  FullAdder U86 (w1563, w1472, IN41[2], w1564, w1565);
  FullAdder U87 (w1565, w1474, IN42[2], w1566, w1567);
  FullAdder U88 (w1567, w1476, IN43[2], w1568, w1569);
  FullAdder U89 (w1569, w1478, IN44[2], w1570, w1571);
  FullAdder U90 (w1571, w1480, IN45[2], w1572, w1573);
  FullAdder U91 (w1573, w1482, IN46[2], w1574, w1575);
  FullAdder U92 (w1575, w1484, IN47[2], w1576, w1577);
  FullAdder U93 (w1577, w1485, IN48[0], w1578, w1579);
  HalfAdder U94 (w1488, IN3[3], Out1[3], w1581);
  FullAdder U95 (w1581, w1490, IN4[3], w1582, w1583);
  FullAdder U96 (w1583, w1492, IN5[3], w1584, w1585);
  FullAdder U97 (w1585, w1494, IN6[3], w1586, w1587);
  FullAdder U98 (w1587, w1496, IN7[3], w1588, w1589);
  FullAdder U99 (w1589, w1498, IN8[3], w1590, w1591);
  FullAdder U100 (w1591, w1500, IN9[3], w1592, w1593);
  FullAdder U101 (w1593, w1502, IN10[3], w1594, w1595);
  FullAdder U102 (w1595, w1504, IN11[3], w1596, w1597);
  FullAdder U103 (w1597, w1506, IN12[3], w1598, w1599);
  FullAdder U104 (w1599, w1508, IN13[3], w1600, w1601);
  FullAdder U105 (w1601, w1510, IN14[3], w1602, w1603);
  FullAdder U106 (w1603, w1512, IN15[3], w1604, w1605);
  FullAdder U107 (w1605, w1514, IN16[3], w1606, w1607);
  FullAdder U108 (w1607, w1516, IN17[3], w1608, w1609);
  FullAdder U109 (w1609, w1518, IN18[3], w1610, w1611);
  FullAdder U110 (w1611, w1520, IN19[3], w1612, w1613);
  FullAdder U111 (w1613, w1522, IN20[3], w1614, w1615);
  FullAdder U112 (w1615, w1524, IN21[3], w1616, w1617);
  FullAdder U113 (w1617, w1526, IN22[3], w1618, w1619);
  FullAdder U114 (w1619, w1528, IN23[3], w1620, w1621);
  FullAdder U115 (w1621, w1530, IN24[3], w1622, w1623);
  FullAdder U116 (w1623, w1532, IN25[3], w1624, w1625);
  FullAdder U117 (w1625, w1534, IN26[3], w1626, w1627);
  FullAdder U118 (w1627, w1536, IN27[3], w1628, w1629);
  FullAdder U119 (w1629, w1538, IN28[3], w1630, w1631);
  FullAdder U120 (w1631, w1540, IN29[3], w1632, w1633);
  FullAdder U121 (w1633, w1542, IN30[3], w1634, w1635);
  FullAdder U122 (w1635, w1544, IN31[3], w1636, w1637);
  FullAdder U123 (w1637, w1546, IN32[3], w1638, w1639);
  FullAdder U124 (w1639, w1548, IN33[3], w1640, w1641);
  FullAdder U125 (w1641, w1550, IN34[3], w1642, w1643);
  FullAdder U126 (w1643, w1552, IN35[3], w1644, w1645);
  FullAdder U127 (w1645, w1554, IN36[3], w1646, w1647);
  FullAdder U128 (w1647, w1556, IN37[3], w1648, w1649);
  FullAdder U129 (w1649, w1558, IN38[3], w1650, w1651);
  FullAdder U130 (w1651, w1560, IN39[3], w1652, w1653);
  FullAdder U131 (w1653, w1562, IN40[3], w1654, w1655);
  FullAdder U132 (w1655, w1564, IN41[3], w1656, w1657);
  FullAdder U133 (w1657, w1566, IN42[3], w1658, w1659);
  FullAdder U134 (w1659, w1568, IN43[3], w1660, w1661);
  FullAdder U135 (w1661, w1570, IN44[3], w1662, w1663);
  FullAdder U136 (w1663, w1572, IN45[3], w1664, w1665);
  FullAdder U137 (w1665, w1574, IN46[3], w1666, w1667);
  FullAdder U138 (w1667, w1576, IN47[3], w1668, w1669);
  FullAdder U139 (w1669, w1578, IN48[1], w1670, w1671);
  FullAdder U140 (w1671, w1579, IN49[0], w1672, w1673);
  HalfAdder U141 (w1582, IN4[4], Out1[4], w1675);
  FullAdder U142 (w1675, w1584, IN5[4], w1676, w1677);
  FullAdder U143 (w1677, w1586, IN6[4], w1678, w1679);
  FullAdder U144 (w1679, w1588, IN7[4], w1680, w1681);
  FullAdder U145 (w1681, w1590, IN8[4], w1682, w1683);
  FullAdder U146 (w1683, w1592, IN9[4], w1684, w1685);
  FullAdder U147 (w1685, w1594, IN10[4], w1686, w1687);
  FullAdder U148 (w1687, w1596, IN11[4], w1688, w1689);
  FullAdder U149 (w1689, w1598, IN12[4], w1690, w1691);
  FullAdder U150 (w1691, w1600, IN13[4], w1692, w1693);
  FullAdder U151 (w1693, w1602, IN14[4], w1694, w1695);
  FullAdder U152 (w1695, w1604, IN15[4], w1696, w1697);
  FullAdder U153 (w1697, w1606, IN16[4], w1698, w1699);
  FullAdder U154 (w1699, w1608, IN17[4], w1700, w1701);
  FullAdder U155 (w1701, w1610, IN18[4], w1702, w1703);
  FullAdder U156 (w1703, w1612, IN19[4], w1704, w1705);
  FullAdder U157 (w1705, w1614, IN20[4], w1706, w1707);
  FullAdder U158 (w1707, w1616, IN21[4], w1708, w1709);
  FullAdder U159 (w1709, w1618, IN22[4], w1710, w1711);
  FullAdder U160 (w1711, w1620, IN23[4], w1712, w1713);
  FullAdder U161 (w1713, w1622, IN24[4], w1714, w1715);
  FullAdder U162 (w1715, w1624, IN25[4], w1716, w1717);
  FullAdder U163 (w1717, w1626, IN26[4], w1718, w1719);
  FullAdder U164 (w1719, w1628, IN27[4], w1720, w1721);
  FullAdder U165 (w1721, w1630, IN28[4], w1722, w1723);
  FullAdder U166 (w1723, w1632, IN29[4], w1724, w1725);
  FullAdder U167 (w1725, w1634, IN30[4], w1726, w1727);
  FullAdder U168 (w1727, w1636, IN31[4], w1728, w1729);
  FullAdder U169 (w1729, w1638, IN32[4], w1730, w1731);
  FullAdder U170 (w1731, w1640, IN33[4], w1732, w1733);
  FullAdder U171 (w1733, w1642, IN34[4], w1734, w1735);
  FullAdder U172 (w1735, w1644, IN35[4], w1736, w1737);
  FullAdder U173 (w1737, w1646, IN36[4], w1738, w1739);
  FullAdder U174 (w1739, w1648, IN37[4], w1740, w1741);
  FullAdder U175 (w1741, w1650, IN38[4], w1742, w1743);
  FullAdder U176 (w1743, w1652, IN39[4], w1744, w1745);
  FullAdder U177 (w1745, w1654, IN40[4], w1746, w1747);
  FullAdder U178 (w1747, w1656, IN41[4], w1748, w1749);
  FullAdder U179 (w1749, w1658, IN42[4], w1750, w1751);
  FullAdder U180 (w1751, w1660, IN43[4], w1752, w1753);
  FullAdder U181 (w1753, w1662, IN44[4], w1754, w1755);
  FullAdder U182 (w1755, w1664, IN45[4], w1756, w1757);
  FullAdder U183 (w1757, w1666, IN46[4], w1758, w1759);
  FullAdder U184 (w1759, w1668, IN47[4], w1760, w1761);
  FullAdder U185 (w1761, w1670, IN48[2], w1762, w1763);
  FullAdder U186 (w1763, w1672, IN49[1], w1764, w1765);
  FullAdder U187 (w1765, w1673, IN50[0], w1766, w1767);
  HalfAdder U188 (w1676, IN5[5], Out1[5], w1769);
  FullAdder U189 (w1769, w1678, IN6[5], w1770, w1771);
  FullAdder U190 (w1771, w1680, IN7[5], w1772, w1773);
  FullAdder U191 (w1773, w1682, IN8[5], w1774, w1775);
  FullAdder U192 (w1775, w1684, IN9[5], w1776, w1777);
  FullAdder U193 (w1777, w1686, IN10[5], w1778, w1779);
  FullAdder U194 (w1779, w1688, IN11[5], w1780, w1781);
  FullAdder U195 (w1781, w1690, IN12[5], w1782, w1783);
  FullAdder U196 (w1783, w1692, IN13[5], w1784, w1785);
  FullAdder U197 (w1785, w1694, IN14[5], w1786, w1787);
  FullAdder U198 (w1787, w1696, IN15[5], w1788, w1789);
  FullAdder U199 (w1789, w1698, IN16[5], w1790, w1791);
  FullAdder U200 (w1791, w1700, IN17[5], w1792, w1793);
  FullAdder U201 (w1793, w1702, IN18[5], w1794, w1795);
  FullAdder U202 (w1795, w1704, IN19[5], w1796, w1797);
  FullAdder U203 (w1797, w1706, IN20[5], w1798, w1799);
  FullAdder U204 (w1799, w1708, IN21[5], w1800, w1801);
  FullAdder U205 (w1801, w1710, IN22[5], w1802, w1803);
  FullAdder U206 (w1803, w1712, IN23[5], w1804, w1805);
  FullAdder U207 (w1805, w1714, IN24[5], w1806, w1807);
  FullAdder U208 (w1807, w1716, IN25[5], w1808, w1809);
  FullAdder U209 (w1809, w1718, IN26[5], w1810, w1811);
  FullAdder U210 (w1811, w1720, IN27[5], w1812, w1813);
  FullAdder U211 (w1813, w1722, IN28[5], w1814, w1815);
  FullAdder U212 (w1815, w1724, IN29[5], w1816, w1817);
  FullAdder U213 (w1817, w1726, IN30[5], w1818, w1819);
  FullAdder U214 (w1819, w1728, IN31[5], w1820, w1821);
  FullAdder U215 (w1821, w1730, IN32[5], w1822, w1823);
  FullAdder U216 (w1823, w1732, IN33[5], w1824, w1825);
  FullAdder U217 (w1825, w1734, IN34[5], w1826, w1827);
  FullAdder U218 (w1827, w1736, IN35[5], w1828, w1829);
  FullAdder U219 (w1829, w1738, IN36[5], w1830, w1831);
  FullAdder U220 (w1831, w1740, IN37[5], w1832, w1833);
  FullAdder U221 (w1833, w1742, IN38[5], w1834, w1835);
  FullAdder U222 (w1835, w1744, IN39[5], w1836, w1837);
  FullAdder U223 (w1837, w1746, IN40[5], w1838, w1839);
  FullAdder U224 (w1839, w1748, IN41[5], w1840, w1841);
  FullAdder U225 (w1841, w1750, IN42[5], w1842, w1843);
  FullAdder U226 (w1843, w1752, IN43[5], w1844, w1845);
  FullAdder U227 (w1845, w1754, IN44[5], w1846, w1847);
  FullAdder U228 (w1847, w1756, IN45[5], w1848, w1849);
  FullAdder U229 (w1849, w1758, IN46[5], w1850, w1851);
  FullAdder U230 (w1851, w1760, IN47[5], w1852, w1853);
  FullAdder U231 (w1853, w1762, IN48[3], w1854, w1855);
  FullAdder U232 (w1855, w1764, IN49[2], w1856, w1857);
  FullAdder U233 (w1857, w1766, IN50[1], w1858, w1859);
  FullAdder U234 (w1859, w1767, IN51[0], w1860, w1861);
  HalfAdder U235 (w1770, IN6[6], Out1[6], w1863);
  FullAdder U236 (w1863, w1772, IN7[6], w1864, w1865);
  FullAdder U237 (w1865, w1774, IN8[6], w1866, w1867);
  FullAdder U238 (w1867, w1776, IN9[6], w1868, w1869);
  FullAdder U239 (w1869, w1778, IN10[6], w1870, w1871);
  FullAdder U240 (w1871, w1780, IN11[6], w1872, w1873);
  FullAdder U241 (w1873, w1782, IN12[6], w1874, w1875);
  FullAdder U242 (w1875, w1784, IN13[6], w1876, w1877);
  FullAdder U243 (w1877, w1786, IN14[6], w1878, w1879);
  FullAdder U244 (w1879, w1788, IN15[6], w1880, w1881);
  FullAdder U245 (w1881, w1790, IN16[6], w1882, w1883);
  FullAdder U246 (w1883, w1792, IN17[6], w1884, w1885);
  FullAdder U247 (w1885, w1794, IN18[6], w1886, w1887);
  FullAdder U248 (w1887, w1796, IN19[6], w1888, w1889);
  FullAdder U249 (w1889, w1798, IN20[6], w1890, w1891);
  FullAdder U250 (w1891, w1800, IN21[6], w1892, w1893);
  FullAdder U251 (w1893, w1802, IN22[6], w1894, w1895);
  FullAdder U252 (w1895, w1804, IN23[6], w1896, w1897);
  FullAdder U253 (w1897, w1806, IN24[6], w1898, w1899);
  FullAdder U254 (w1899, w1808, IN25[6], w1900, w1901);
  FullAdder U255 (w1901, w1810, IN26[6], w1902, w1903);
  FullAdder U256 (w1903, w1812, IN27[6], w1904, w1905);
  FullAdder U257 (w1905, w1814, IN28[6], w1906, w1907);
  FullAdder U258 (w1907, w1816, IN29[6], w1908, w1909);
  FullAdder U259 (w1909, w1818, IN30[6], w1910, w1911);
  FullAdder U260 (w1911, w1820, IN31[6], w1912, w1913);
  FullAdder U261 (w1913, w1822, IN32[6], w1914, w1915);
  FullAdder U262 (w1915, w1824, IN33[6], w1916, w1917);
  FullAdder U263 (w1917, w1826, IN34[6], w1918, w1919);
  FullAdder U264 (w1919, w1828, IN35[6], w1920, w1921);
  FullAdder U265 (w1921, w1830, IN36[6], w1922, w1923);
  FullAdder U266 (w1923, w1832, IN37[6], w1924, w1925);
  FullAdder U267 (w1925, w1834, IN38[6], w1926, w1927);
  FullAdder U268 (w1927, w1836, IN39[6], w1928, w1929);
  FullAdder U269 (w1929, w1838, IN40[6], w1930, w1931);
  FullAdder U270 (w1931, w1840, IN41[6], w1932, w1933);
  FullAdder U271 (w1933, w1842, IN42[6], w1934, w1935);
  FullAdder U272 (w1935, w1844, IN43[6], w1936, w1937);
  FullAdder U273 (w1937, w1846, IN44[6], w1938, w1939);
  FullAdder U274 (w1939, w1848, IN45[6], w1940, w1941);
  FullAdder U275 (w1941, w1850, IN46[6], w1942, w1943);
  FullAdder U276 (w1943, w1852, IN47[6], w1944, w1945);
  FullAdder U277 (w1945, w1854, IN48[4], w1946, w1947);
  FullAdder U278 (w1947, w1856, IN49[3], w1948, w1949);
  FullAdder U279 (w1949, w1858, IN50[2], w1950, w1951);
  FullAdder U280 (w1951, w1860, IN51[1], w1952, w1953);
  FullAdder U281 (w1953, w1861, IN52[0], w1954, w1955);
  HalfAdder U282 (w1864, IN7[7], Out1[7], w1957);
  FullAdder U283 (w1957, w1866, IN8[7], w1958, w1959);
  FullAdder U284 (w1959, w1868, IN9[7], w1960, w1961);
  FullAdder U285 (w1961, w1870, IN10[7], w1962, w1963);
  FullAdder U286 (w1963, w1872, IN11[7], w1964, w1965);
  FullAdder U287 (w1965, w1874, IN12[7], w1966, w1967);
  FullAdder U288 (w1967, w1876, IN13[7], w1968, w1969);
  FullAdder U289 (w1969, w1878, IN14[7], w1970, w1971);
  FullAdder U290 (w1971, w1880, IN15[7], w1972, w1973);
  FullAdder U291 (w1973, w1882, IN16[7], w1974, w1975);
  FullAdder U292 (w1975, w1884, IN17[7], w1976, w1977);
  FullAdder U293 (w1977, w1886, IN18[7], w1978, w1979);
  FullAdder U294 (w1979, w1888, IN19[7], w1980, w1981);
  FullAdder U295 (w1981, w1890, IN20[7], w1982, w1983);
  FullAdder U296 (w1983, w1892, IN21[7], w1984, w1985);
  FullAdder U297 (w1985, w1894, IN22[7], w1986, w1987);
  FullAdder U298 (w1987, w1896, IN23[7], w1988, w1989);
  FullAdder U299 (w1989, w1898, IN24[7], w1990, w1991);
  FullAdder U300 (w1991, w1900, IN25[7], w1992, w1993);
  FullAdder U301 (w1993, w1902, IN26[7], w1994, w1995);
  FullAdder U302 (w1995, w1904, IN27[7], w1996, w1997);
  FullAdder U303 (w1997, w1906, IN28[7], w1998, w1999);
  FullAdder U304 (w1999, w1908, IN29[7], w2000, w2001);
  FullAdder U305 (w2001, w1910, IN30[7], w2002, w2003);
  FullAdder U306 (w2003, w1912, IN31[7], w2004, w2005);
  FullAdder U307 (w2005, w1914, IN32[7], w2006, w2007);
  FullAdder U308 (w2007, w1916, IN33[7], w2008, w2009);
  FullAdder U309 (w2009, w1918, IN34[7], w2010, w2011);
  FullAdder U310 (w2011, w1920, IN35[7], w2012, w2013);
  FullAdder U311 (w2013, w1922, IN36[7], w2014, w2015);
  FullAdder U312 (w2015, w1924, IN37[7], w2016, w2017);
  FullAdder U313 (w2017, w1926, IN38[7], w2018, w2019);
  FullAdder U314 (w2019, w1928, IN39[7], w2020, w2021);
  FullAdder U315 (w2021, w1930, IN40[7], w2022, w2023);
  FullAdder U316 (w2023, w1932, IN41[7], w2024, w2025);
  FullAdder U317 (w2025, w1934, IN42[7], w2026, w2027);
  FullAdder U318 (w2027, w1936, IN43[7], w2028, w2029);
  FullAdder U319 (w2029, w1938, IN44[7], w2030, w2031);
  FullAdder U320 (w2031, w1940, IN45[7], w2032, w2033);
  FullAdder U321 (w2033, w1942, IN46[7], w2034, w2035);
  FullAdder U322 (w2035, w1944, IN47[7], w2036, w2037);
  FullAdder U323 (w2037, w1946, IN48[5], w2038, w2039);
  FullAdder U324 (w2039, w1948, IN49[4], w2040, w2041);
  FullAdder U325 (w2041, w1950, IN50[3], w2042, w2043);
  FullAdder U326 (w2043, w1952, IN51[2], w2044, w2045);
  FullAdder U327 (w2045, w1954, IN52[1], w2046, w2047);
  FullAdder U328 (w2047, w1955, IN53[0], w2048, w2049);
  HalfAdder U329 (w1958, IN8[8], Out1[8], w2051);
  FullAdder U330 (w2051, w1960, IN9[8], w2052, w2053);
  FullAdder U331 (w2053, w1962, IN10[8], w2054, w2055);
  FullAdder U332 (w2055, w1964, IN11[8], w2056, w2057);
  FullAdder U333 (w2057, w1966, IN12[8], w2058, w2059);
  FullAdder U334 (w2059, w1968, IN13[8], w2060, w2061);
  FullAdder U335 (w2061, w1970, IN14[8], w2062, w2063);
  FullAdder U336 (w2063, w1972, IN15[8], w2064, w2065);
  FullAdder U337 (w2065, w1974, IN16[8], w2066, w2067);
  FullAdder U338 (w2067, w1976, IN17[8], w2068, w2069);
  FullAdder U339 (w2069, w1978, IN18[8], w2070, w2071);
  FullAdder U340 (w2071, w1980, IN19[8], w2072, w2073);
  FullAdder U341 (w2073, w1982, IN20[8], w2074, w2075);
  FullAdder U342 (w2075, w1984, IN21[8], w2076, w2077);
  FullAdder U343 (w2077, w1986, IN22[8], w2078, w2079);
  FullAdder U344 (w2079, w1988, IN23[8], w2080, w2081);
  FullAdder U345 (w2081, w1990, IN24[8], w2082, w2083);
  FullAdder U346 (w2083, w1992, IN25[8], w2084, w2085);
  FullAdder U347 (w2085, w1994, IN26[8], w2086, w2087);
  FullAdder U348 (w2087, w1996, IN27[8], w2088, w2089);
  FullAdder U349 (w2089, w1998, IN28[8], w2090, w2091);
  FullAdder U350 (w2091, w2000, IN29[8], w2092, w2093);
  FullAdder U351 (w2093, w2002, IN30[8], w2094, w2095);
  FullAdder U352 (w2095, w2004, IN31[8], w2096, w2097);
  FullAdder U353 (w2097, w2006, IN32[8], w2098, w2099);
  FullAdder U354 (w2099, w2008, IN33[8], w2100, w2101);
  FullAdder U355 (w2101, w2010, IN34[8], w2102, w2103);
  FullAdder U356 (w2103, w2012, IN35[8], w2104, w2105);
  FullAdder U357 (w2105, w2014, IN36[8], w2106, w2107);
  FullAdder U358 (w2107, w2016, IN37[8], w2108, w2109);
  FullAdder U359 (w2109, w2018, IN38[8], w2110, w2111);
  FullAdder U360 (w2111, w2020, IN39[8], w2112, w2113);
  FullAdder U361 (w2113, w2022, IN40[8], w2114, w2115);
  FullAdder U362 (w2115, w2024, IN41[8], w2116, w2117);
  FullAdder U363 (w2117, w2026, IN42[8], w2118, w2119);
  FullAdder U364 (w2119, w2028, IN43[8], w2120, w2121);
  FullAdder U365 (w2121, w2030, IN44[8], w2122, w2123);
  FullAdder U366 (w2123, w2032, IN45[8], w2124, w2125);
  FullAdder U367 (w2125, w2034, IN46[8], w2126, w2127);
  FullAdder U368 (w2127, w2036, IN47[8], w2128, w2129);
  FullAdder U369 (w2129, w2038, IN48[6], w2130, w2131);
  FullAdder U370 (w2131, w2040, IN49[5], w2132, w2133);
  FullAdder U371 (w2133, w2042, IN50[4], w2134, w2135);
  FullAdder U372 (w2135, w2044, IN51[3], w2136, w2137);
  FullAdder U373 (w2137, w2046, IN52[2], w2138, w2139);
  FullAdder U374 (w2139, w2048, IN53[1], w2140, w2141);
  FullAdder U375 (w2141, w2049, IN54[0], w2142, w2143);
  HalfAdder U376 (w2052, IN9[9], Out1[9], w2145);
  FullAdder U377 (w2145, w2054, IN10[9], w2146, w2147);
  FullAdder U378 (w2147, w2056, IN11[9], w2148, w2149);
  FullAdder U379 (w2149, w2058, IN12[9], w2150, w2151);
  FullAdder U380 (w2151, w2060, IN13[9], w2152, w2153);
  FullAdder U381 (w2153, w2062, IN14[9], w2154, w2155);
  FullAdder U382 (w2155, w2064, IN15[9], w2156, w2157);
  FullAdder U383 (w2157, w2066, IN16[9], w2158, w2159);
  FullAdder U384 (w2159, w2068, IN17[9], w2160, w2161);
  FullAdder U385 (w2161, w2070, IN18[9], w2162, w2163);
  FullAdder U386 (w2163, w2072, IN19[9], w2164, w2165);
  FullAdder U387 (w2165, w2074, IN20[9], w2166, w2167);
  FullAdder U388 (w2167, w2076, IN21[9], w2168, w2169);
  FullAdder U389 (w2169, w2078, IN22[9], w2170, w2171);
  FullAdder U390 (w2171, w2080, IN23[9], w2172, w2173);
  FullAdder U391 (w2173, w2082, IN24[9], w2174, w2175);
  FullAdder U392 (w2175, w2084, IN25[9], w2176, w2177);
  FullAdder U393 (w2177, w2086, IN26[9], w2178, w2179);
  FullAdder U394 (w2179, w2088, IN27[9], w2180, w2181);
  FullAdder U395 (w2181, w2090, IN28[9], w2182, w2183);
  FullAdder U396 (w2183, w2092, IN29[9], w2184, w2185);
  FullAdder U397 (w2185, w2094, IN30[9], w2186, w2187);
  FullAdder U398 (w2187, w2096, IN31[9], w2188, w2189);
  FullAdder U399 (w2189, w2098, IN32[9], w2190, w2191);
  FullAdder U400 (w2191, w2100, IN33[9], w2192, w2193);
  FullAdder U401 (w2193, w2102, IN34[9], w2194, w2195);
  FullAdder U402 (w2195, w2104, IN35[9], w2196, w2197);
  FullAdder U403 (w2197, w2106, IN36[9], w2198, w2199);
  FullAdder U404 (w2199, w2108, IN37[9], w2200, w2201);
  FullAdder U405 (w2201, w2110, IN38[9], w2202, w2203);
  FullAdder U406 (w2203, w2112, IN39[9], w2204, w2205);
  FullAdder U407 (w2205, w2114, IN40[9], w2206, w2207);
  FullAdder U408 (w2207, w2116, IN41[9], w2208, w2209);
  FullAdder U409 (w2209, w2118, IN42[9], w2210, w2211);
  FullAdder U410 (w2211, w2120, IN43[9], w2212, w2213);
  FullAdder U411 (w2213, w2122, IN44[9], w2214, w2215);
  FullAdder U412 (w2215, w2124, IN45[9], w2216, w2217);
  FullAdder U413 (w2217, w2126, IN46[9], w2218, w2219);
  FullAdder U414 (w2219, w2128, IN47[9], w2220, w2221);
  FullAdder U415 (w2221, w2130, IN48[7], w2222, w2223);
  FullAdder U416 (w2223, w2132, IN49[6], w2224, w2225);
  FullAdder U417 (w2225, w2134, IN50[5], w2226, w2227);
  FullAdder U418 (w2227, w2136, IN51[4], w2228, w2229);
  FullAdder U419 (w2229, w2138, IN52[3], w2230, w2231);
  FullAdder U420 (w2231, w2140, IN53[2], w2232, w2233);
  FullAdder U421 (w2233, w2142, IN54[1], w2234, w2235);
  FullAdder U422 (w2235, w2143, IN55[0], w2236, w2237);
  HalfAdder U423 (w2146, IN10[10], Out1[10], w2239);
  FullAdder U424 (w2239, w2148, IN11[10], w2240, w2241);
  FullAdder U425 (w2241, w2150, IN12[10], w2242, w2243);
  FullAdder U426 (w2243, w2152, IN13[10], w2244, w2245);
  FullAdder U427 (w2245, w2154, IN14[10], w2246, w2247);
  FullAdder U428 (w2247, w2156, IN15[10], w2248, w2249);
  FullAdder U429 (w2249, w2158, IN16[10], w2250, w2251);
  FullAdder U430 (w2251, w2160, IN17[10], w2252, w2253);
  FullAdder U431 (w2253, w2162, IN18[10], w2254, w2255);
  FullAdder U432 (w2255, w2164, IN19[10], w2256, w2257);
  FullAdder U433 (w2257, w2166, IN20[10], w2258, w2259);
  FullAdder U434 (w2259, w2168, IN21[10], w2260, w2261);
  FullAdder U435 (w2261, w2170, IN22[10], w2262, w2263);
  FullAdder U436 (w2263, w2172, IN23[10], w2264, w2265);
  FullAdder U437 (w2265, w2174, IN24[10], w2266, w2267);
  FullAdder U438 (w2267, w2176, IN25[10], w2268, w2269);
  FullAdder U439 (w2269, w2178, IN26[10], w2270, w2271);
  FullAdder U440 (w2271, w2180, IN27[10], w2272, w2273);
  FullAdder U441 (w2273, w2182, IN28[10], w2274, w2275);
  FullAdder U442 (w2275, w2184, IN29[10], w2276, w2277);
  FullAdder U443 (w2277, w2186, IN30[10], w2278, w2279);
  FullAdder U444 (w2279, w2188, IN31[10], w2280, w2281);
  FullAdder U445 (w2281, w2190, IN32[10], w2282, w2283);
  FullAdder U446 (w2283, w2192, IN33[10], w2284, w2285);
  FullAdder U447 (w2285, w2194, IN34[10], w2286, w2287);
  FullAdder U448 (w2287, w2196, IN35[10], w2288, w2289);
  FullAdder U449 (w2289, w2198, IN36[10], w2290, w2291);
  FullAdder U450 (w2291, w2200, IN37[10], w2292, w2293);
  FullAdder U451 (w2293, w2202, IN38[10], w2294, w2295);
  FullAdder U452 (w2295, w2204, IN39[10], w2296, w2297);
  FullAdder U453 (w2297, w2206, IN40[10], w2298, w2299);
  FullAdder U454 (w2299, w2208, IN41[10], w2300, w2301);
  FullAdder U455 (w2301, w2210, IN42[10], w2302, w2303);
  FullAdder U456 (w2303, w2212, IN43[10], w2304, w2305);
  FullAdder U457 (w2305, w2214, IN44[10], w2306, w2307);
  FullAdder U458 (w2307, w2216, IN45[10], w2308, w2309);
  FullAdder U459 (w2309, w2218, IN46[10], w2310, w2311);
  FullAdder U460 (w2311, w2220, IN47[10], w2312, w2313);
  FullAdder U461 (w2313, w2222, IN48[8], w2314, w2315);
  FullAdder U462 (w2315, w2224, IN49[7], w2316, w2317);
  FullAdder U463 (w2317, w2226, IN50[6], w2318, w2319);
  FullAdder U464 (w2319, w2228, IN51[5], w2320, w2321);
  FullAdder U465 (w2321, w2230, IN52[4], w2322, w2323);
  FullAdder U466 (w2323, w2232, IN53[3], w2324, w2325);
  FullAdder U467 (w2325, w2234, IN54[2], w2326, w2327);
  FullAdder U468 (w2327, w2236, IN55[1], w2328, w2329);
  FullAdder U469 (w2329, w2237, IN56[0], w2330, w2331);
  HalfAdder U470 (w2240, IN11[11], Out1[11], w2333);
  FullAdder U471 (w2333, w2242, IN12[11], w2334, w2335);
  FullAdder U472 (w2335, w2244, IN13[11], w2336, w2337);
  FullAdder U473 (w2337, w2246, IN14[11], w2338, w2339);
  FullAdder U474 (w2339, w2248, IN15[11], w2340, w2341);
  FullAdder U475 (w2341, w2250, IN16[11], w2342, w2343);
  FullAdder U476 (w2343, w2252, IN17[11], w2344, w2345);
  FullAdder U477 (w2345, w2254, IN18[11], w2346, w2347);
  FullAdder U478 (w2347, w2256, IN19[11], w2348, w2349);
  FullAdder U479 (w2349, w2258, IN20[11], w2350, w2351);
  FullAdder U480 (w2351, w2260, IN21[11], w2352, w2353);
  FullAdder U481 (w2353, w2262, IN22[11], w2354, w2355);
  FullAdder U482 (w2355, w2264, IN23[11], w2356, w2357);
  FullAdder U483 (w2357, w2266, IN24[11], w2358, w2359);
  FullAdder U484 (w2359, w2268, IN25[11], w2360, w2361);
  FullAdder U485 (w2361, w2270, IN26[11], w2362, w2363);
  FullAdder U486 (w2363, w2272, IN27[11], w2364, w2365);
  FullAdder U487 (w2365, w2274, IN28[11], w2366, w2367);
  FullAdder U488 (w2367, w2276, IN29[11], w2368, w2369);
  FullAdder U489 (w2369, w2278, IN30[11], w2370, w2371);
  FullAdder U490 (w2371, w2280, IN31[11], w2372, w2373);
  FullAdder U491 (w2373, w2282, IN32[11], w2374, w2375);
  FullAdder U492 (w2375, w2284, IN33[11], w2376, w2377);
  FullAdder U493 (w2377, w2286, IN34[11], w2378, w2379);
  FullAdder U494 (w2379, w2288, IN35[11], w2380, w2381);
  FullAdder U495 (w2381, w2290, IN36[11], w2382, w2383);
  FullAdder U496 (w2383, w2292, IN37[11], w2384, w2385);
  FullAdder U497 (w2385, w2294, IN38[11], w2386, w2387);
  FullAdder U498 (w2387, w2296, IN39[11], w2388, w2389);
  FullAdder U499 (w2389, w2298, IN40[11], w2390, w2391);
  FullAdder U500 (w2391, w2300, IN41[11], w2392, w2393);
  FullAdder U501 (w2393, w2302, IN42[11], w2394, w2395);
  FullAdder U502 (w2395, w2304, IN43[11], w2396, w2397);
  FullAdder U503 (w2397, w2306, IN44[11], w2398, w2399);
  FullAdder U504 (w2399, w2308, IN45[11], w2400, w2401);
  FullAdder U505 (w2401, w2310, IN46[11], w2402, w2403);
  FullAdder U506 (w2403, w2312, IN47[11], w2404, w2405);
  FullAdder U507 (w2405, w2314, IN48[9], w2406, w2407);
  FullAdder U508 (w2407, w2316, IN49[8], w2408, w2409);
  FullAdder U509 (w2409, w2318, IN50[7], w2410, w2411);
  FullAdder U510 (w2411, w2320, IN51[6], w2412, w2413);
  FullAdder U511 (w2413, w2322, IN52[5], w2414, w2415);
  FullAdder U512 (w2415, w2324, IN53[4], w2416, w2417);
  FullAdder U513 (w2417, w2326, IN54[3], w2418, w2419);
  FullAdder U514 (w2419, w2328, IN55[2], w2420, w2421);
  FullAdder U515 (w2421, w2330, IN56[1], w2422, w2423);
  FullAdder U516 (w2423, w2331, IN57[0], w2424, w2425);
  HalfAdder U517 (w2334, IN12[12], Out1[12], w2427);
  FullAdder U518 (w2427, w2336, IN13[12], w2428, w2429);
  FullAdder U519 (w2429, w2338, IN14[12], w2430, w2431);
  FullAdder U520 (w2431, w2340, IN15[12], w2432, w2433);
  FullAdder U521 (w2433, w2342, IN16[12], w2434, w2435);
  FullAdder U522 (w2435, w2344, IN17[12], w2436, w2437);
  FullAdder U523 (w2437, w2346, IN18[12], w2438, w2439);
  FullAdder U524 (w2439, w2348, IN19[12], w2440, w2441);
  FullAdder U525 (w2441, w2350, IN20[12], w2442, w2443);
  FullAdder U526 (w2443, w2352, IN21[12], w2444, w2445);
  FullAdder U527 (w2445, w2354, IN22[12], w2446, w2447);
  FullAdder U528 (w2447, w2356, IN23[12], w2448, w2449);
  FullAdder U529 (w2449, w2358, IN24[12], w2450, w2451);
  FullAdder U530 (w2451, w2360, IN25[12], w2452, w2453);
  FullAdder U531 (w2453, w2362, IN26[12], w2454, w2455);
  FullAdder U532 (w2455, w2364, IN27[12], w2456, w2457);
  FullAdder U533 (w2457, w2366, IN28[12], w2458, w2459);
  FullAdder U534 (w2459, w2368, IN29[12], w2460, w2461);
  FullAdder U535 (w2461, w2370, IN30[12], w2462, w2463);
  FullAdder U536 (w2463, w2372, IN31[12], w2464, w2465);
  FullAdder U537 (w2465, w2374, IN32[12], w2466, w2467);
  FullAdder U538 (w2467, w2376, IN33[12], w2468, w2469);
  FullAdder U539 (w2469, w2378, IN34[12], w2470, w2471);
  FullAdder U540 (w2471, w2380, IN35[12], w2472, w2473);
  FullAdder U541 (w2473, w2382, IN36[12], w2474, w2475);
  FullAdder U542 (w2475, w2384, IN37[12], w2476, w2477);
  FullAdder U543 (w2477, w2386, IN38[12], w2478, w2479);
  FullAdder U544 (w2479, w2388, IN39[12], w2480, w2481);
  FullAdder U545 (w2481, w2390, IN40[12], w2482, w2483);
  FullAdder U546 (w2483, w2392, IN41[12], w2484, w2485);
  FullAdder U547 (w2485, w2394, IN42[12], w2486, w2487);
  FullAdder U548 (w2487, w2396, IN43[12], w2488, w2489);
  FullAdder U549 (w2489, w2398, IN44[12], w2490, w2491);
  FullAdder U550 (w2491, w2400, IN45[12], w2492, w2493);
  FullAdder U551 (w2493, w2402, IN46[12], w2494, w2495);
  FullAdder U552 (w2495, w2404, IN47[12], w2496, w2497);
  FullAdder U553 (w2497, w2406, IN48[10], w2498, w2499);
  FullAdder U554 (w2499, w2408, IN49[9], w2500, w2501);
  FullAdder U555 (w2501, w2410, IN50[8], w2502, w2503);
  FullAdder U556 (w2503, w2412, IN51[7], w2504, w2505);
  FullAdder U557 (w2505, w2414, IN52[6], w2506, w2507);
  FullAdder U558 (w2507, w2416, IN53[5], w2508, w2509);
  FullAdder U559 (w2509, w2418, IN54[4], w2510, w2511);
  FullAdder U560 (w2511, w2420, IN55[3], w2512, w2513);
  FullAdder U561 (w2513, w2422, IN56[2], w2514, w2515);
  FullAdder U562 (w2515, w2424, IN57[1], w2516, w2517);
  FullAdder U563 (w2517, w2425, IN58[0], w2518, w2519);
  HalfAdder U564 (w2428, IN13[13], Out1[13], w2521);
  FullAdder U565 (w2521, w2430, IN14[13], w2522, w2523);
  FullAdder U566 (w2523, w2432, IN15[13], w2524, w2525);
  FullAdder U567 (w2525, w2434, IN16[13], w2526, w2527);
  FullAdder U568 (w2527, w2436, IN17[13], w2528, w2529);
  FullAdder U569 (w2529, w2438, IN18[13], w2530, w2531);
  FullAdder U570 (w2531, w2440, IN19[13], w2532, w2533);
  FullAdder U571 (w2533, w2442, IN20[13], w2534, w2535);
  FullAdder U572 (w2535, w2444, IN21[13], w2536, w2537);
  FullAdder U573 (w2537, w2446, IN22[13], w2538, w2539);
  FullAdder U574 (w2539, w2448, IN23[13], w2540, w2541);
  FullAdder U575 (w2541, w2450, IN24[13], w2542, w2543);
  FullAdder U576 (w2543, w2452, IN25[13], w2544, w2545);
  FullAdder U577 (w2545, w2454, IN26[13], w2546, w2547);
  FullAdder U578 (w2547, w2456, IN27[13], w2548, w2549);
  FullAdder U579 (w2549, w2458, IN28[13], w2550, w2551);
  FullAdder U580 (w2551, w2460, IN29[13], w2552, w2553);
  FullAdder U581 (w2553, w2462, IN30[13], w2554, w2555);
  FullAdder U582 (w2555, w2464, IN31[13], w2556, w2557);
  FullAdder U583 (w2557, w2466, IN32[13], w2558, w2559);
  FullAdder U584 (w2559, w2468, IN33[13], w2560, w2561);
  FullAdder U585 (w2561, w2470, IN34[13], w2562, w2563);
  FullAdder U586 (w2563, w2472, IN35[13], w2564, w2565);
  FullAdder U587 (w2565, w2474, IN36[13], w2566, w2567);
  FullAdder U588 (w2567, w2476, IN37[13], w2568, w2569);
  FullAdder U589 (w2569, w2478, IN38[13], w2570, w2571);
  FullAdder U590 (w2571, w2480, IN39[13], w2572, w2573);
  FullAdder U591 (w2573, w2482, IN40[13], w2574, w2575);
  FullAdder U592 (w2575, w2484, IN41[13], w2576, w2577);
  FullAdder U593 (w2577, w2486, IN42[13], w2578, w2579);
  FullAdder U594 (w2579, w2488, IN43[13], w2580, w2581);
  FullAdder U595 (w2581, w2490, IN44[13], w2582, w2583);
  FullAdder U596 (w2583, w2492, IN45[13], w2584, w2585);
  FullAdder U597 (w2585, w2494, IN46[13], w2586, w2587);
  FullAdder U598 (w2587, w2496, IN47[13], w2588, w2589);
  FullAdder U599 (w2589, w2498, IN48[11], w2590, w2591);
  FullAdder U600 (w2591, w2500, IN49[10], w2592, w2593);
  FullAdder U601 (w2593, w2502, IN50[9], w2594, w2595);
  FullAdder U602 (w2595, w2504, IN51[8], w2596, w2597);
  FullAdder U603 (w2597, w2506, IN52[7], w2598, w2599);
  FullAdder U604 (w2599, w2508, IN53[6], w2600, w2601);
  FullAdder U605 (w2601, w2510, IN54[5], w2602, w2603);
  FullAdder U606 (w2603, w2512, IN55[4], w2604, w2605);
  FullAdder U607 (w2605, w2514, IN56[3], w2606, w2607);
  FullAdder U608 (w2607, w2516, IN57[2], w2608, w2609);
  FullAdder U609 (w2609, w2518, IN58[1], w2610, w2611);
  FullAdder U610 (w2611, w2519, IN59[0], w2612, w2613);
  HalfAdder U611 (w2522, IN14[14], Out1[14], w2615);
  FullAdder U612 (w2615, w2524, IN15[14], w2616, w2617);
  FullAdder U613 (w2617, w2526, IN16[14], w2618, w2619);
  FullAdder U614 (w2619, w2528, IN17[14], w2620, w2621);
  FullAdder U615 (w2621, w2530, IN18[14], w2622, w2623);
  FullAdder U616 (w2623, w2532, IN19[14], w2624, w2625);
  FullAdder U617 (w2625, w2534, IN20[14], w2626, w2627);
  FullAdder U618 (w2627, w2536, IN21[14], w2628, w2629);
  FullAdder U619 (w2629, w2538, IN22[14], w2630, w2631);
  FullAdder U620 (w2631, w2540, IN23[14], w2632, w2633);
  FullAdder U621 (w2633, w2542, IN24[14], w2634, w2635);
  FullAdder U622 (w2635, w2544, IN25[14], w2636, w2637);
  FullAdder U623 (w2637, w2546, IN26[14], w2638, w2639);
  FullAdder U624 (w2639, w2548, IN27[14], w2640, w2641);
  FullAdder U625 (w2641, w2550, IN28[14], w2642, w2643);
  FullAdder U626 (w2643, w2552, IN29[14], w2644, w2645);
  FullAdder U627 (w2645, w2554, IN30[14], w2646, w2647);
  FullAdder U628 (w2647, w2556, IN31[14], w2648, w2649);
  FullAdder U629 (w2649, w2558, IN32[14], w2650, w2651);
  FullAdder U630 (w2651, w2560, IN33[14], w2652, w2653);
  FullAdder U631 (w2653, w2562, IN34[14], w2654, w2655);
  FullAdder U632 (w2655, w2564, IN35[14], w2656, w2657);
  FullAdder U633 (w2657, w2566, IN36[14], w2658, w2659);
  FullAdder U634 (w2659, w2568, IN37[14], w2660, w2661);
  FullAdder U635 (w2661, w2570, IN38[14], w2662, w2663);
  FullAdder U636 (w2663, w2572, IN39[14], w2664, w2665);
  FullAdder U637 (w2665, w2574, IN40[14], w2666, w2667);
  FullAdder U638 (w2667, w2576, IN41[14], w2668, w2669);
  FullAdder U639 (w2669, w2578, IN42[14], w2670, w2671);
  FullAdder U640 (w2671, w2580, IN43[14], w2672, w2673);
  FullAdder U641 (w2673, w2582, IN44[14], w2674, w2675);
  FullAdder U642 (w2675, w2584, IN45[14], w2676, w2677);
  FullAdder U643 (w2677, w2586, IN46[14], w2678, w2679);
  FullAdder U644 (w2679, w2588, IN47[14], w2680, w2681);
  FullAdder U645 (w2681, w2590, IN48[12], w2682, w2683);
  FullAdder U646 (w2683, w2592, IN49[11], w2684, w2685);
  FullAdder U647 (w2685, w2594, IN50[10], w2686, w2687);
  FullAdder U648 (w2687, w2596, IN51[9], w2688, w2689);
  FullAdder U649 (w2689, w2598, IN52[8], w2690, w2691);
  FullAdder U650 (w2691, w2600, IN53[7], w2692, w2693);
  FullAdder U651 (w2693, w2602, IN54[6], w2694, w2695);
  FullAdder U652 (w2695, w2604, IN55[5], w2696, w2697);
  FullAdder U653 (w2697, w2606, IN56[4], w2698, w2699);
  FullAdder U654 (w2699, w2608, IN57[3], w2700, w2701);
  FullAdder U655 (w2701, w2610, IN58[2], w2702, w2703);
  FullAdder U656 (w2703, w2612, IN59[1], w2704, w2705);
  FullAdder U657 (w2705, w2613, IN60[0], w2706, w2707);
  HalfAdder U658 (w2616, IN15[15], Out1[15], w2709);
  FullAdder U659 (w2709, w2618, IN16[15], w2710, w2711);
  FullAdder U660 (w2711, w2620, IN17[15], w2712, w2713);
  FullAdder U661 (w2713, w2622, IN18[15], w2714, w2715);
  FullAdder U662 (w2715, w2624, IN19[15], w2716, w2717);
  FullAdder U663 (w2717, w2626, IN20[15], w2718, w2719);
  FullAdder U664 (w2719, w2628, IN21[15], w2720, w2721);
  FullAdder U665 (w2721, w2630, IN22[15], w2722, w2723);
  FullAdder U666 (w2723, w2632, IN23[15], w2724, w2725);
  FullAdder U667 (w2725, w2634, IN24[15], w2726, w2727);
  FullAdder U668 (w2727, w2636, IN25[15], w2728, w2729);
  FullAdder U669 (w2729, w2638, IN26[15], w2730, w2731);
  FullAdder U670 (w2731, w2640, IN27[15], w2732, w2733);
  FullAdder U671 (w2733, w2642, IN28[15], w2734, w2735);
  FullAdder U672 (w2735, w2644, IN29[15], w2736, w2737);
  FullAdder U673 (w2737, w2646, IN30[15], w2738, w2739);
  FullAdder U674 (w2739, w2648, IN31[15], w2740, w2741);
  FullAdder U675 (w2741, w2650, IN32[15], w2742, w2743);
  FullAdder U676 (w2743, w2652, IN33[15], w2744, w2745);
  FullAdder U677 (w2745, w2654, IN34[15], w2746, w2747);
  FullAdder U678 (w2747, w2656, IN35[15], w2748, w2749);
  FullAdder U679 (w2749, w2658, IN36[15], w2750, w2751);
  FullAdder U680 (w2751, w2660, IN37[15], w2752, w2753);
  FullAdder U681 (w2753, w2662, IN38[15], w2754, w2755);
  FullAdder U682 (w2755, w2664, IN39[15], w2756, w2757);
  FullAdder U683 (w2757, w2666, IN40[15], w2758, w2759);
  FullAdder U684 (w2759, w2668, IN41[15], w2760, w2761);
  FullAdder U685 (w2761, w2670, IN42[15], w2762, w2763);
  FullAdder U686 (w2763, w2672, IN43[15], w2764, w2765);
  FullAdder U687 (w2765, w2674, IN44[15], w2766, w2767);
  FullAdder U688 (w2767, w2676, IN45[15], w2768, w2769);
  FullAdder U689 (w2769, w2678, IN46[15], w2770, w2771);
  FullAdder U690 (w2771, w2680, IN47[15], w2772, w2773);
  FullAdder U691 (w2773, w2682, IN48[13], w2774, w2775);
  FullAdder U692 (w2775, w2684, IN49[12], w2776, w2777);
  FullAdder U693 (w2777, w2686, IN50[11], w2778, w2779);
  FullAdder U694 (w2779, w2688, IN51[10], w2780, w2781);
  FullAdder U695 (w2781, w2690, IN52[9], w2782, w2783);
  FullAdder U696 (w2783, w2692, IN53[8], w2784, w2785);
  FullAdder U697 (w2785, w2694, IN54[7], w2786, w2787);
  FullAdder U698 (w2787, w2696, IN55[6], w2788, w2789);
  FullAdder U699 (w2789, w2698, IN56[5], w2790, w2791);
  FullAdder U700 (w2791, w2700, IN57[4], w2792, w2793);
  FullAdder U701 (w2793, w2702, IN58[3], w2794, w2795);
  FullAdder U702 (w2795, w2704, IN59[2], w2796, w2797);
  FullAdder U703 (w2797, w2706, IN60[1], w2798, w2799);
  FullAdder U704 (w2799, w2707, IN61[0], w2800, w2801);
  HalfAdder U705 (w2710, IN16[16], Out1[16], w2803);
  FullAdder U706 (w2803, w2712, IN17[16], w2804, w2805);
  FullAdder U707 (w2805, w2714, IN18[16], w2806, w2807);
  FullAdder U708 (w2807, w2716, IN19[16], w2808, w2809);
  FullAdder U709 (w2809, w2718, IN20[16], w2810, w2811);
  FullAdder U710 (w2811, w2720, IN21[16], w2812, w2813);
  FullAdder U711 (w2813, w2722, IN22[16], w2814, w2815);
  FullAdder U712 (w2815, w2724, IN23[16], w2816, w2817);
  FullAdder U713 (w2817, w2726, IN24[16], w2818, w2819);
  FullAdder U714 (w2819, w2728, IN25[16], w2820, w2821);
  FullAdder U715 (w2821, w2730, IN26[16], w2822, w2823);
  FullAdder U716 (w2823, w2732, IN27[16], w2824, w2825);
  FullAdder U717 (w2825, w2734, IN28[16], w2826, w2827);
  FullAdder U718 (w2827, w2736, IN29[16], w2828, w2829);
  FullAdder U719 (w2829, w2738, IN30[16], w2830, w2831);
  FullAdder U720 (w2831, w2740, IN31[16], w2832, w2833);
  FullAdder U721 (w2833, w2742, IN32[16], w2834, w2835);
  FullAdder U722 (w2835, w2744, IN33[16], w2836, w2837);
  FullAdder U723 (w2837, w2746, IN34[16], w2838, w2839);
  FullAdder U724 (w2839, w2748, IN35[16], w2840, w2841);
  FullAdder U725 (w2841, w2750, IN36[16], w2842, w2843);
  FullAdder U726 (w2843, w2752, IN37[16], w2844, w2845);
  FullAdder U727 (w2845, w2754, IN38[16], w2846, w2847);
  FullAdder U728 (w2847, w2756, IN39[16], w2848, w2849);
  FullAdder U729 (w2849, w2758, IN40[16], w2850, w2851);
  FullAdder U730 (w2851, w2760, IN41[16], w2852, w2853);
  FullAdder U731 (w2853, w2762, IN42[16], w2854, w2855);
  FullAdder U732 (w2855, w2764, IN43[16], w2856, w2857);
  FullAdder U733 (w2857, w2766, IN44[16], w2858, w2859);
  FullAdder U734 (w2859, w2768, IN45[16], w2860, w2861);
  FullAdder U735 (w2861, w2770, IN46[16], w2862, w2863);
  FullAdder U736 (w2863, w2772, IN47[16], w2864, w2865);
  FullAdder U737 (w2865, w2774, IN48[14], w2866, w2867);
  FullAdder U738 (w2867, w2776, IN49[13], w2868, w2869);
  FullAdder U739 (w2869, w2778, IN50[12], w2870, w2871);
  FullAdder U740 (w2871, w2780, IN51[11], w2872, w2873);
  FullAdder U741 (w2873, w2782, IN52[10], w2874, w2875);
  FullAdder U742 (w2875, w2784, IN53[9], w2876, w2877);
  FullAdder U743 (w2877, w2786, IN54[8], w2878, w2879);
  FullAdder U744 (w2879, w2788, IN55[7], w2880, w2881);
  FullAdder U745 (w2881, w2790, IN56[6], w2882, w2883);
  FullAdder U746 (w2883, w2792, IN57[5], w2884, w2885);
  FullAdder U747 (w2885, w2794, IN58[4], w2886, w2887);
  FullAdder U748 (w2887, w2796, IN59[3], w2888, w2889);
  FullAdder U749 (w2889, w2798, IN60[2], w2890, w2891);
  FullAdder U750 (w2891, w2800, IN61[1], w2892, w2893);
  FullAdder U751 (w2893, w2801, IN62[0], w2894, w2895);
  HalfAdder U752 (w2804, IN17[17], Out1[17], w2897);
  FullAdder U753 (w2897, w2806, IN18[17], w2898, w2899);
  FullAdder U754 (w2899, w2808, IN19[17], w2900, w2901);
  FullAdder U755 (w2901, w2810, IN20[17], w2902, w2903);
  FullAdder U756 (w2903, w2812, IN21[17], w2904, w2905);
  FullAdder U757 (w2905, w2814, IN22[17], w2906, w2907);
  FullAdder U758 (w2907, w2816, IN23[17], w2908, w2909);
  FullAdder U759 (w2909, w2818, IN24[17], w2910, w2911);
  FullAdder U760 (w2911, w2820, IN25[17], w2912, w2913);
  FullAdder U761 (w2913, w2822, IN26[17], w2914, w2915);
  FullAdder U762 (w2915, w2824, IN27[17], w2916, w2917);
  FullAdder U763 (w2917, w2826, IN28[17], w2918, w2919);
  FullAdder U764 (w2919, w2828, IN29[17], w2920, w2921);
  FullAdder U765 (w2921, w2830, IN30[17], w2922, w2923);
  FullAdder U766 (w2923, w2832, IN31[17], w2924, w2925);
  FullAdder U767 (w2925, w2834, IN32[17], w2926, w2927);
  FullAdder U768 (w2927, w2836, IN33[17], w2928, w2929);
  FullAdder U769 (w2929, w2838, IN34[17], w2930, w2931);
  FullAdder U770 (w2931, w2840, IN35[17], w2932, w2933);
  FullAdder U771 (w2933, w2842, IN36[17], w2934, w2935);
  FullAdder U772 (w2935, w2844, IN37[17], w2936, w2937);
  FullAdder U773 (w2937, w2846, IN38[17], w2938, w2939);
  FullAdder U774 (w2939, w2848, IN39[17], w2940, w2941);
  FullAdder U775 (w2941, w2850, IN40[17], w2942, w2943);
  FullAdder U776 (w2943, w2852, IN41[17], w2944, w2945);
  FullAdder U777 (w2945, w2854, IN42[17], w2946, w2947);
  FullAdder U778 (w2947, w2856, IN43[17], w2948, w2949);
  FullAdder U779 (w2949, w2858, IN44[17], w2950, w2951);
  FullAdder U780 (w2951, w2860, IN45[17], w2952, w2953);
  FullAdder U781 (w2953, w2862, IN46[17], w2954, w2955);
  FullAdder U782 (w2955, w2864, IN47[17], w2956, w2957);
  FullAdder U783 (w2957, w2866, IN48[15], w2958, w2959);
  FullAdder U784 (w2959, w2868, IN49[14], w2960, w2961);
  FullAdder U785 (w2961, w2870, IN50[13], w2962, w2963);
  FullAdder U786 (w2963, w2872, IN51[12], w2964, w2965);
  FullAdder U787 (w2965, w2874, IN52[11], w2966, w2967);
  FullAdder U788 (w2967, w2876, IN53[10], w2968, w2969);
  FullAdder U789 (w2969, w2878, IN54[9], w2970, w2971);
  FullAdder U790 (w2971, w2880, IN55[8], w2972, w2973);
  FullAdder U791 (w2973, w2882, IN56[7], w2974, w2975);
  FullAdder U792 (w2975, w2884, IN57[6], w2976, w2977);
  FullAdder U793 (w2977, w2886, IN58[5], w2978, w2979);
  FullAdder U794 (w2979, w2888, IN59[4], w2980, w2981);
  FullAdder U795 (w2981, w2890, IN60[3], w2982, w2983);
  FullAdder U796 (w2983, w2892, IN61[2], w2984, w2985);
  FullAdder U797 (w2985, w2894, IN62[1], w2986, w2987);
  FullAdder U798 (w2987, w2895, IN63[0], w2988, w2989);
  HalfAdder U799 (w2898, IN18[18], Out1[18], w2991);
  FullAdder U800 (w2991, w2900, IN19[18], w2992, w2993);
  FullAdder U801 (w2993, w2902, IN20[18], w2994, w2995);
  FullAdder U802 (w2995, w2904, IN21[18], w2996, w2997);
  FullAdder U803 (w2997, w2906, IN22[18], w2998, w2999);
  FullAdder U804 (w2999, w2908, IN23[18], w3000, w3001);
  FullAdder U805 (w3001, w2910, IN24[18], w3002, w3003);
  FullAdder U806 (w3003, w2912, IN25[18], w3004, w3005);
  FullAdder U807 (w3005, w2914, IN26[18], w3006, w3007);
  FullAdder U808 (w3007, w2916, IN27[18], w3008, w3009);
  FullAdder U809 (w3009, w2918, IN28[18], w3010, w3011);
  FullAdder U810 (w3011, w2920, IN29[18], w3012, w3013);
  FullAdder U811 (w3013, w2922, IN30[18], w3014, w3015);
  FullAdder U812 (w3015, w2924, IN31[18], w3016, w3017);
  FullAdder U813 (w3017, w2926, IN32[18], w3018, w3019);
  FullAdder U814 (w3019, w2928, IN33[18], w3020, w3021);
  FullAdder U815 (w3021, w2930, IN34[18], w3022, w3023);
  FullAdder U816 (w3023, w2932, IN35[18], w3024, w3025);
  FullAdder U817 (w3025, w2934, IN36[18], w3026, w3027);
  FullAdder U818 (w3027, w2936, IN37[18], w3028, w3029);
  FullAdder U819 (w3029, w2938, IN38[18], w3030, w3031);
  FullAdder U820 (w3031, w2940, IN39[18], w3032, w3033);
  FullAdder U821 (w3033, w2942, IN40[18], w3034, w3035);
  FullAdder U822 (w3035, w2944, IN41[18], w3036, w3037);
  FullAdder U823 (w3037, w2946, IN42[18], w3038, w3039);
  FullAdder U824 (w3039, w2948, IN43[18], w3040, w3041);
  FullAdder U825 (w3041, w2950, IN44[18], w3042, w3043);
  FullAdder U826 (w3043, w2952, IN45[18], w3044, w3045);
  FullAdder U827 (w3045, w2954, IN46[18], w3046, w3047);
  FullAdder U828 (w3047, w2956, IN47[18], w3048, w3049);
  FullAdder U829 (w3049, w2958, IN48[16], w3050, w3051);
  FullAdder U830 (w3051, w2960, IN49[15], w3052, w3053);
  FullAdder U831 (w3053, w2962, IN50[14], w3054, w3055);
  FullAdder U832 (w3055, w2964, IN51[13], w3056, w3057);
  FullAdder U833 (w3057, w2966, IN52[12], w3058, w3059);
  FullAdder U834 (w3059, w2968, IN53[11], w3060, w3061);
  FullAdder U835 (w3061, w2970, IN54[10], w3062, w3063);
  FullAdder U836 (w3063, w2972, IN55[9], w3064, w3065);
  FullAdder U837 (w3065, w2974, IN56[8], w3066, w3067);
  FullAdder U838 (w3067, w2976, IN57[7], w3068, w3069);
  FullAdder U839 (w3069, w2978, IN58[6], w3070, w3071);
  FullAdder U840 (w3071, w2980, IN59[5], w3072, w3073);
  FullAdder U841 (w3073, w2982, IN60[4], w3074, w3075);
  FullAdder U842 (w3075, w2984, IN61[3], w3076, w3077);
  FullAdder U843 (w3077, w2986, IN62[2], w3078, w3079);
  FullAdder U844 (w3079, w2988, IN63[1], w3080, w3081);
  FullAdder U845 (w3081, w2989, IN64[0], w3082, w3083);
  HalfAdder U846 (w2992, IN19[19], Out1[19], w3085);
  FullAdder U847 (w3085, w2994, IN20[19], w3086, w3087);
  FullAdder U848 (w3087, w2996, IN21[19], w3088, w3089);
  FullAdder U849 (w3089, w2998, IN22[19], w3090, w3091);
  FullAdder U850 (w3091, w3000, IN23[19], w3092, w3093);
  FullAdder U851 (w3093, w3002, IN24[19], w3094, w3095);
  FullAdder U852 (w3095, w3004, IN25[19], w3096, w3097);
  FullAdder U853 (w3097, w3006, IN26[19], w3098, w3099);
  FullAdder U854 (w3099, w3008, IN27[19], w3100, w3101);
  FullAdder U855 (w3101, w3010, IN28[19], w3102, w3103);
  FullAdder U856 (w3103, w3012, IN29[19], w3104, w3105);
  FullAdder U857 (w3105, w3014, IN30[19], w3106, w3107);
  FullAdder U858 (w3107, w3016, IN31[19], w3108, w3109);
  FullAdder U859 (w3109, w3018, IN32[19], w3110, w3111);
  FullAdder U860 (w3111, w3020, IN33[19], w3112, w3113);
  FullAdder U861 (w3113, w3022, IN34[19], w3114, w3115);
  FullAdder U862 (w3115, w3024, IN35[19], w3116, w3117);
  FullAdder U863 (w3117, w3026, IN36[19], w3118, w3119);
  FullAdder U864 (w3119, w3028, IN37[19], w3120, w3121);
  FullAdder U865 (w3121, w3030, IN38[19], w3122, w3123);
  FullAdder U866 (w3123, w3032, IN39[19], w3124, w3125);
  FullAdder U867 (w3125, w3034, IN40[19], w3126, w3127);
  FullAdder U868 (w3127, w3036, IN41[19], w3128, w3129);
  FullAdder U869 (w3129, w3038, IN42[19], w3130, w3131);
  FullAdder U870 (w3131, w3040, IN43[19], w3132, w3133);
  FullAdder U871 (w3133, w3042, IN44[19], w3134, w3135);
  FullAdder U872 (w3135, w3044, IN45[19], w3136, w3137);
  FullAdder U873 (w3137, w3046, IN46[19], w3138, w3139);
  FullAdder U874 (w3139, w3048, IN47[19], w3140, w3141);
  FullAdder U875 (w3141, w3050, IN48[17], w3142, w3143);
  FullAdder U876 (w3143, w3052, IN49[16], w3144, w3145);
  FullAdder U877 (w3145, w3054, IN50[15], w3146, w3147);
  FullAdder U878 (w3147, w3056, IN51[14], w3148, w3149);
  FullAdder U879 (w3149, w3058, IN52[13], w3150, w3151);
  FullAdder U880 (w3151, w3060, IN53[12], w3152, w3153);
  FullAdder U881 (w3153, w3062, IN54[11], w3154, w3155);
  FullAdder U882 (w3155, w3064, IN55[10], w3156, w3157);
  FullAdder U883 (w3157, w3066, IN56[9], w3158, w3159);
  FullAdder U884 (w3159, w3068, IN57[8], w3160, w3161);
  FullAdder U885 (w3161, w3070, IN58[7], w3162, w3163);
  FullAdder U886 (w3163, w3072, IN59[6], w3164, w3165);
  FullAdder U887 (w3165, w3074, IN60[5], w3166, w3167);
  FullAdder U888 (w3167, w3076, IN61[4], w3168, w3169);
  FullAdder U889 (w3169, w3078, IN62[3], w3170, w3171);
  FullAdder U890 (w3171, w3080, IN63[2], w3172, w3173);
  FullAdder U891 (w3173, w3082, IN64[1], w3174, w3175);
  FullAdder U892 (w3175, w3083, IN65[0], w3176, w3177);
  HalfAdder U893 (w3086, IN20[20], Out1[20], w3179);
  FullAdder U894 (w3179, w3088, IN21[20], w3180, w3181);
  FullAdder U895 (w3181, w3090, IN22[20], w3182, w3183);
  FullAdder U896 (w3183, w3092, IN23[20], w3184, w3185);
  FullAdder U897 (w3185, w3094, IN24[20], w3186, w3187);
  FullAdder U898 (w3187, w3096, IN25[20], w3188, w3189);
  FullAdder U899 (w3189, w3098, IN26[20], w3190, w3191);
  FullAdder U900 (w3191, w3100, IN27[20], w3192, w3193);
  FullAdder U901 (w3193, w3102, IN28[20], w3194, w3195);
  FullAdder U902 (w3195, w3104, IN29[20], w3196, w3197);
  FullAdder U903 (w3197, w3106, IN30[20], w3198, w3199);
  FullAdder U904 (w3199, w3108, IN31[20], w3200, w3201);
  FullAdder U905 (w3201, w3110, IN32[20], w3202, w3203);
  FullAdder U906 (w3203, w3112, IN33[20], w3204, w3205);
  FullAdder U907 (w3205, w3114, IN34[20], w3206, w3207);
  FullAdder U908 (w3207, w3116, IN35[20], w3208, w3209);
  FullAdder U909 (w3209, w3118, IN36[20], w3210, w3211);
  FullAdder U910 (w3211, w3120, IN37[20], w3212, w3213);
  FullAdder U911 (w3213, w3122, IN38[20], w3214, w3215);
  FullAdder U912 (w3215, w3124, IN39[20], w3216, w3217);
  FullAdder U913 (w3217, w3126, IN40[20], w3218, w3219);
  FullAdder U914 (w3219, w3128, IN41[20], w3220, w3221);
  FullAdder U915 (w3221, w3130, IN42[20], w3222, w3223);
  FullAdder U916 (w3223, w3132, IN43[20], w3224, w3225);
  FullAdder U917 (w3225, w3134, IN44[20], w3226, w3227);
  FullAdder U918 (w3227, w3136, IN45[20], w3228, w3229);
  FullAdder U919 (w3229, w3138, IN46[20], w3230, w3231);
  FullAdder U920 (w3231, w3140, IN47[20], w3232, w3233);
  FullAdder U921 (w3233, w3142, IN48[18], w3234, w3235);
  FullAdder U922 (w3235, w3144, IN49[17], w3236, w3237);
  FullAdder U923 (w3237, w3146, IN50[16], w3238, w3239);
  FullAdder U924 (w3239, w3148, IN51[15], w3240, w3241);
  FullAdder U925 (w3241, w3150, IN52[14], w3242, w3243);
  FullAdder U926 (w3243, w3152, IN53[13], w3244, w3245);
  FullAdder U927 (w3245, w3154, IN54[12], w3246, w3247);
  FullAdder U928 (w3247, w3156, IN55[11], w3248, w3249);
  FullAdder U929 (w3249, w3158, IN56[10], w3250, w3251);
  FullAdder U930 (w3251, w3160, IN57[9], w3252, w3253);
  FullAdder U931 (w3253, w3162, IN58[8], w3254, w3255);
  FullAdder U932 (w3255, w3164, IN59[7], w3256, w3257);
  FullAdder U933 (w3257, w3166, IN60[6], w3258, w3259);
  FullAdder U934 (w3259, w3168, IN61[5], w3260, w3261);
  FullAdder U935 (w3261, w3170, IN62[4], w3262, w3263);
  FullAdder U936 (w3263, w3172, IN63[3], w3264, w3265);
  FullAdder U937 (w3265, w3174, IN64[2], w3266, w3267);
  FullAdder U938 (w3267, w3176, IN65[1], w3268, w3269);
  FullAdder U939 (w3269, w3177, IN66[0], w3270, w3271);
  HalfAdder U940 (w3180, IN21[21], Out1[21], w3273);
  FullAdder U941 (w3273, w3182, IN22[21], w3274, w3275);
  FullAdder U942 (w3275, w3184, IN23[21], w3276, w3277);
  FullAdder U943 (w3277, w3186, IN24[21], w3278, w3279);
  FullAdder U944 (w3279, w3188, IN25[21], w3280, w3281);
  FullAdder U945 (w3281, w3190, IN26[21], w3282, w3283);
  FullAdder U946 (w3283, w3192, IN27[21], w3284, w3285);
  FullAdder U947 (w3285, w3194, IN28[21], w3286, w3287);
  FullAdder U948 (w3287, w3196, IN29[21], w3288, w3289);
  FullAdder U949 (w3289, w3198, IN30[21], w3290, w3291);
  FullAdder U950 (w3291, w3200, IN31[21], w3292, w3293);
  FullAdder U951 (w3293, w3202, IN32[21], w3294, w3295);
  FullAdder U952 (w3295, w3204, IN33[21], w3296, w3297);
  FullAdder U953 (w3297, w3206, IN34[21], w3298, w3299);
  FullAdder U954 (w3299, w3208, IN35[21], w3300, w3301);
  FullAdder U955 (w3301, w3210, IN36[21], w3302, w3303);
  FullAdder U956 (w3303, w3212, IN37[21], w3304, w3305);
  FullAdder U957 (w3305, w3214, IN38[21], w3306, w3307);
  FullAdder U958 (w3307, w3216, IN39[21], w3308, w3309);
  FullAdder U959 (w3309, w3218, IN40[21], w3310, w3311);
  FullAdder U960 (w3311, w3220, IN41[21], w3312, w3313);
  FullAdder U961 (w3313, w3222, IN42[21], w3314, w3315);
  FullAdder U962 (w3315, w3224, IN43[21], w3316, w3317);
  FullAdder U963 (w3317, w3226, IN44[21], w3318, w3319);
  FullAdder U964 (w3319, w3228, IN45[21], w3320, w3321);
  FullAdder U965 (w3321, w3230, IN46[21], w3322, w3323);
  FullAdder U966 (w3323, w3232, IN47[21], w3324, w3325);
  FullAdder U967 (w3325, w3234, IN48[19], w3326, w3327);
  FullAdder U968 (w3327, w3236, IN49[18], w3328, w3329);
  FullAdder U969 (w3329, w3238, IN50[17], w3330, w3331);
  FullAdder U970 (w3331, w3240, IN51[16], w3332, w3333);
  FullAdder U971 (w3333, w3242, IN52[15], w3334, w3335);
  FullAdder U972 (w3335, w3244, IN53[14], w3336, w3337);
  FullAdder U973 (w3337, w3246, IN54[13], w3338, w3339);
  FullAdder U974 (w3339, w3248, IN55[12], w3340, w3341);
  FullAdder U975 (w3341, w3250, IN56[11], w3342, w3343);
  FullAdder U976 (w3343, w3252, IN57[10], w3344, w3345);
  FullAdder U977 (w3345, w3254, IN58[9], w3346, w3347);
  FullAdder U978 (w3347, w3256, IN59[8], w3348, w3349);
  FullAdder U979 (w3349, w3258, IN60[7], w3350, w3351);
  FullAdder U980 (w3351, w3260, IN61[6], w3352, w3353);
  FullAdder U981 (w3353, w3262, IN62[5], w3354, w3355);
  FullAdder U982 (w3355, w3264, IN63[4], w3356, w3357);
  FullAdder U983 (w3357, w3266, IN64[3], w3358, w3359);
  FullAdder U984 (w3359, w3268, IN65[2], w3360, w3361);
  FullAdder U985 (w3361, w3270, IN66[1], w3362, w3363);
  FullAdder U986 (w3363, w3271, IN67[0], w3364, w3365);
  HalfAdder U987 (w3274, IN22[22], Out1[22], w3367);
  FullAdder U988 (w3367, w3276, IN23[22], w3368, w3369);
  FullAdder U989 (w3369, w3278, IN24[22], w3370, w3371);
  FullAdder U990 (w3371, w3280, IN25[22], w3372, w3373);
  FullAdder U991 (w3373, w3282, IN26[22], w3374, w3375);
  FullAdder U992 (w3375, w3284, IN27[22], w3376, w3377);
  FullAdder U993 (w3377, w3286, IN28[22], w3378, w3379);
  FullAdder U994 (w3379, w3288, IN29[22], w3380, w3381);
  FullAdder U995 (w3381, w3290, IN30[22], w3382, w3383);
  FullAdder U996 (w3383, w3292, IN31[22], w3384, w3385);
  FullAdder U997 (w3385, w3294, IN32[22], w3386, w3387);
  FullAdder U998 (w3387, w3296, IN33[22], w3388, w3389);
  FullAdder U999 (w3389, w3298, IN34[22], w3390, w3391);
  FullAdder U1000 (w3391, w3300, IN35[22], w3392, w3393);
  FullAdder U1001 (w3393, w3302, IN36[22], w3394, w3395);
  FullAdder U1002 (w3395, w3304, IN37[22], w3396, w3397);
  FullAdder U1003 (w3397, w3306, IN38[22], w3398, w3399);
  FullAdder U1004 (w3399, w3308, IN39[22], w3400, w3401);
  FullAdder U1005 (w3401, w3310, IN40[22], w3402, w3403);
  FullAdder U1006 (w3403, w3312, IN41[22], w3404, w3405);
  FullAdder U1007 (w3405, w3314, IN42[22], w3406, w3407);
  FullAdder U1008 (w3407, w3316, IN43[22], w3408, w3409);
  FullAdder U1009 (w3409, w3318, IN44[22], w3410, w3411);
  FullAdder U1010 (w3411, w3320, IN45[22], w3412, w3413);
  FullAdder U1011 (w3413, w3322, IN46[22], w3414, w3415);
  FullAdder U1012 (w3415, w3324, IN47[22], w3416, w3417);
  FullAdder U1013 (w3417, w3326, IN48[20], w3418, w3419);
  FullAdder U1014 (w3419, w3328, IN49[19], w3420, w3421);
  FullAdder U1015 (w3421, w3330, IN50[18], w3422, w3423);
  FullAdder U1016 (w3423, w3332, IN51[17], w3424, w3425);
  FullAdder U1017 (w3425, w3334, IN52[16], w3426, w3427);
  FullAdder U1018 (w3427, w3336, IN53[15], w3428, w3429);
  FullAdder U1019 (w3429, w3338, IN54[14], w3430, w3431);
  FullAdder U1020 (w3431, w3340, IN55[13], w3432, w3433);
  FullAdder U1021 (w3433, w3342, IN56[12], w3434, w3435);
  FullAdder U1022 (w3435, w3344, IN57[11], w3436, w3437);
  FullAdder U1023 (w3437, w3346, IN58[10], w3438, w3439);
  FullAdder U1024 (w3439, w3348, IN59[9], w3440, w3441);
  FullAdder U1025 (w3441, w3350, IN60[8], w3442, w3443);
  FullAdder U1026 (w3443, w3352, IN61[7], w3444, w3445);
  FullAdder U1027 (w3445, w3354, IN62[6], w3446, w3447);
  FullAdder U1028 (w3447, w3356, IN63[5], w3448, w3449);
  FullAdder U1029 (w3449, w3358, IN64[4], w3450, w3451);
  FullAdder U1030 (w3451, w3360, IN65[3], w3452, w3453);
  FullAdder U1031 (w3453, w3362, IN66[2], w3454, w3455);
  FullAdder U1032 (w3455, w3364, IN67[1], w3456, w3457);
  FullAdder U1033 (w3457, w3365, IN68[0], w3458, w3459);
  HalfAdder U1034 (w3368, IN23[23], Out1[23], w3461);
  FullAdder U1035 (w3461, w3370, IN24[23], w3462, w3463);
  FullAdder U1036 (w3463, w3372, IN25[23], w3464, w3465);
  FullAdder U1037 (w3465, w3374, IN26[23], w3466, w3467);
  FullAdder U1038 (w3467, w3376, IN27[23], w3468, w3469);
  FullAdder U1039 (w3469, w3378, IN28[23], w3470, w3471);
  FullAdder U1040 (w3471, w3380, IN29[23], w3472, w3473);
  FullAdder U1041 (w3473, w3382, IN30[23], w3474, w3475);
  FullAdder U1042 (w3475, w3384, IN31[23], w3476, w3477);
  FullAdder U1043 (w3477, w3386, IN32[23], w3478, w3479);
  FullAdder U1044 (w3479, w3388, IN33[23], w3480, w3481);
  FullAdder U1045 (w3481, w3390, IN34[23], w3482, w3483);
  FullAdder U1046 (w3483, w3392, IN35[23], w3484, w3485);
  FullAdder U1047 (w3485, w3394, IN36[23], w3486, w3487);
  FullAdder U1048 (w3487, w3396, IN37[23], w3488, w3489);
  FullAdder U1049 (w3489, w3398, IN38[23], w3490, w3491);
  FullAdder U1050 (w3491, w3400, IN39[23], w3492, w3493);
  FullAdder U1051 (w3493, w3402, IN40[23], w3494, w3495);
  FullAdder U1052 (w3495, w3404, IN41[23], w3496, w3497);
  FullAdder U1053 (w3497, w3406, IN42[23], w3498, w3499);
  FullAdder U1054 (w3499, w3408, IN43[23], w3500, w3501);
  FullAdder U1055 (w3501, w3410, IN44[23], w3502, w3503);
  FullAdder U1056 (w3503, w3412, IN45[23], w3504, w3505);
  FullAdder U1057 (w3505, w3414, IN46[23], w3506, w3507);
  FullAdder U1058 (w3507, w3416, IN47[23], w3508, w3509);
  FullAdder U1059 (w3509, w3418, IN48[21], w3510, w3511);
  FullAdder U1060 (w3511, w3420, IN49[20], w3512, w3513);
  FullAdder U1061 (w3513, w3422, IN50[19], w3514, w3515);
  FullAdder U1062 (w3515, w3424, IN51[18], w3516, w3517);
  FullAdder U1063 (w3517, w3426, IN52[17], w3518, w3519);
  FullAdder U1064 (w3519, w3428, IN53[16], w3520, w3521);
  FullAdder U1065 (w3521, w3430, IN54[15], w3522, w3523);
  FullAdder U1066 (w3523, w3432, IN55[14], w3524, w3525);
  FullAdder U1067 (w3525, w3434, IN56[13], w3526, w3527);
  FullAdder U1068 (w3527, w3436, IN57[12], w3528, w3529);
  FullAdder U1069 (w3529, w3438, IN58[11], w3530, w3531);
  FullAdder U1070 (w3531, w3440, IN59[10], w3532, w3533);
  FullAdder U1071 (w3533, w3442, IN60[9], w3534, w3535);
  FullAdder U1072 (w3535, w3444, IN61[8], w3536, w3537);
  FullAdder U1073 (w3537, w3446, IN62[7], w3538, w3539);
  FullAdder U1074 (w3539, w3448, IN63[6], w3540, w3541);
  FullAdder U1075 (w3541, w3450, IN64[5], w3542, w3543);
  FullAdder U1076 (w3543, w3452, IN65[4], w3544, w3545);
  FullAdder U1077 (w3545, w3454, IN66[3], w3546, w3547);
  FullAdder U1078 (w3547, w3456, IN67[2], w3548, w3549);
  FullAdder U1079 (w3549, w3458, IN68[1], w3550, w3551);
  FullAdder U1080 (w3551, w3459, IN69[0], w3552, w3553);
  HalfAdder U1081 (w3462, IN24[24], Out1[24], w3555);
  FullAdder U1082 (w3555, w3464, IN25[24], w3556, w3557);
  FullAdder U1083 (w3557, w3466, IN26[24], w3558, w3559);
  FullAdder U1084 (w3559, w3468, IN27[24], w3560, w3561);
  FullAdder U1085 (w3561, w3470, IN28[24], w3562, w3563);
  FullAdder U1086 (w3563, w3472, IN29[24], w3564, w3565);
  FullAdder U1087 (w3565, w3474, IN30[24], w3566, w3567);
  FullAdder U1088 (w3567, w3476, IN31[24], w3568, w3569);
  FullAdder U1089 (w3569, w3478, IN32[24], w3570, w3571);
  FullAdder U1090 (w3571, w3480, IN33[24], w3572, w3573);
  FullAdder U1091 (w3573, w3482, IN34[24], w3574, w3575);
  FullAdder U1092 (w3575, w3484, IN35[24], w3576, w3577);
  FullAdder U1093 (w3577, w3486, IN36[24], w3578, w3579);
  FullAdder U1094 (w3579, w3488, IN37[24], w3580, w3581);
  FullAdder U1095 (w3581, w3490, IN38[24], w3582, w3583);
  FullAdder U1096 (w3583, w3492, IN39[24], w3584, w3585);
  FullAdder U1097 (w3585, w3494, IN40[24], w3586, w3587);
  FullAdder U1098 (w3587, w3496, IN41[24], w3588, w3589);
  FullAdder U1099 (w3589, w3498, IN42[24], w3590, w3591);
  FullAdder U1100 (w3591, w3500, IN43[24], w3592, w3593);
  FullAdder U1101 (w3593, w3502, IN44[24], w3594, w3595);
  FullAdder U1102 (w3595, w3504, IN45[24], w3596, w3597);
  FullAdder U1103 (w3597, w3506, IN46[24], w3598, w3599);
  FullAdder U1104 (w3599, w3508, IN47[24], w3600, w3601);
  FullAdder U1105 (w3601, w3510, IN48[22], w3602, w3603);
  FullAdder U1106 (w3603, w3512, IN49[21], w3604, w3605);
  FullAdder U1107 (w3605, w3514, IN50[20], w3606, w3607);
  FullAdder U1108 (w3607, w3516, IN51[19], w3608, w3609);
  FullAdder U1109 (w3609, w3518, IN52[18], w3610, w3611);
  FullAdder U1110 (w3611, w3520, IN53[17], w3612, w3613);
  FullAdder U1111 (w3613, w3522, IN54[16], w3614, w3615);
  FullAdder U1112 (w3615, w3524, IN55[15], w3616, w3617);
  FullAdder U1113 (w3617, w3526, IN56[14], w3618, w3619);
  FullAdder U1114 (w3619, w3528, IN57[13], w3620, w3621);
  FullAdder U1115 (w3621, w3530, IN58[12], w3622, w3623);
  FullAdder U1116 (w3623, w3532, IN59[11], w3624, w3625);
  FullAdder U1117 (w3625, w3534, IN60[10], w3626, w3627);
  FullAdder U1118 (w3627, w3536, IN61[9], w3628, w3629);
  FullAdder U1119 (w3629, w3538, IN62[8], w3630, w3631);
  FullAdder U1120 (w3631, w3540, IN63[7], w3632, w3633);
  FullAdder U1121 (w3633, w3542, IN64[6], w3634, w3635);
  FullAdder U1122 (w3635, w3544, IN65[5], w3636, w3637);
  FullAdder U1123 (w3637, w3546, IN66[4], w3638, w3639);
  FullAdder U1124 (w3639, w3548, IN67[3], w3640, w3641);
  FullAdder U1125 (w3641, w3550, IN68[2], w3642, w3643);
  FullAdder U1126 (w3643, w3552, IN69[1], w3644, w3645);
  FullAdder U1127 (w3645, w3553, IN70[0], w3646, w3647);
  HalfAdder U1128 (w3556, IN25[25], Out1[25], w3649);
  FullAdder U1129 (w3649, w3558, IN26[25], w3650, w3651);
  FullAdder U1130 (w3651, w3560, IN27[25], w3652, w3653);
  FullAdder U1131 (w3653, w3562, IN28[25], w3654, w3655);
  FullAdder U1132 (w3655, w3564, IN29[25], w3656, w3657);
  FullAdder U1133 (w3657, w3566, IN30[25], w3658, w3659);
  FullAdder U1134 (w3659, w3568, IN31[25], w3660, w3661);
  FullAdder U1135 (w3661, w3570, IN32[25], w3662, w3663);
  FullAdder U1136 (w3663, w3572, IN33[25], w3664, w3665);
  FullAdder U1137 (w3665, w3574, IN34[25], w3666, w3667);
  FullAdder U1138 (w3667, w3576, IN35[25], w3668, w3669);
  FullAdder U1139 (w3669, w3578, IN36[25], w3670, w3671);
  FullAdder U1140 (w3671, w3580, IN37[25], w3672, w3673);
  FullAdder U1141 (w3673, w3582, IN38[25], w3674, w3675);
  FullAdder U1142 (w3675, w3584, IN39[25], w3676, w3677);
  FullAdder U1143 (w3677, w3586, IN40[25], w3678, w3679);
  FullAdder U1144 (w3679, w3588, IN41[25], w3680, w3681);
  FullAdder U1145 (w3681, w3590, IN42[25], w3682, w3683);
  FullAdder U1146 (w3683, w3592, IN43[25], w3684, w3685);
  FullAdder U1147 (w3685, w3594, IN44[25], w3686, w3687);
  FullAdder U1148 (w3687, w3596, IN45[25], w3688, w3689);
  FullAdder U1149 (w3689, w3598, IN46[25], w3690, w3691);
  FullAdder U1150 (w3691, w3600, IN47[25], w3692, w3693);
  FullAdder U1151 (w3693, w3602, IN48[23], w3694, w3695);
  FullAdder U1152 (w3695, w3604, IN49[22], w3696, w3697);
  FullAdder U1153 (w3697, w3606, IN50[21], w3698, w3699);
  FullAdder U1154 (w3699, w3608, IN51[20], w3700, w3701);
  FullAdder U1155 (w3701, w3610, IN52[19], w3702, w3703);
  FullAdder U1156 (w3703, w3612, IN53[18], w3704, w3705);
  FullAdder U1157 (w3705, w3614, IN54[17], w3706, w3707);
  FullAdder U1158 (w3707, w3616, IN55[16], w3708, w3709);
  FullAdder U1159 (w3709, w3618, IN56[15], w3710, w3711);
  FullAdder U1160 (w3711, w3620, IN57[14], w3712, w3713);
  FullAdder U1161 (w3713, w3622, IN58[13], w3714, w3715);
  FullAdder U1162 (w3715, w3624, IN59[12], w3716, w3717);
  FullAdder U1163 (w3717, w3626, IN60[11], w3718, w3719);
  FullAdder U1164 (w3719, w3628, IN61[10], w3720, w3721);
  FullAdder U1165 (w3721, w3630, IN62[9], w3722, w3723);
  FullAdder U1166 (w3723, w3632, IN63[8], w3724, w3725);
  FullAdder U1167 (w3725, w3634, IN64[7], w3726, w3727);
  FullAdder U1168 (w3727, w3636, IN65[6], w3728, w3729);
  FullAdder U1169 (w3729, w3638, IN66[5], w3730, w3731);
  FullAdder U1170 (w3731, w3640, IN67[4], w3732, w3733);
  FullAdder U1171 (w3733, w3642, IN68[3], w3734, w3735);
  FullAdder U1172 (w3735, w3644, IN69[2], w3736, w3737);
  FullAdder U1173 (w3737, w3646, IN70[1], w3738, w3739);
  FullAdder U1174 (w3739, w3647, IN71[0], w3740, w3741);
  HalfAdder U1175 (w3650, IN26[26], Out1[26], w3743);
  FullAdder U1176 (w3743, w3652, IN27[26], w3744, w3745);
  FullAdder U1177 (w3745, w3654, IN28[26], w3746, w3747);
  FullAdder U1178 (w3747, w3656, IN29[26], w3748, w3749);
  FullAdder U1179 (w3749, w3658, IN30[26], w3750, w3751);
  FullAdder U1180 (w3751, w3660, IN31[26], w3752, w3753);
  FullAdder U1181 (w3753, w3662, IN32[26], w3754, w3755);
  FullAdder U1182 (w3755, w3664, IN33[26], w3756, w3757);
  FullAdder U1183 (w3757, w3666, IN34[26], w3758, w3759);
  FullAdder U1184 (w3759, w3668, IN35[26], w3760, w3761);
  FullAdder U1185 (w3761, w3670, IN36[26], w3762, w3763);
  FullAdder U1186 (w3763, w3672, IN37[26], w3764, w3765);
  FullAdder U1187 (w3765, w3674, IN38[26], w3766, w3767);
  FullAdder U1188 (w3767, w3676, IN39[26], w3768, w3769);
  FullAdder U1189 (w3769, w3678, IN40[26], w3770, w3771);
  FullAdder U1190 (w3771, w3680, IN41[26], w3772, w3773);
  FullAdder U1191 (w3773, w3682, IN42[26], w3774, w3775);
  FullAdder U1192 (w3775, w3684, IN43[26], w3776, w3777);
  FullAdder U1193 (w3777, w3686, IN44[26], w3778, w3779);
  FullAdder U1194 (w3779, w3688, IN45[26], w3780, w3781);
  FullAdder U1195 (w3781, w3690, IN46[26], w3782, w3783);
  FullAdder U1196 (w3783, w3692, IN47[26], w3784, w3785);
  FullAdder U1197 (w3785, w3694, IN48[24], w3786, w3787);
  FullAdder U1198 (w3787, w3696, IN49[23], w3788, w3789);
  FullAdder U1199 (w3789, w3698, IN50[22], w3790, w3791);
  FullAdder U1200 (w3791, w3700, IN51[21], w3792, w3793);
  FullAdder U1201 (w3793, w3702, IN52[20], w3794, w3795);
  FullAdder U1202 (w3795, w3704, IN53[19], w3796, w3797);
  FullAdder U1203 (w3797, w3706, IN54[18], w3798, w3799);
  FullAdder U1204 (w3799, w3708, IN55[17], w3800, w3801);
  FullAdder U1205 (w3801, w3710, IN56[16], w3802, w3803);
  FullAdder U1206 (w3803, w3712, IN57[15], w3804, w3805);
  FullAdder U1207 (w3805, w3714, IN58[14], w3806, w3807);
  FullAdder U1208 (w3807, w3716, IN59[13], w3808, w3809);
  FullAdder U1209 (w3809, w3718, IN60[12], w3810, w3811);
  FullAdder U1210 (w3811, w3720, IN61[11], w3812, w3813);
  FullAdder U1211 (w3813, w3722, IN62[10], w3814, w3815);
  FullAdder U1212 (w3815, w3724, IN63[9], w3816, w3817);
  FullAdder U1213 (w3817, w3726, IN64[8], w3818, w3819);
  FullAdder U1214 (w3819, w3728, IN65[7], w3820, w3821);
  FullAdder U1215 (w3821, w3730, IN66[6], w3822, w3823);
  FullAdder U1216 (w3823, w3732, IN67[5], w3824, w3825);
  FullAdder U1217 (w3825, w3734, IN68[4], w3826, w3827);
  FullAdder U1218 (w3827, w3736, IN69[3], w3828, w3829);
  FullAdder U1219 (w3829, w3738, IN70[2], w3830, w3831);
  FullAdder U1220 (w3831, w3740, IN71[1], w3832, w3833);
  FullAdder U1221 (w3833, w3741, IN72[0], w3834, w3835);
  HalfAdder U1222 (w3744, IN27[27], Out1[27], w3837);
  FullAdder U1223 (w3837, w3746, IN28[27], w3838, w3839);
  FullAdder U1224 (w3839, w3748, IN29[27], w3840, w3841);
  FullAdder U1225 (w3841, w3750, IN30[27], w3842, w3843);
  FullAdder U1226 (w3843, w3752, IN31[27], w3844, w3845);
  FullAdder U1227 (w3845, w3754, IN32[27], w3846, w3847);
  FullAdder U1228 (w3847, w3756, IN33[27], w3848, w3849);
  FullAdder U1229 (w3849, w3758, IN34[27], w3850, w3851);
  FullAdder U1230 (w3851, w3760, IN35[27], w3852, w3853);
  FullAdder U1231 (w3853, w3762, IN36[27], w3854, w3855);
  FullAdder U1232 (w3855, w3764, IN37[27], w3856, w3857);
  FullAdder U1233 (w3857, w3766, IN38[27], w3858, w3859);
  FullAdder U1234 (w3859, w3768, IN39[27], w3860, w3861);
  FullAdder U1235 (w3861, w3770, IN40[27], w3862, w3863);
  FullAdder U1236 (w3863, w3772, IN41[27], w3864, w3865);
  FullAdder U1237 (w3865, w3774, IN42[27], w3866, w3867);
  FullAdder U1238 (w3867, w3776, IN43[27], w3868, w3869);
  FullAdder U1239 (w3869, w3778, IN44[27], w3870, w3871);
  FullAdder U1240 (w3871, w3780, IN45[27], w3872, w3873);
  FullAdder U1241 (w3873, w3782, IN46[27], w3874, w3875);
  FullAdder U1242 (w3875, w3784, IN47[27], w3876, w3877);
  FullAdder U1243 (w3877, w3786, IN48[25], w3878, w3879);
  FullAdder U1244 (w3879, w3788, IN49[24], w3880, w3881);
  FullAdder U1245 (w3881, w3790, IN50[23], w3882, w3883);
  FullAdder U1246 (w3883, w3792, IN51[22], w3884, w3885);
  FullAdder U1247 (w3885, w3794, IN52[21], w3886, w3887);
  FullAdder U1248 (w3887, w3796, IN53[20], w3888, w3889);
  FullAdder U1249 (w3889, w3798, IN54[19], w3890, w3891);
  FullAdder U1250 (w3891, w3800, IN55[18], w3892, w3893);
  FullAdder U1251 (w3893, w3802, IN56[17], w3894, w3895);
  FullAdder U1252 (w3895, w3804, IN57[16], w3896, w3897);
  FullAdder U1253 (w3897, w3806, IN58[15], w3898, w3899);
  FullAdder U1254 (w3899, w3808, IN59[14], w3900, w3901);
  FullAdder U1255 (w3901, w3810, IN60[13], w3902, w3903);
  FullAdder U1256 (w3903, w3812, IN61[12], w3904, w3905);
  FullAdder U1257 (w3905, w3814, IN62[11], w3906, w3907);
  FullAdder U1258 (w3907, w3816, IN63[10], w3908, w3909);
  FullAdder U1259 (w3909, w3818, IN64[9], w3910, w3911);
  FullAdder U1260 (w3911, w3820, IN65[8], w3912, w3913);
  FullAdder U1261 (w3913, w3822, IN66[7], w3914, w3915);
  FullAdder U1262 (w3915, w3824, IN67[6], w3916, w3917);
  FullAdder U1263 (w3917, w3826, IN68[5], w3918, w3919);
  FullAdder U1264 (w3919, w3828, IN69[4], w3920, w3921);
  FullAdder U1265 (w3921, w3830, IN70[3], w3922, w3923);
  FullAdder U1266 (w3923, w3832, IN71[2], w3924, w3925);
  FullAdder U1267 (w3925, w3834, IN72[1], w3926, w3927);
  FullAdder U1268 (w3927, w3835, IN73[0], w3928, w3929);
  HalfAdder U1269 (w3838, IN28[28], Out1[28], w3931);
  FullAdder U1270 (w3931, w3840, IN29[28], Out1[29], w3933);
  FullAdder U1271 (w3933, w3842, IN30[28], Out1[30], w3935);
  FullAdder U1272 (w3935, w3844, IN31[28], Out1[31], w3937);
  FullAdder U1273 (w3937, w3846, IN32[28], Out1[32], w3939);
  FullAdder U1274 (w3939, w3848, IN33[28], Out1[33], w3941);
  FullAdder U1275 (w3941, w3850, IN34[28], Out1[34], w3943);
  FullAdder U1276 (w3943, w3852, IN35[28], Out1[35], w3945);
  FullAdder U1277 (w3945, w3854, IN36[28], Out1[36], w3947);
  FullAdder U1278 (w3947, w3856, IN37[28], Out1[37], w3949);
  FullAdder U1279 (w3949, w3858, IN38[28], Out1[38], w3951);
  FullAdder U1280 (w3951, w3860, IN39[28], Out1[39], w3953);
  FullAdder U1281 (w3953, w3862, IN40[28], Out1[40], w3955);
  FullAdder U1282 (w3955, w3864, IN41[28], Out1[41], w3957);
  FullAdder U1283 (w3957, w3866, IN42[28], Out1[42], w3959);
  FullAdder U1284 (w3959, w3868, IN43[28], Out1[43], w3961);
  FullAdder U1285 (w3961, w3870, IN44[28], Out1[44], w3963);
  FullAdder U1286 (w3963, w3872, IN45[28], Out1[45], w3965);
  FullAdder U1287 (w3965, w3874, IN46[28], Out1[46], w3967);
  FullAdder U1288 (w3967, w3876, IN47[28], Out1[47], w3969);
  FullAdder U1289 (w3969, w3878, IN48[26], Out1[48], w3971);
  FullAdder U1290 (w3971, w3880, IN49[25], Out1[49], w3973);
  FullAdder U1291 (w3973, w3882, IN50[24], Out1[50], w3975);
  FullAdder U1292 (w3975, w3884, IN51[23], Out1[51], w3977);
  FullAdder U1293 (w3977, w3886, IN52[22], Out1[52], w3979);
  FullAdder U1294 (w3979, w3888, IN53[21], Out1[53], w3981);
  FullAdder U1295 (w3981, w3890, IN54[20], Out1[54], w3983);
  FullAdder U1296 (w3983, w3892, IN55[19], Out1[55], w3985);
  FullAdder U1297 (w3985, w3894, IN56[18], Out1[56], w3987);
  FullAdder U1298 (w3987, w3896, IN57[17], Out1[57], w3989);
  FullAdder U1299 (w3989, w3898, IN58[16], Out1[58], w3991);
  FullAdder U1300 (w3991, w3900, IN59[15], Out1[59], w3993);
  FullAdder U1301 (w3993, w3902, IN60[14], Out1[60], w3995);
  FullAdder U1302 (w3995, w3904, IN61[13], Out1[61], w3997);
  FullAdder U1303 (w3997, w3906, IN62[12], Out1[62], w3999);
  FullAdder U1304 (w3999, w3908, IN63[11], Out1[63], w4001);
  FullAdder U1305 (w4001, w3910, IN64[10], Out1[64], w4003);
  FullAdder U1306 (w4003, w3912, IN65[9], Out1[65], w4005);
  FullAdder U1307 (w4005, w3914, IN66[8], Out1[66], w4007);
  FullAdder U1308 (w4007, w3916, IN67[7], Out1[67], w4009);
  FullAdder U1309 (w4009, w3918, IN68[6], Out1[68], w4011);
  FullAdder U1310 (w4011, w3920, IN69[5], Out1[69], w4013);
  FullAdder U1311 (w4013, w3922, IN70[4], Out1[70], w4015);
  FullAdder U1312 (w4015, w3924, IN71[3], Out1[71], w4017);
  FullAdder U1313 (w4017, w3926, IN72[2], Out1[72], w4019);
  FullAdder U1314 (w4019, w3928, IN73[1], Out1[73], w4021);
  FullAdder U1315 (w4021, w3929, IN74[0], Out1[74], Out1[75]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN48[27];
  assign Out2[1] = IN49[26];
  assign Out2[2] = IN50[25];
  assign Out2[3] = IN51[24];
  assign Out2[4] = IN52[23];
  assign Out2[5] = IN53[22];
  assign Out2[6] = IN54[21];
  assign Out2[7] = IN55[20];
  assign Out2[8] = IN56[19];
  assign Out2[9] = IN57[18];
  assign Out2[10] = IN58[17];
  assign Out2[11] = IN59[16];
  assign Out2[12] = IN60[15];
  assign Out2[13] = IN61[14];
  assign Out2[14] = IN62[13];
  assign Out2[15] = IN63[12];
  assign Out2[16] = IN64[11];
  assign Out2[17] = IN65[10];
  assign Out2[18] = IN66[9];
  assign Out2[19] = IN67[8];
  assign Out2[20] = IN68[7];
  assign Out2[21] = IN69[6];
  assign Out2[22] = IN70[5];
  assign Out2[23] = IN71[4];
  assign Out2[24] = IN72[3];
  assign Out2[25] = IN73[2];
  assign Out2[26] = IN74[1];
  assign Out2[27] = IN75[0];

endmodule
module RC_28_28(IN1, IN2, Out);
  input [27:0] IN1;
  input [27:0] IN2;
  output [28:0] Out;
  wire w57;
  wire w59;
  wire w61;
  wire w63;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w57);
  FullAdder U1 (IN1[1], IN2[1], w57, Out[1], w59);
  FullAdder U2 (IN1[2], IN2[2], w59, Out[2], w61);
  FullAdder U3 (IN1[3], IN2[3], w61, Out[3], w63);
  FullAdder U4 (IN1[4], IN2[4], w63, Out[4], w65);
  FullAdder U5 (IN1[5], IN2[5], w65, Out[5], w67);
  FullAdder U6 (IN1[6], IN2[6], w67, Out[6], w69);
  FullAdder U7 (IN1[7], IN2[7], w69, Out[7], w71);
  FullAdder U8 (IN1[8], IN2[8], w71, Out[8], w73);
  FullAdder U9 (IN1[9], IN2[9], w73, Out[9], w75);
  FullAdder U10 (IN1[10], IN2[10], w75, Out[10], w77);
  FullAdder U11 (IN1[11], IN2[11], w77, Out[11], w79);
  FullAdder U12 (IN1[12], IN2[12], w79, Out[12], w81);
  FullAdder U13 (IN1[13], IN2[13], w81, Out[13], w83);
  FullAdder U14 (IN1[14], IN2[14], w83, Out[14], w85);
  FullAdder U15 (IN1[15], IN2[15], w85, Out[15], w87);
  FullAdder U16 (IN1[16], IN2[16], w87, Out[16], w89);
  FullAdder U17 (IN1[17], IN2[17], w89, Out[17], w91);
  FullAdder U18 (IN1[18], IN2[18], w91, Out[18], w93);
  FullAdder U19 (IN1[19], IN2[19], w93, Out[19], w95);
  FullAdder U20 (IN1[20], IN2[20], w95, Out[20], w97);
  FullAdder U21 (IN1[21], IN2[21], w97, Out[21], w99);
  FullAdder U22 (IN1[22], IN2[22], w99, Out[22], w101);
  FullAdder U23 (IN1[23], IN2[23], w101, Out[23], w103);
  FullAdder U24 (IN1[24], IN2[24], w103, Out[24], w105);
  FullAdder U25 (IN1[25], IN2[25], w105, Out[25], w107);
  FullAdder U26 (IN1[26], IN2[26], w107, Out[26], w109);
  FullAdder U27 (IN1[27], IN2[27], w109, Out[27], Out[28]);

endmodule
module NR_48_29(IN1, IN2, Out);
  input [47:0] IN1;
  input [28:0] IN2;
  output [76:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [28:0] P29;
  wire [28:0] P30;
  wire [28:0] P31;
  wire [28:0] P32;
  wire [28:0] P33;
  wire [28:0] P34;
  wire [28:0] P35;
  wire [28:0] P36;
  wire [28:0] P37;
  wire [28:0] P38;
  wire [28:0] P39;
  wire [28:0] P40;
  wire [28:0] P41;
  wire [28:0] P42;
  wire [28:0] P43;
  wire [28:0] P44;
  wire [28:0] P45;
  wire [28:0] P46;
  wire [28:0] P47;
  wire [27:0] P48;
  wire [26:0] P49;
  wire [25:0] P50;
  wire [24:0] P51;
  wire [23:0] P52;
  wire [22:0] P53;
  wire [21:0] P54;
  wire [20:0] P55;
  wire [19:0] P56;
  wire [18:0] P57;
  wire [17:0] P58;
  wire [16:0] P59;
  wire [15:0] P60;
  wire [14:0] P61;
  wire [13:0] P62;
  wire [12:0] P63;
  wire [11:0] P64;
  wire [10:0] P65;
  wire [9:0] P66;
  wire [8:0] P67;
  wire [7:0] P68;
  wire [6:0] P69;
  wire [5:0] P70;
  wire [4:0] P71;
  wire [3:0] P72;
  wire [2:0] P73;
  wire [1:0] P74;
  wire [0:0] P75;
  wire [75:0] R1;
  wire [27:0] R2;
  wire [76:0] aOut;
  U_SP_48_29 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, R1, R2);
  RC_28_28 S2 (R1[75:48], R2, aOut[76:48]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign Out = aOut[76:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
