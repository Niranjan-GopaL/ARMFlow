//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 7
  second input length: 60
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_7_60(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65);
  input [6:0] IN1;
  input [59:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [6:0] P37;
  output [6:0] P38;
  output [6:0] P39;
  output [6:0] P40;
  output [6:0] P41;
  output [6:0] P42;
  output [6:0] P43;
  output [6:0] P44;
  output [6:0] P45;
  output [6:0] P46;
  output [6:0] P47;
  output [6:0] P48;
  output [6:0] P49;
  output [6:0] P50;
  output [6:0] P51;
  output [6:0] P52;
  output [6:0] P53;
  output [6:0] P54;
  output [6:0] P55;
  output [6:0] P56;
  output [6:0] P57;
  output [6:0] P58;
  output [6:0] P59;
  output [5:0] P60;
  output [4:0] P61;
  output [3:0] P62;
  output [2:0] P63;
  output [1:0] P64;
  output [0:0] P65;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P59[0] = IN1[0]&IN2[59];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[1] = IN1[1]&IN2[58];
  assign P60[0] = IN1[1]&IN2[59];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[2] = IN1[2]&IN2[57];
  assign P60[1] = IN1[2]&IN2[58];
  assign P61[0] = IN1[2]&IN2[59];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[3] = IN1[3]&IN2[56];
  assign P60[2] = IN1[3]&IN2[57];
  assign P61[1] = IN1[3]&IN2[58];
  assign P62[0] = IN1[3]&IN2[59];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[4] = IN1[4]&IN2[55];
  assign P60[3] = IN1[4]&IN2[56];
  assign P61[2] = IN1[4]&IN2[57];
  assign P62[1] = IN1[4]&IN2[58];
  assign P63[0] = IN1[4]&IN2[59];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[5] = IN1[5]&IN2[54];
  assign P60[4] = IN1[5]&IN2[55];
  assign P61[3] = IN1[5]&IN2[56];
  assign P62[2] = IN1[5]&IN2[57];
  assign P63[1] = IN1[5]&IN2[58];
  assign P64[0] = IN1[5]&IN2[59];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[6] = IN1[6]&IN2[53];
  assign P60[5] = IN1[6]&IN2[54];
  assign P61[4] = IN1[6]&IN2[55];
  assign P62[3] = IN1[6]&IN2[56];
  assign P63[2] = IN1[6]&IN2[57];
  assign P64[1] = IN1[6]&IN2[58];
  assign P65[0] = IN1[6]&IN2[59];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [6:0] IN37;
  input [6:0] IN38;
  input [6:0] IN39;
  input [6:0] IN40;
  input [6:0] IN41;
  input [6:0] IN42;
  input [6:0] IN43;
  input [6:0] IN44;
  input [6:0] IN45;
  input [6:0] IN46;
  input [6:0] IN47;
  input [6:0] IN48;
  input [6:0] IN49;
  input [6:0] IN50;
  input [6:0] IN51;
  input [6:0] IN52;
  input [6:0] IN53;
  input [6:0] IN54;
  input [6:0] IN55;
  input [6:0] IN56;
  input [6:0] IN57;
  input [6:0] IN58;
  input [6:0] IN59;
  input [5:0] IN60;
  input [4:0] IN61;
  input [3:0] IN62;
  input [2:0] IN63;
  input [1:0] IN64;
  input [0:0] IN65;
  output [65:0] Out1;
  output [58:0] Out2;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1117;
  wire w1119;
  wire w1121;
  wire w1123;
  wire w1125;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w421);
  FullAdder U1 (w421, IN2[0], IN2[1], w422, w423);
  FullAdder U2 (w423, IN3[0], IN3[1], w424, w425);
  FullAdder U3 (w425, IN4[0], IN4[1], w426, w427);
  FullAdder U4 (w427, IN5[0], IN5[1], w428, w429);
  FullAdder U5 (w429, IN6[0], IN6[1], w430, w431);
  HalfAdder U6 (w422, IN2[2], Out1[2], w433);
  FullAdder U7 (w433, w424, IN3[2], w434, w435);
  FullAdder U8 (w435, w426, IN4[2], w436, w437);
  FullAdder U9 (w437, w428, IN5[2], w438, w439);
  FullAdder U10 (w439, w430, IN6[2], w440, w441);
  FullAdder U11 (w441, w431, IN7[0], w442, w443);
  HalfAdder U12 (w434, IN3[3], Out1[3], w445);
  FullAdder U13 (w445, w436, IN4[3], w446, w447);
  FullAdder U14 (w447, w438, IN5[3], w448, w449);
  FullAdder U15 (w449, w440, IN6[3], w450, w451);
  FullAdder U16 (w451, w442, IN7[1], w452, w453);
  FullAdder U17 (w453, w443, IN8[0], w454, w455);
  HalfAdder U18 (w446, IN4[4], Out1[4], w457);
  FullAdder U19 (w457, w448, IN5[4], w458, w459);
  FullAdder U20 (w459, w450, IN6[4], w460, w461);
  FullAdder U21 (w461, w452, IN7[2], w462, w463);
  FullAdder U22 (w463, w454, IN8[1], w464, w465);
  FullAdder U23 (w465, w455, IN9[0], w466, w467);
  HalfAdder U24 (w458, IN5[5], Out1[5], w469);
  FullAdder U25 (w469, w460, IN6[5], w470, w471);
  FullAdder U26 (w471, w462, IN7[3], w472, w473);
  FullAdder U27 (w473, w464, IN8[2], w474, w475);
  FullAdder U28 (w475, w466, IN9[1], w476, w477);
  FullAdder U29 (w477, w467, IN10[0], w478, w479);
  HalfAdder U30 (w470, IN6[6], Out1[6], w481);
  FullAdder U31 (w481, w472, IN7[4], w482, w483);
  FullAdder U32 (w483, w474, IN8[3], w484, w485);
  FullAdder U33 (w485, w476, IN9[2], w486, w487);
  FullAdder U34 (w487, w478, IN10[1], w488, w489);
  FullAdder U35 (w489, w479, IN11[0], w490, w491);
  HalfAdder U36 (w482, IN7[5], Out1[7], w493);
  FullAdder U37 (w493, w484, IN8[4], w494, w495);
  FullAdder U38 (w495, w486, IN9[3], w496, w497);
  FullAdder U39 (w497, w488, IN10[2], w498, w499);
  FullAdder U40 (w499, w490, IN11[1], w500, w501);
  FullAdder U41 (w501, w491, IN12[0], w502, w503);
  HalfAdder U42 (w494, IN8[5], Out1[8], w505);
  FullAdder U43 (w505, w496, IN9[4], w506, w507);
  FullAdder U44 (w507, w498, IN10[3], w508, w509);
  FullAdder U45 (w509, w500, IN11[2], w510, w511);
  FullAdder U46 (w511, w502, IN12[1], w512, w513);
  FullAdder U47 (w513, w503, IN13[0], w514, w515);
  HalfAdder U48 (w506, IN9[5], Out1[9], w517);
  FullAdder U49 (w517, w508, IN10[4], w518, w519);
  FullAdder U50 (w519, w510, IN11[3], w520, w521);
  FullAdder U51 (w521, w512, IN12[2], w522, w523);
  FullAdder U52 (w523, w514, IN13[1], w524, w525);
  FullAdder U53 (w525, w515, IN14[0], w526, w527);
  HalfAdder U54 (w518, IN10[5], Out1[10], w529);
  FullAdder U55 (w529, w520, IN11[4], w530, w531);
  FullAdder U56 (w531, w522, IN12[3], w532, w533);
  FullAdder U57 (w533, w524, IN13[2], w534, w535);
  FullAdder U58 (w535, w526, IN14[1], w536, w537);
  FullAdder U59 (w537, w527, IN15[0], w538, w539);
  HalfAdder U60 (w530, IN11[5], Out1[11], w541);
  FullAdder U61 (w541, w532, IN12[4], w542, w543);
  FullAdder U62 (w543, w534, IN13[3], w544, w545);
  FullAdder U63 (w545, w536, IN14[2], w546, w547);
  FullAdder U64 (w547, w538, IN15[1], w548, w549);
  FullAdder U65 (w549, w539, IN16[0], w550, w551);
  HalfAdder U66 (w542, IN12[5], Out1[12], w553);
  FullAdder U67 (w553, w544, IN13[4], w554, w555);
  FullAdder U68 (w555, w546, IN14[3], w556, w557);
  FullAdder U69 (w557, w548, IN15[2], w558, w559);
  FullAdder U70 (w559, w550, IN16[1], w560, w561);
  FullAdder U71 (w561, w551, IN17[0], w562, w563);
  HalfAdder U72 (w554, IN13[5], Out1[13], w565);
  FullAdder U73 (w565, w556, IN14[4], w566, w567);
  FullAdder U74 (w567, w558, IN15[3], w568, w569);
  FullAdder U75 (w569, w560, IN16[2], w570, w571);
  FullAdder U76 (w571, w562, IN17[1], w572, w573);
  FullAdder U77 (w573, w563, IN18[0], w574, w575);
  HalfAdder U78 (w566, IN14[5], Out1[14], w577);
  FullAdder U79 (w577, w568, IN15[4], w578, w579);
  FullAdder U80 (w579, w570, IN16[3], w580, w581);
  FullAdder U81 (w581, w572, IN17[2], w582, w583);
  FullAdder U82 (w583, w574, IN18[1], w584, w585);
  FullAdder U83 (w585, w575, IN19[0], w586, w587);
  HalfAdder U84 (w578, IN15[5], Out1[15], w589);
  FullAdder U85 (w589, w580, IN16[4], w590, w591);
  FullAdder U86 (w591, w582, IN17[3], w592, w593);
  FullAdder U87 (w593, w584, IN18[2], w594, w595);
  FullAdder U88 (w595, w586, IN19[1], w596, w597);
  FullAdder U89 (w597, w587, IN20[0], w598, w599);
  HalfAdder U90 (w590, IN16[5], Out1[16], w601);
  FullAdder U91 (w601, w592, IN17[4], w602, w603);
  FullAdder U92 (w603, w594, IN18[3], w604, w605);
  FullAdder U93 (w605, w596, IN19[2], w606, w607);
  FullAdder U94 (w607, w598, IN20[1], w608, w609);
  FullAdder U95 (w609, w599, IN21[0], w610, w611);
  HalfAdder U96 (w602, IN17[5], Out1[17], w613);
  FullAdder U97 (w613, w604, IN18[4], w614, w615);
  FullAdder U98 (w615, w606, IN19[3], w616, w617);
  FullAdder U99 (w617, w608, IN20[2], w618, w619);
  FullAdder U100 (w619, w610, IN21[1], w620, w621);
  FullAdder U101 (w621, w611, IN22[0], w622, w623);
  HalfAdder U102 (w614, IN18[5], Out1[18], w625);
  FullAdder U103 (w625, w616, IN19[4], w626, w627);
  FullAdder U104 (w627, w618, IN20[3], w628, w629);
  FullAdder U105 (w629, w620, IN21[2], w630, w631);
  FullAdder U106 (w631, w622, IN22[1], w632, w633);
  FullAdder U107 (w633, w623, IN23[0], w634, w635);
  HalfAdder U108 (w626, IN19[5], Out1[19], w637);
  FullAdder U109 (w637, w628, IN20[4], w638, w639);
  FullAdder U110 (w639, w630, IN21[3], w640, w641);
  FullAdder U111 (w641, w632, IN22[2], w642, w643);
  FullAdder U112 (w643, w634, IN23[1], w644, w645);
  FullAdder U113 (w645, w635, IN24[0], w646, w647);
  HalfAdder U114 (w638, IN20[5], Out1[20], w649);
  FullAdder U115 (w649, w640, IN21[4], w650, w651);
  FullAdder U116 (w651, w642, IN22[3], w652, w653);
  FullAdder U117 (w653, w644, IN23[2], w654, w655);
  FullAdder U118 (w655, w646, IN24[1], w656, w657);
  FullAdder U119 (w657, w647, IN25[0], w658, w659);
  HalfAdder U120 (w650, IN21[5], Out1[21], w661);
  FullAdder U121 (w661, w652, IN22[4], w662, w663);
  FullAdder U122 (w663, w654, IN23[3], w664, w665);
  FullAdder U123 (w665, w656, IN24[2], w666, w667);
  FullAdder U124 (w667, w658, IN25[1], w668, w669);
  FullAdder U125 (w669, w659, IN26[0], w670, w671);
  HalfAdder U126 (w662, IN22[5], Out1[22], w673);
  FullAdder U127 (w673, w664, IN23[4], w674, w675);
  FullAdder U128 (w675, w666, IN24[3], w676, w677);
  FullAdder U129 (w677, w668, IN25[2], w678, w679);
  FullAdder U130 (w679, w670, IN26[1], w680, w681);
  FullAdder U131 (w681, w671, IN27[0], w682, w683);
  HalfAdder U132 (w674, IN23[5], Out1[23], w685);
  FullAdder U133 (w685, w676, IN24[4], w686, w687);
  FullAdder U134 (w687, w678, IN25[3], w688, w689);
  FullAdder U135 (w689, w680, IN26[2], w690, w691);
  FullAdder U136 (w691, w682, IN27[1], w692, w693);
  FullAdder U137 (w693, w683, IN28[0], w694, w695);
  HalfAdder U138 (w686, IN24[5], Out1[24], w697);
  FullAdder U139 (w697, w688, IN25[4], w698, w699);
  FullAdder U140 (w699, w690, IN26[3], w700, w701);
  FullAdder U141 (w701, w692, IN27[2], w702, w703);
  FullAdder U142 (w703, w694, IN28[1], w704, w705);
  FullAdder U143 (w705, w695, IN29[0], w706, w707);
  HalfAdder U144 (w698, IN25[5], Out1[25], w709);
  FullAdder U145 (w709, w700, IN26[4], w710, w711);
  FullAdder U146 (w711, w702, IN27[3], w712, w713);
  FullAdder U147 (w713, w704, IN28[2], w714, w715);
  FullAdder U148 (w715, w706, IN29[1], w716, w717);
  FullAdder U149 (w717, w707, IN30[0], w718, w719);
  HalfAdder U150 (w710, IN26[5], Out1[26], w721);
  FullAdder U151 (w721, w712, IN27[4], w722, w723);
  FullAdder U152 (w723, w714, IN28[3], w724, w725);
  FullAdder U153 (w725, w716, IN29[2], w726, w727);
  FullAdder U154 (w727, w718, IN30[1], w728, w729);
  FullAdder U155 (w729, w719, IN31[0], w730, w731);
  HalfAdder U156 (w722, IN27[5], Out1[27], w733);
  FullAdder U157 (w733, w724, IN28[4], w734, w735);
  FullAdder U158 (w735, w726, IN29[3], w736, w737);
  FullAdder U159 (w737, w728, IN30[2], w738, w739);
  FullAdder U160 (w739, w730, IN31[1], w740, w741);
  FullAdder U161 (w741, w731, IN32[0], w742, w743);
  HalfAdder U162 (w734, IN28[5], Out1[28], w745);
  FullAdder U163 (w745, w736, IN29[4], w746, w747);
  FullAdder U164 (w747, w738, IN30[3], w748, w749);
  FullAdder U165 (w749, w740, IN31[2], w750, w751);
  FullAdder U166 (w751, w742, IN32[1], w752, w753);
  FullAdder U167 (w753, w743, IN33[0], w754, w755);
  HalfAdder U168 (w746, IN29[5], Out1[29], w757);
  FullAdder U169 (w757, w748, IN30[4], w758, w759);
  FullAdder U170 (w759, w750, IN31[3], w760, w761);
  FullAdder U171 (w761, w752, IN32[2], w762, w763);
  FullAdder U172 (w763, w754, IN33[1], w764, w765);
  FullAdder U173 (w765, w755, IN34[0], w766, w767);
  HalfAdder U174 (w758, IN30[5], Out1[30], w769);
  FullAdder U175 (w769, w760, IN31[4], w770, w771);
  FullAdder U176 (w771, w762, IN32[3], w772, w773);
  FullAdder U177 (w773, w764, IN33[2], w774, w775);
  FullAdder U178 (w775, w766, IN34[1], w776, w777);
  FullAdder U179 (w777, w767, IN35[0], w778, w779);
  HalfAdder U180 (w770, IN31[5], Out1[31], w781);
  FullAdder U181 (w781, w772, IN32[4], w782, w783);
  FullAdder U182 (w783, w774, IN33[3], w784, w785);
  FullAdder U183 (w785, w776, IN34[2], w786, w787);
  FullAdder U184 (w787, w778, IN35[1], w788, w789);
  FullAdder U185 (w789, w779, IN36[0], w790, w791);
  HalfAdder U186 (w782, IN32[5], Out1[32], w793);
  FullAdder U187 (w793, w784, IN33[4], w794, w795);
  FullAdder U188 (w795, w786, IN34[3], w796, w797);
  FullAdder U189 (w797, w788, IN35[2], w798, w799);
  FullAdder U190 (w799, w790, IN36[1], w800, w801);
  FullAdder U191 (w801, w791, IN37[0], w802, w803);
  HalfAdder U192 (w794, IN33[5], Out1[33], w805);
  FullAdder U193 (w805, w796, IN34[4], w806, w807);
  FullAdder U194 (w807, w798, IN35[3], w808, w809);
  FullAdder U195 (w809, w800, IN36[2], w810, w811);
  FullAdder U196 (w811, w802, IN37[1], w812, w813);
  FullAdder U197 (w813, w803, IN38[0], w814, w815);
  HalfAdder U198 (w806, IN34[5], Out1[34], w817);
  FullAdder U199 (w817, w808, IN35[4], w818, w819);
  FullAdder U200 (w819, w810, IN36[3], w820, w821);
  FullAdder U201 (w821, w812, IN37[2], w822, w823);
  FullAdder U202 (w823, w814, IN38[1], w824, w825);
  FullAdder U203 (w825, w815, IN39[0], w826, w827);
  HalfAdder U204 (w818, IN35[5], Out1[35], w829);
  FullAdder U205 (w829, w820, IN36[4], w830, w831);
  FullAdder U206 (w831, w822, IN37[3], w832, w833);
  FullAdder U207 (w833, w824, IN38[2], w834, w835);
  FullAdder U208 (w835, w826, IN39[1], w836, w837);
  FullAdder U209 (w837, w827, IN40[0], w838, w839);
  HalfAdder U210 (w830, IN36[5], Out1[36], w841);
  FullAdder U211 (w841, w832, IN37[4], w842, w843);
  FullAdder U212 (w843, w834, IN38[3], w844, w845);
  FullAdder U213 (w845, w836, IN39[2], w846, w847);
  FullAdder U214 (w847, w838, IN40[1], w848, w849);
  FullAdder U215 (w849, w839, IN41[0], w850, w851);
  HalfAdder U216 (w842, IN37[5], Out1[37], w853);
  FullAdder U217 (w853, w844, IN38[4], w854, w855);
  FullAdder U218 (w855, w846, IN39[3], w856, w857);
  FullAdder U219 (w857, w848, IN40[2], w858, w859);
  FullAdder U220 (w859, w850, IN41[1], w860, w861);
  FullAdder U221 (w861, w851, IN42[0], w862, w863);
  HalfAdder U222 (w854, IN38[5], Out1[38], w865);
  FullAdder U223 (w865, w856, IN39[4], w866, w867);
  FullAdder U224 (w867, w858, IN40[3], w868, w869);
  FullAdder U225 (w869, w860, IN41[2], w870, w871);
  FullAdder U226 (w871, w862, IN42[1], w872, w873);
  FullAdder U227 (w873, w863, IN43[0], w874, w875);
  HalfAdder U228 (w866, IN39[5], Out1[39], w877);
  FullAdder U229 (w877, w868, IN40[4], w878, w879);
  FullAdder U230 (w879, w870, IN41[3], w880, w881);
  FullAdder U231 (w881, w872, IN42[2], w882, w883);
  FullAdder U232 (w883, w874, IN43[1], w884, w885);
  FullAdder U233 (w885, w875, IN44[0], w886, w887);
  HalfAdder U234 (w878, IN40[5], Out1[40], w889);
  FullAdder U235 (w889, w880, IN41[4], w890, w891);
  FullAdder U236 (w891, w882, IN42[3], w892, w893);
  FullAdder U237 (w893, w884, IN43[2], w894, w895);
  FullAdder U238 (w895, w886, IN44[1], w896, w897);
  FullAdder U239 (w897, w887, IN45[0], w898, w899);
  HalfAdder U240 (w890, IN41[5], Out1[41], w901);
  FullAdder U241 (w901, w892, IN42[4], w902, w903);
  FullAdder U242 (w903, w894, IN43[3], w904, w905);
  FullAdder U243 (w905, w896, IN44[2], w906, w907);
  FullAdder U244 (w907, w898, IN45[1], w908, w909);
  FullAdder U245 (w909, w899, IN46[0], w910, w911);
  HalfAdder U246 (w902, IN42[5], Out1[42], w913);
  FullAdder U247 (w913, w904, IN43[4], w914, w915);
  FullAdder U248 (w915, w906, IN44[3], w916, w917);
  FullAdder U249 (w917, w908, IN45[2], w918, w919);
  FullAdder U250 (w919, w910, IN46[1], w920, w921);
  FullAdder U251 (w921, w911, IN47[0], w922, w923);
  HalfAdder U252 (w914, IN43[5], Out1[43], w925);
  FullAdder U253 (w925, w916, IN44[4], w926, w927);
  FullAdder U254 (w927, w918, IN45[3], w928, w929);
  FullAdder U255 (w929, w920, IN46[2], w930, w931);
  FullAdder U256 (w931, w922, IN47[1], w932, w933);
  FullAdder U257 (w933, w923, IN48[0], w934, w935);
  HalfAdder U258 (w926, IN44[5], Out1[44], w937);
  FullAdder U259 (w937, w928, IN45[4], w938, w939);
  FullAdder U260 (w939, w930, IN46[3], w940, w941);
  FullAdder U261 (w941, w932, IN47[2], w942, w943);
  FullAdder U262 (w943, w934, IN48[1], w944, w945);
  FullAdder U263 (w945, w935, IN49[0], w946, w947);
  HalfAdder U264 (w938, IN45[5], Out1[45], w949);
  FullAdder U265 (w949, w940, IN46[4], w950, w951);
  FullAdder U266 (w951, w942, IN47[3], w952, w953);
  FullAdder U267 (w953, w944, IN48[2], w954, w955);
  FullAdder U268 (w955, w946, IN49[1], w956, w957);
  FullAdder U269 (w957, w947, IN50[0], w958, w959);
  HalfAdder U270 (w950, IN46[5], Out1[46], w961);
  FullAdder U271 (w961, w952, IN47[4], w962, w963);
  FullAdder U272 (w963, w954, IN48[3], w964, w965);
  FullAdder U273 (w965, w956, IN49[2], w966, w967);
  FullAdder U274 (w967, w958, IN50[1], w968, w969);
  FullAdder U275 (w969, w959, IN51[0], w970, w971);
  HalfAdder U276 (w962, IN47[5], Out1[47], w973);
  FullAdder U277 (w973, w964, IN48[4], w974, w975);
  FullAdder U278 (w975, w966, IN49[3], w976, w977);
  FullAdder U279 (w977, w968, IN50[2], w978, w979);
  FullAdder U280 (w979, w970, IN51[1], w980, w981);
  FullAdder U281 (w981, w971, IN52[0], w982, w983);
  HalfAdder U282 (w974, IN48[5], Out1[48], w985);
  FullAdder U283 (w985, w976, IN49[4], w986, w987);
  FullAdder U284 (w987, w978, IN50[3], w988, w989);
  FullAdder U285 (w989, w980, IN51[2], w990, w991);
  FullAdder U286 (w991, w982, IN52[1], w992, w993);
  FullAdder U287 (w993, w983, IN53[0], w994, w995);
  HalfAdder U288 (w986, IN49[5], Out1[49], w997);
  FullAdder U289 (w997, w988, IN50[4], w998, w999);
  FullAdder U290 (w999, w990, IN51[3], w1000, w1001);
  FullAdder U291 (w1001, w992, IN52[2], w1002, w1003);
  FullAdder U292 (w1003, w994, IN53[1], w1004, w1005);
  FullAdder U293 (w1005, w995, IN54[0], w1006, w1007);
  HalfAdder U294 (w998, IN50[5], Out1[50], w1009);
  FullAdder U295 (w1009, w1000, IN51[4], w1010, w1011);
  FullAdder U296 (w1011, w1002, IN52[3], w1012, w1013);
  FullAdder U297 (w1013, w1004, IN53[2], w1014, w1015);
  FullAdder U298 (w1015, w1006, IN54[1], w1016, w1017);
  FullAdder U299 (w1017, w1007, IN55[0], w1018, w1019);
  HalfAdder U300 (w1010, IN51[5], Out1[51], w1021);
  FullAdder U301 (w1021, w1012, IN52[4], w1022, w1023);
  FullAdder U302 (w1023, w1014, IN53[3], w1024, w1025);
  FullAdder U303 (w1025, w1016, IN54[2], w1026, w1027);
  FullAdder U304 (w1027, w1018, IN55[1], w1028, w1029);
  FullAdder U305 (w1029, w1019, IN56[0], w1030, w1031);
  HalfAdder U306 (w1022, IN52[5], Out1[52], w1033);
  FullAdder U307 (w1033, w1024, IN53[4], w1034, w1035);
  FullAdder U308 (w1035, w1026, IN54[3], w1036, w1037);
  FullAdder U309 (w1037, w1028, IN55[2], w1038, w1039);
  FullAdder U310 (w1039, w1030, IN56[1], w1040, w1041);
  FullAdder U311 (w1041, w1031, IN57[0], w1042, w1043);
  HalfAdder U312 (w1034, IN53[5], Out1[53], w1045);
  FullAdder U313 (w1045, w1036, IN54[4], w1046, w1047);
  FullAdder U314 (w1047, w1038, IN55[3], w1048, w1049);
  FullAdder U315 (w1049, w1040, IN56[2], w1050, w1051);
  FullAdder U316 (w1051, w1042, IN57[1], w1052, w1053);
  FullAdder U317 (w1053, w1043, IN58[0], w1054, w1055);
  HalfAdder U318 (w1046, IN54[5], Out1[54], w1057);
  FullAdder U319 (w1057, w1048, IN55[4], w1058, w1059);
  FullAdder U320 (w1059, w1050, IN56[3], w1060, w1061);
  FullAdder U321 (w1061, w1052, IN57[2], w1062, w1063);
  FullAdder U322 (w1063, w1054, IN58[1], w1064, w1065);
  FullAdder U323 (w1065, w1055, IN59[0], w1066, w1067);
  HalfAdder U324 (w1058, IN55[5], Out1[55], w1069);
  FullAdder U325 (w1069, w1060, IN56[4], w1070, w1071);
  FullAdder U326 (w1071, w1062, IN57[3], w1072, w1073);
  FullAdder U327 (w1073, w1064, IN58[2], w1074, w1075);
  FullAdder U328 (w1075, w1066, IN59[1], w1076, w1077);
  FullAdder U329 (w1077, w1067, IN60[0], w1078, w1079);
  HalfAdder U330 (w1070, IN56[5], Out1[56], w1081);
  FullAdder U331 (w1081, w1072, IN57[4], w1082, w1083);
  FullAdder U332 (w1083, w1074, IN58[3], w1084, w1085);
  FullAdder U333 (w1085, w1076, IN59[2], w1086, w1087);
  FullAdder U334 (w1087, w1078, IN60[1], w1088, w1089);
  FullAdder U335 (w1089, w1079, IN61[0], w1090, w1091);
  HalfAdder U336 (w1082, IN57[5], Out1[57], w1093);
  FullAdder U337 (w1093, w1084, IN58[4], w1094, w1095);
  FullAdder U338 (w1095, w1086, IN59[3], w1096, w1097);
  FullAdder U339 (w1097, w1088, IN60[2], w1098, w1099);
  FullAdder U340 (w1099, w1090, IN61[1], w1100, w1101);
  FullAdder U341 (w1101, w1091, IN62[0], w1102, w1103);
  HalfAdder U342 (w1094, IN58[5], Out1[58], w1105);
  FullAdder U343 (w1105, w1096, IN59[4], w1106, w1107);
  FullAdder U344 (w1107, w1098, IN60[3], w1108, w1109);
  FullAdder U345 (w1109, w1100, IN61[2], w1110, w1111);
  FullAdder U346 (w1111, w1102, IN62[1], w1112, w1113);
  FullAdder U347 (w1113, w1103, IN63[0], w1114, w1115);
  HalfAdder U348 (w1106, IN59[5], Out1[59], w1117);
  FullAdder U349 (w1117, w1108, IN60[4], Out1[60], w1119);
  FullAdder U350 (w1119, w1110, IN61[3], Out1[61], w1121);
  FullAdder U351 (w1121, w1112, IN62[2], Out1[62], w1123);
  FullAdder U352 (w1123, w1114, IN63[1], Out1[63], w1125);
  FullAdder U353 (w1125, w1115, IN64[0], Out1[64], Out1[65]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN7[6];
  assign Out2[1] = IN8[6];
  assign Out2[2] = IN9[6];
  assign Out2[3] = IN10[6];
  assign Out2[4] = IN11[6];
  assign Out2[5] = IN12[6];
  assign Out2[6] = IN13[6];
  assign Out2[7] = IN14[6];
  assign Out2[8] = IN15[6];
  assign Out2[9] = IN16[6];
  assign Out2[10] = IN17[6];
  assign Out2[11] = IN18[6];
  assign Out2[12] = IN19[6];
  assign Out2[13] = IN20[6];
  assign Out2[14] = IN21[6];
  assign Out2[15] = IN22[6];
  assign Out2[16] = IN23[6];
  assign Out2[17] = IN24[6];
  assign Out2[18] = IN25[6];
  assign Out2[19] = IN26[6];
  assign Out2[20] = IN27[6];
  assign Out2[21] = IN28[6];
  assign Out2[22] = IN29[6];
  assign Out2[23] = IN30[6];
  assign Out2[24] = IN31[6];
  assign Out2[25] = IN32[6];
  assign Out2[26] = IN33[6];
  assign Out2[27] = IN34[6];
  assign Out2[28] = IN35[6];
  assign Out2[29] = IN36[6];
  assign Out2[30] = IN37[6];
  assign Out2[31] = IN38[6];
  assign Out2[32] = IN39[6];
  assign Out2[33] = IN40[6];
  assign Out2[34] = IN41[6];
  assign Out2[35] = IN42[6];
  assign Out2[36] = IN43[6];
  assign Out2[37] = IN44[6];
  assign Out2[38] = IN45[6];
  assign Out2[39] = IN46[6];
  assign Out2[40] = IN47[6];
  assign Out2[41] = IN48[6];
  assign Out2[42] = IN49[6];
  assign Out2[43] = IN50[6];
  assign Out2[44] = IN51[6];
  assign Out2[45] = IN52[6];
  assign Out2[46] = IN53[6];
  assign Out2[47] = IN54[6];
  assign Out2[48] = IN55[6];
  assign Out2[49] = IN56[6];
  assign Out2[50] = IN57[6];
  assign Out2[51] = IN58[6];
  assign Out2[52] = IN59[6];
  assign Out2[53] = IN60[5];
  assign Out2[54] = IN61[4];
  assign Out2[55] = IN62[3];
  assign Out2[56] = IN63[2];
  assign Out2[57] = IN64[1];
  assign Out2[58] = IN65[0];

endmodule
module RC_59_59(IN1, IN2, Out);
  input [58:0] IN1;
  input [58:0] IN2;
  output [59:0] Out;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  wire w231;
  wire w233;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w119);
  FullAdder U1 (IN1[1], IN2[1], w119, Out[1], w121);
  FullAdder U2 (IN1[2], IN2[2], w121, Out[2], w123);
  FullAdder U3 (IN1[3], IN2[3], w123, Out[3], w125);
  FullAdder U4 (IN1[4], IN2[4], w125, Out[4], w127);
  FullAdder U5 (IN1[5], IN2[5], w127, Out[5], w129);
  FullAdder U6 (IN1[6], IN2[6], w129, Out[6], w131);
  FullAdder U7 (IN1[7], IN2[7], w131, Out[7], w133);
  FullAdder U8 (IN1[8], IN2[8], w133, Out[8], w135);
  FullAdder U9 (IN1[9], IN2[9], w135, Out[9], w137);
  FullAdder U10 (IN1[10], IN2[10], w137, Out[10], w139);
  FullAdder U11 (IN1[11], IN2[11], w139, Out[11], w141);
  FullAdder U12 (IN1[12], IN2[12], w141, Out[12], w143);
  FullAdder U13 (IN1[13], IN2[13], w143, Out[13], w145);
  FullAdder U14 (IN1[14], IN2[14], w145, Out[14], w147);
  FullAdder U15 (IN1[15], IN2[15], w147, Out[15], w149);
  FullAdder U16 (IN1[16], IN2[16], w149, Out[16], w151);
  FullAdder U17 (IN1[17], IN2[17], w151, Out[17], w153);
  FullAdder U18 (IN1[18], IN2[18], w153, Out[18], w155);
  FullAdder U19 (IN1[19], IN2[19], w155, Out[19], w157);
  FullAdder U20 (IN1[20], IN2[20], w157, Out[20], w159);
  FullAdder U21 (IN1[21], IN2[21], w159, Out[21], w161);
  FullAdder U22 (IN1[22], IN2[22], w161, Out[22], w163);
  FullAdder U23 (IN1[23], IN2[23], w163, Out[23], w165);
  FullAdder U24 (IN1[24], IN2[24], w165, Out[24], w167);
  FullAdder U25 (IN1[25], IN2[25], w167, Out[25], w169);
  FullAdder U26 (IN1[26], IN2[26], w169, Out[26], w171);
  FullAdder U27 (IN1[27], IN2[27], w171, Out[27], w173);
  FullAdder U28 (IN1[28], IN2[28], w173, Out[28], w175);
  FullAdder U29 (IN1[29], IN2[29], w175, Out[29], w177);
  FullAdder U30 (IN1[30], IN2[30], w177, Out[30], w179);
  FullAdder U31 (IN1[31], IN2[31], w179, Out[31], w181);
  FullAdder U32 (IN1[32], IN2[32], w181, Out[32], w183);
  FullAdder U33 (IN1[33], IN2[33], w183, Out[33], w185);
  FullAdder U34 (IN1[34], IN2[34], w185, Out[34], w187);
  FullAdder U35 (IN1[35], IN2[35], w187, Out[35], w189);
  FullAdder U36 (IN1[36], IN2[36], w189, Out[36], w191);
  FullAdder U37 (IN1[37], IN2[37], w191, Out[37], w193);
  FullAdder U38 (IN1[38], IN2[38], w193, Out[38], w195);
  FullAdder U39 (IN1[39], IN2[39], w195, Out[39], w197);
  FullAdder U40 (IN1[40], IN2[40], w197, Out[40], w199);
  FullAdder U41 (IN1[41], IN2[41], w199, Out[41], w201);
  FullAdder U42 (IN1[42], IN2[42], w201, Out[42], w203);
  FullAdder U43 (IN1[43], IN2[43], w203, Out[43], w205);
  FullAdder U44 (IN1[44], IN2[44], w205, Out[44], w207);
  FullAdder U45 (IN1[45], IN2[45], w207, Out[45], w209);
  FullAdder U46 (IN1[46], IN2[46], w209, Out[46], w211);
  FullAdder U47 (IN1[47], IN2[47], w211, Out[47], w213);
  FullAdder U48 (IN1[48], IN2[48], w213, Out[48], w215);
  FullAdder U49 (IN1[49], IN2[49], w215, Out[49], w217);
  FullAdder U50 (IN1[50], IN2[50], w217, Out[50], w219);
  FullAdder U51 (IN1[51], IN2[51], w219, Out[51], w221);
  FullAdder U52 (IN1[52], IN2[52], w221, Out[52], w223);
  FullAdder U53 (IN1[53], IN2[53], w223, Out[53], w225);
  FullAdder U54 (IN1[54], IN2[54], w225, Out[54], w227);
  FullAdder U55 (IN1[55], IN2[55], w227, Out[55], w229);
  FullAdder U56 (IN1[56], IN2[56], w229, Out[56], w231);
  FullAdder U57 (IN1[57], IN2[57], w231, Out[57], w233);
  FullAdder U58 (IN1[58], IN2[58], w233, Out[58], Out[59]);

endmodule
module NR_7_60(IN1, IN2, Out);
  input [6:0] IN1;
  input [59:0] IN2;
  output [66:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [6:0] P37;
  wire [6:0] P38;
  wire [6:0] P39;
  wire [6:0] P40;
  wire [6:0] P41;
  wire [6:0] P42;
  wire [6:0] P43;
  wire [6:0] P44;
  wire [6:0] P45;
  wire [6:0] P46;
  wire [6:0] P47;
  wire [6:0] P48;
  wire [6:0] P49;
  wire [6:0] P50;
  wire [6:0] P51;
  wire [6:0] P52;
  wire [6:0] P53;
  wire [6:0] P54;
  wire [6:0] P55;
  wire [6:0] P56;
  wire [6:0] P57;
  wire [6:0] P58;
  wire [6:0] P59;
  wire [5:0] P60;
  wire [4:0] P61;
  wire [3:0] P62;
  wire [2:0] P63;
  wire [1:0] P64;
  wire [0:0] P65;
  wire [65:0] R1;
  wire [58:0] R2;
  wire [66:0] aOut;
  U_SP_7_60 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, R1, R2);
  RC_59_59 S2 (R1[65:7], R2, aOut[66:7]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign Out = aOut[66:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
