//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 7
  second input length: 59
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_7_59(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64);
  input [6:0] IN1;
  input [58:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [6:0] P37;
  output [6:0] P38;
  output [6:0] P39;
  output [6:0] P40;
  output [6:0] P41;
  output [6:0] P42;
  output [6:0] P43;
  output [6:0] P44;
  output [6:0] P45;
  output [6:0] P46;
  output [6:0] P47;
  output [6:0] P48;
  output [6:0] P49;
  output [6:0] P50;
  output [6:0] P51;
  output [6:0] P52;
  output [6:0] P53;
  output [6:0] P54;
  output [6:0] P55;
  output [6:0] P56;
  output [6:0] P57;
  output [6:0] P58;
  output [5:0] P59;
  output [4:0] P60;
  output [3:0] P61;
  output [2:0] P62;
  output [1:0] P63;
  output [0:0] P64;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[0] = IN1[1]&IN2[58];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[1] = IN1[2]&IN2[57];
  assign P60[0] = IN1[2]&IN2[58];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[2] = IN1[3]&IN2[56];
  assign P60[1] = IN1[3]&IN2[57];
  assign P61[0] = IN1[3]&IN2[58];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[3] = IN1[4]&IN2[55];
  assign P60[2] = IN1[4]&IN2[56];
  assign P61[1] = IN1[4]&IN2[57];
  assign P62[0] = IN1[4]&IN2[58];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[4] = IN1[5]&IN2[54];
  assign P60[3] = IN1[5]&IN2[55];
  assign P61[2] = IN1[5]&IN2[56];
  assign P62[1] = IN1[5]&IN2[57];
  assign P63[0] = IN1[5]&IN2[58];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[5] = IN1[6]&IN2[53];
  assign P60[4] = IN1[6]&IN2[54];
  assign P61[3] = IN1[6]&IN2[55];
  assign P62[2] = IN1[6]&IN2[56];
  assign P63[1] = IN1[6]&IN2[57];
  assign P64[0] = IN1[6]&IN2[58];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [6:0] IN37;
  input [6:0] IN38;
  input [6:0] IN39;
  input [6:0] IN40;
  input [6:0] IN41;
  input [6:0] IN42;
  input [6:0] IN43;
  input [6:0] IN44;
  input [6:0] IN45;
  input [6:0] IN46;
  input [6:0] IN47;
  input [6:0] IN48;
  input [6:0] IN49;
  input [6:0] IN50;
  input [6:0] IN51;
  input [6:0] IN52;
  input [6:0] IN53;
  input [6:0] IN54;
  input [6:0] IN55;
  input [6:0] IN56;
  input [6:0] IN57;
  input [6:0] IN58;
  input [5:0] IN59;
  input [4:0] IN60;
  input [3:0] IN61;
  input [2:0] IN62;
  input [1:0] IN63;
  input [0:0] IN64;
  output [64:0] Out1;
  output [57:0] Out2;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1098;
  wire w1100;
  wire w1102;
  wire w1104;
  wire w1106;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w414);
  FullAdder U1 (w414, IN2[0], IN2[1], w415, w416);
  FullAdder U2 (w416, IN3[0], IN3[1], w417, w418);
  FullAdder U3 (w418, IN4[0], IN4[1], w419, w420);
  FullAdder U4 (w420, IN5[0], IN5[1], w421, w422);
  FullAdder U5 (w422, IN6[0], IN6[1], w423, w424);
  HalfAdder U6 (w415, IN2[2], Out1[2], w426);
  FullAdder U7 (w426, w417, IN3[2], w427, w428);
  FullAdder U8 (w428, w419, IN4[2], w429, w430);
  FullAdder U9 (w430, w421, IN5[2], w431, w432);
  FullAdder U10 (w432, w423, IN6[2], w433, w434);
  FullAdder U11 (w434, w424, IN7[0], w435, w436);
  HalfAdder U12 (w427, IN3[3], Out1[3], w438);
  FullAdder U13 (w438, w429, IN4[3], w439, w440);
  FullAdder U14 (w440, w431, IN5[3], w441, w442);
  FullAdder U15 (w442, w433, IN6[3], w443, w444);
  FullAdder U16 (w444, w435, IN7[1], w445, w446);
  FullAdder U17 (w446, w436, IN8[0], w447, w448);
  HalfAdder U18 (w439, IN4[4], Out1[4], w450);
  FullAdder U19 (w450, w441, IN5[4], w451, w452);
  FullAdder U20 (w452, w443, IN6[4], w453, w454);
  FullAdder U21 (w454, w445, IN7[2], w455, w456);
  FullAdder U22 (w456, w447, IN8[1], w457, w458);
  FullAdder U23 (w458, w448, IN9[0], w459, w460);
  HalfAdder U24 (w451, IN5[5], Out1[5], w462);
  FullAdder U25 (w462, w453, IN6[5], w463, w464);
  FullAdder U26 (w464, w455, IN7[3], w465, w466);
  FullAdder U27 (w466, w457, IN8[2], w467, w468);
  FullAdder U28 (w468, w459, IN9[1], w469, w470);
  FullAdder U29 (w470, w460, IN10[0], w471, w472);
  HalfAdder U30 (w463, IN6[6], Out1[6], w474);
  FullAdder U31 (w474, w465, IN7[4], w475, w476);
  FullAdder U32 (w476, w467, IN8[3], w477, w478);
  FullAdder U33 (w478, w469, IN9[2], w479, w480);
  FullAdder U34 (w480, w471, IN10[1], w481, w482);
  FullAdder U35 (w482, w472, IN11[0], w483, w484);
  HalfAdder U36 (w475, IN7[5], Out1[7], w486);
  FullAdder U37 (w486, w477, IN8[4], w487, w488);
  FullAdder U38 (w488, w479, IN9[3], w489, w490);
  FullAdder U39 (w490, w481, IN10[2], w491, w492);
  FullAdder U40 (w492, w483, IN11[1], w493, w494);
  FullAdder U41 (w494, w484, IN12[0], w495, w496);
  HalfAdder U42 (w487, IN8[5], Out1[8], w498);
  FullAdder U43 (w498, w489, IN9[4], w499, w500);
  FullAdder U44 (w500, w491, IN10[3], w501, w502);
  FullAdder U45 (w502, w493, IN11[2], w503, w504);
  FullAdder U46 (w504, w495, IN12[1], w505, w506);
  FullAdder U47 (w506, w496, IN13[0], w507, w508);
  HalfAdder U48 (w499, IN9[5], Out1[9], w510);
  FullAdder U49 (w510, w501, IN10[4], w511, w512);
  FullAdder U50 (w512, w503, IN11[3], w513, w514);
  FullAdder U51 (w514, w505, IN12[2], w515, w516);
  FullAdder U52 (w516, w507, IN13[1], w517, w518);
  FullAdder U53 (w518, w508, IN14[0], w519, w520);
  HalfAdder U54 (w511, IN10[5], Out1[10], w522);
  FullAdder U55 (w522, w513, IN11[4], w523, w524);
  FullAdder U56 (w524, w515, IN12[3], w525, w526);
  FullAdder U57 (w526, w517, IN13[2], w527, w528);
  FullAdder U58 (w528, w519, IN14[1], w529, w530);
  FullAdder U59 (w530, w520, IN15[0], w531, w532);
  HalfAdder U60 (w523, IN11[5], Out1[11], w534);
  FullAdder U61 (w534, w525, IN12[4], w535, w536);
  FullAdder U62 (w536, w527, IN13[3], w537, w538);
  FullAdder U63 (w538, w529, IN14[2], w539, w540);
  FullAdder U64 (w540, w531, IN15[1], w541, w542);
  FullAdder U65 (w542, w532, IN16[0], w543, w544);
  HalfAdder U66 (w535, IN12[5], Out1[12], w546);
  FullAdder U67 (w546, w537, IN13[4], w547, w548);
  FullAdder U68 (w548, w539, IN14[3], w549, w550);
  FullAdder U69 (w550, w541, IN15[2], w551, w552);
  FullAdder U70 (w552, w543, IN16[1], w553, w554);
  FullAdder U71 (w554, w544, IN17[0], w555, w556);
  HalfAdder U72 (w547, IN13[5], Out1[13], w558);
  FullAdder U73 (w558, w549, IN14[4], w559, w560);
  FullAdder U74 (w560, w551, IN15[3], w561, w562);
  FullAdder U75 (w562, w553, IN16[2], w563, w564);
  FullAdder U76 (w564, w555, IN17[1], w565, w566);
  FullAdder U77 (w566, w556, IN18[0], w567, w568);
  HalfAdder U78 (w559, IN14[5], Out1[14], w570);
  FullAdder U79 (w570, w561, IN15[4], w571, w572);
  FullAdder U80 (w572, w563, IN16[3], w573, w574);
  FullAdder U81 (w574, w565, IN17[2], w575, w576);
  FullAdder U82 (w576, w567, IN18[1], w577, w578);
  FullAdder U83 (w578, w568, IN19[0], w579, w580);
  HalfAdder U84 (w571, IN15[5], Out1[15], w582);
  FullAdder U85 (w582, w573, IN16[4], w583, w584);
  FullAdder U86 (w584, w575, IN17[3], w585, w586);
  FullAdder U87 (w586, w577, IN18[2], w587, w588);
  FullAdder U88 (w588, w579, IN19[1], w589, w590);
  FullAdder U89 (w590, w580, IN20[0], w591, w592);
  HalfAdder U90 (w583, IN16[5], Out1[16], w594);
  FullAdder U91 (w594, w585, IN17[4], w595, w596);
  FullAdder U92 (w596, w587, IN18[3], w597, w598);
  FullAdder U93 (w598, w589, IN19[2], w599, w600);
  FullAdder U94 (w600, w591, IN20[1], w601, w602);
  FullAdder U95 (w602, w592, IN21[0], w603, w604);
  HalfAdder U96 (w595, IN17[5], Out1[17], w606);
  FullAdder U97 (w606, w597, IN18[4], w607, w608);
  FullAdder U98 (w608, w599, IN19[3], w609, w610);
  FullAdder U99 (w610, w601, IN20[2], w611, w612);
  FullAdder U100 (w612, w603, IN21[1], w613, w614);
  FullAdder U101 (w614, w604, IN22[0], w615, w616);
  HalfAdder U102 (w607, IN18[5], Out1[18], w618);
  FullAdder U103 (w618, w609, IN19[4], w619, w620);
  FullAdder U104 (w620, w611, IN20[3], w621, w622);
  FullAdder U105 (w622, w613, IN21[2], w623, w624);
  FullAdder U106 (w624, w615, IN22[1], w625, w626);
  FullAdder U107 (w626, w616, IN23[0], w627, w628);
  HalfAdder U108 (w619, IN19[5], Out1[19], w630);
  FullAdder U109 (w630, w621, IN20[4], w631, w632);
  FullAdder U110 (w632, w623, IN21[3], w633, w634);
  FullAdder U111 (w634, w625, IN22[2], w635, w636);
  FullAdder U112 (w636, w627, IN23[1], w637, w638);
  FullAdder U113 (w638, w628, IN24[0], w639, w640);
  HalfAdder U114 (w631, IN20[5], Out1[20], w642);
  FullAdder U115 (w642, w633, IN21[4], w643, w644);
  FullAdder U116 (w644, w635, IN22[3], w645, w646);
  FullAdder U117 (w646, w637, IN23[2], w647, w648);
  FullAdder U118 (w648, w639, IN24[1], w649, w650);
  FullAdder U119 (w650, w640, IN25[0], w651, w652);
  HalfAdder U120 (w643, IN21[5], Out1[21], w654);
  FullAdder U121 (w654, w645, IN22[4], w655, w656);
  FullAdder U122 (w656, w647, IN23[3], w657, w658);
  FullAdder U123 (w658, w649, IN24[2], w659, w660);
  FullAdder U124 (w660, w651, IN25[1], w661, w662);
  FullAdder U125 (w662, w652, IN26[0], w663, w664);
  HalfAdder U126 (w655, IN22[5], Out1[22], w666);
  FullAdder U127 (w666, w657, IN23[4], w667, w668);
  FullAdder U128 (w668, w659, IN24[3], w669, w670);
  FullAdder U129 (w670, w661, IN25[2], w671, w672);
  FullAdder U130 (w672, w663, IN26[1], w673, w674);
  FullAdder U131 (w674, w664, IN27[0], w675, w676);
  HalfAdder U132 (w667, IN23[5], Out1[23], w678);
  FullAdder U133 (w678, w669, IN24[4], w679, w680);
  FullAdder U134 (w680, w671, IN25[3], w681, w682);
  FullAdder U135 (w682, w673, IN26[2], w683, w684);
  FullAdder U136 (w684, w675, IN27[1], w685, w686);
  FullAdder U137 (w686, w676, IN28[0], w687, w688);
  HalfAdder U138 (w679, IN24[5], Out1[24], w690);
  FullAdder U139 (w690, w681, IN25[4], w691, w692);
  FullAdder U140 (w692, w683, IN26[3], w693, w694);
  FullAdder U141 (w694, w685, IN27[2], w695, w696);
  FullAdder U142 (w696, w687, IN28[1], w697, w698);
  FullAdder U143 (w698, w688, IN29[0], w699, w700);
  HalfAdder U144 (w691, IN25[5], Out1[25], w702);
  FullAdder U145 (w702, w693, IN26[4], w703, w704);
  FullAdder U146 (w704, w695, IN27[3], w705, w706);
  FullAdder U147 (w706, w697, IN28[2], w707, w708);
  FullAdder U148 (w708, w699, IN29[1], w709, w710);
  FullAdder U149 (w710, w700, IN30[0], w711, w712);
  HalfAdder U150 (w703, IN26[5], Out1[26], w714);
  FullAdder U151 (w714, w705, IN27[4], w715, w716);
  FullAdder U152 (w716, w707, IN28[3], w717, w718);
  FullAdder U153 (w718, w709, IN29[2], w719, w720);
  FullAdder U154 (w720, w711, IN30[1], w721, w722);
  FullAdder U155 (w722, w712, IN31[0], w723, w724);
  HalfAdder U156 (w715, IN27[5], Out1[27], w726);
  FullAdder U157 (w726, w717, IN28[4], w727, w728);
  FullAdder U158 (w728, w719, IN29[3], w729, w730);
  FullAdder U159 (w730, w721, IN30[2], w731, w732);
  FullAdder U160 (w732, w723, IN31[1], w733, w734);
  FullAdder U161 (w734, w724, IN32[0], w735, w736);
  HalfAdder U162 (w727, IN28[5], Out1[28], w738);
  FullAdder U163 (w738, w729, IN29[4], w739, w740);
  FullAdder U164 (w740, w731, IN30[3], w741, w742);
  FullAdder U165 (w742, w733, IN31[2], w743, w744);
  FullAdder U166 (w744, w735, IN32[1], w745, w746);
  FullAdder U167 (w746, w736, IN33[0], w747, w748);
  HalfAdder U168 (w739, IN29[5], Out1[29], w750);
  FullAdder U169 (w750, w741, IN30[4], w751, w752);
  FullAdder U170 (w752, w743, IN31[3], w753, w754);
  FullAdder U171 (w754, w745, IN32[2], w755, w756);
  FullAdder U172 (w756, w747, IN33[1], w757, w758);
  FullAdder U173 (w758, w748, IN34[0], w759, w760);
  HalfAdder U174 (w751, IN30[5], Out1[30], w762);
  FullAdder U175 (w762, w753, IN31[4], w763, w764);
  FullAdder U176 (w764, w755, IN32[3], w765, w766);
  FullAdder U177 (w766, w757, IN33[2], w767, w768);
  FullAdder U178 (w768, w759, IN34[1], w769, w770);
  FullAdder U179 (w770, w760, IN35[0], w771, w772);
  HalfAdder U180 (w763, IN31[5], Out1[31], w774);
  FullAdder U181 (w774, w765, IN32[4], w775, w776);
  FullAdder U182 (w776, w767, IN33[3], w777, w778);
  FullAdder U183 (w778, w769, IN34[2], w779, w780);
  FullAdder U184 (w780, w771, IN35[1], w781, w782);
  FullAdder U185 (w782, w772, IN36[0], w783, w784);
  HalfAdder U186 (w775, IN32[5], Out1[32], w786);
  FullAdder U187 (w786, w777, IN33[4], w787, w788);
  FullAdder U188 (w788, w779, IN34[3], w789, w790);
  FullAdder U189 (w790, w781, IN35[2], w791, w792);
  FullAdder U190 (w792, w783, IN36[1], w793, w794);
  FullAdder U191 (w794, w784, IN37[0], w795, w796);
  HalfAdder U192 (w787, IN33[5], Out1[33], w798);
  FullAdder U193 (w798, w789, IN34[4], w799, w800);
  FullAdder U194 (w800, w791, IN35[3], w801, w802);
  FullAdder U195 (w802, w793, IN36[2], w803, w804);
  FullAdder U196 (w804, w795, IN37[1], w805, w806);
  FullAdder U197 (w806, w796, IN38[0], w807, w808);
  HalfAdder U198 (w799, IN34[5], Out1[34], w810);
  FullAdder U199 (w810, w801, IN35[4], w811, w812);
  FullAdder U200 (w812, w803, IN36[3], w813, w814);
  FullAdder U201 (w814, w805, IN37[2], w815, w816);
  FullAdder U202 (w816, w807, IN38[1], w817, w818);
  FullAdder U203 (w818, w808, IN39[0], w819, w820);
  HalfAdder U204 (w811, IN35[5], Out1[35], w822);
  FullAdder U205 (w822, w813, IN36[4], w823, w824);
  FullAdder U206 (w824, w815, IN37[3], w825, w826);
  FullAdder U207 (w826, w817, IN38[2], w827, w828);
  FullAdder U208 (w828, w819, IN39[1], w829, w830);
  FullAdder U209 (w830, w820, IN40[0], w831, w832);
  HalfAdder U210 (w823, IN36[5], Out1[36], w834);
  FullAdder U211 (w834, w825, IN37[4], w835, w836);
  FullAdder U212 (w836, w827, IN38[3], w837, w838);
  FullAdder U213 (w838, w829, IN39[2], w839, w840);
  FullAdder U214 (w840, w831, IN40[1], w841, w842);
  FullAdder U215 (w842, w832, IN41[0], w843, w844);
  HalfAdder U216 (w835, IN37[5], Out1[37], w846);
  FullAdder U217 (w846, w837, IN38[4], w847, w848);
  FullAdder U218 (w848, w839, IN39[3], w849, w850);
  FullAdder U219 (w850, w841, IN40[2], w851, w852);
  FullAdder U220 (w852, w843, IN41[1], w853, w854);
  FullAdder U221 (w854, w844, IN42[0], w855, w856);
  HalfAdder U222 (w847, IN38[5], Out1[38], w858);
  FullAdder U223 (w858, w849, IN39[4], w859, w860);
  FullAdder U224 (w860, w851, IN40[3], w861, w862);
  FullAdder U225 (w862, w853, IN41[2], w863, w864);
  FullAdder U226 (w864, w855, IN42[1], w865, w866);
  FullAdder U227 (w866, w856, IN43[0], w867, w868);
  HalfAdder U228 (w859, IN39[5], Out1[39], w870);
  FullAdder U229 (w870, w861, IN40[4], w871, w872);
  FullAdder U230 (w872, w863, IN41[3], w873, w874);
  FullAdder U231 (w874, w865, IN42[2], w875, w876);
  FullAdder U232 (w876, w867, IN43[1], w877, w878);
  FullAdder U233 (w878, w868, IN44[0], w879, w880);
  HalfAdder U234 (w871, IN40[5], Out1[40], w882);
  FullAdder U235 (w882, w873, IN41[4], w883, w884);
  FullAdder U236 (w884, w875, IN42[3], w885, w886);
  FullAdder U237 (w886, w877, IN43[2], w887, w888);
  FullAdder U238 (w888, w879, IN44[1], w889, w890);
  FullAdder U239 (w890, w880, IN45[0], w891, w892);
  HalfAdder U240 (w883, IN41[5], Out1[41], w894);
  FullAdder U241 (w894, w885, IN42[4], w895, w896);
  FullAdder U242 (w896, w887, IN43[3], w897, w898);
  FullAdder U243 (w898, w889, IN44[2], w899, w900);
  FullAdder U244 (w900, w891, IN45[1], w901, w902);
  FullAdder U245 (w902, w892, IN46[0], w903, w904);
  HalfAdder U246 (w895, IN42[5], Out1[42], w906);
  FullAdder U247 (w906, w897, IN43[4], w907, w908);
  FullAdder U248 (w908, w899, IN44[3], w909, w910);
  FullAdder U249 (w910, w901, IN45[2], w911, w912);
  FullAdder U250 (w912, w903, IN46[1], w913, w914);
  FullAdder U251 (w914, w904, IN47[0], w915, w916);
  HalfAdder U252 (w907, IN43[5], Out1[43], w918);
  FullAdder U253 (w918, w909, IN44[4], w919, w920);
  FullAdder U254 (w920, w911, IN45[3], w921, w922);
  FullAdder U255 (w922, w913, IN46[2], w923, w924);
  FullAdder U256 (w924, w915, IN47[1], w925, w926);
  FullAdder U257 (w926, w916, IN48[0], w927, w928);
  HalfAdder U258 (w919, IN44[5], Out1[44], w930);
  FullAdder U259 (w930, w921, IN45[4], w931, w932);
  FullAdder U260 (w932, w923, IN46[3], w933, w934);
  FullAdder U261 (w934, w925, IN47[2], w935, w936);
  FullAdder U262 (w936, w927, IN48[1], w937, w938);
  FullAdder U263 (w938, w928, IN49[0], w939, w940);
  HalfAdder U264 (w931, IN45[5], Out1[45], w942);
  FullAdder U265 (w942, w933, IN46[4], w943, w944);
  FullAdder U266 (w944, w935, IN47[3], w945, w946);
  FullAdder U267 (w946, w937, IN48[2], w947, w948);
  FullAdder U268 (w948, w939, IN49[1], w949, w950);
  FullAdder U269 (w950, w940, IN50[0], w951, w952);
  HalfAdder U270 (w943, IN46[5], Out1[46], w954);
  FullAdder U271 (w954, w945, IN47[4], w955, w956);
  FullAdder U272 (w956, w947, IN48[3], w957, w958);
  FullAdder U273 (w958, w949, IN49[2], w959, w960);
  FullAdder U274 (w960, w951, IN50[1], w961, w962);
  FullAdder U275 (w962, w952, IN51[0], w963, w964);
  HalfAdder U276 (w955, IN47[5], Out1[47], w966);
  FullAdder U277 (w966, w957, IN48[4], w967, w968);
  FullAdder U278 (w968, w959, IN49[3], w969, w970);
  FullAdder U279 (w970, w961, IN50[2], w971, w972);
  FullAdder U280 (w972, w963, IN51[1], w973, w974);
  FullAdder U281 (w974, w964, IN52[0], w975, w976);
  HalfAdder U282 (w967, IN48[5], Out1[48], w978);
  FullAdder U283 (w978, w969, IN49[4], w979, w980);
  FullAdder U284 (w980, w971, IN50[3], w981, w982);
  FullAdder U285 (w982, w973, IN51[2], w983, w984);
  FullAdder U286 (w984, w975, IN52[1], w985, w986);
  FullAdder U287 (w986, w976, IN53[0], w987, w988);
  HalfAdder U288 (w979, IN49[5], Out1[49], w990);
  FullAdder U289 (w990, w981, IN50[4], w991, w992);
  FullAdder U290 (w992, w983, IN51[3], w993, w994);
  FullAdder U291 (w994, w985, IN52[2], w995, w996);
  FullAdder U292 (w996, w987, IN53[1], w997, w998);
  FullAdder U293 (w998, w988, IN54[0], w999, w1000);
  HalfAdder U294 (w991, IN50[5], Out1[50], w1002);
  FullAdder U295 (w1002, w993, IN51[4], w1003, w1004);
  FullAdder U296 (w1004, w995, IN52[3], w1005, w1006);
  FullAdder U297 (w1006, w997, IN53[2], w1007, w1008);
  FullAdder U298 (w1008, w999, IN54[1], w1009, w1010);
  FullAdder U299 (w1010, w1000, IN55[0], w1011, w1012);
  HalfAdder U300 (w1003, IN51[5], Out1[51], w1014);
  FullAdder U301 (w1014, w1005, IN52[4], w1015, w1016);
  FullAdder U302 (w1016, w1007, IN53[3], w1017, w1018);
  FullAdder U303 (w1018, w1009, IN54[2], w1019, w1020);
  FullAdder U304 (w1020, w1011, IN55[1], w1021, w1022);
  FullAdder U305 (w1022, w1012, IN56[0], w1023, w1024);
  HalfAdder U306 (w1015, IN52[5], Out1[52], w1026);
  FullAdder U307 (w1026, w1017, IN53[4], w1027, w1028);
  FullAdder U308 (w1028, w1019, IN54[3], w1029, w1030);
  FullAdder U309 (w1030, w1021, IN55[2], w1031, w1032);
  FullAdder U310 (w1032, w1023, IN56[1], w1033, w1034);
  FullAdder U311 (w1034, w1024, IN57[0], w1035, w1036);
  HalfAdder U312 (w1027, IN53[5], Out1[53], w1038);
  FullAdder U313 (w1038, w1029, IN54[4], w1039, w1040);
  FullAdder U314 (w1040, w1031, IN55[3], w1041, w1042);
  FullAdder U315 (w1042, w1033, IN56[2], w1043, w1044);
  FullAdder U316 (w1044, w1035, IN57[1], w1045, w1046);
  FullAdder U317 (w1046, w1036, IN58[0], w1047, w1048);
  HalfAdder U318 (w1039, IN54[5], Out1[54], w1050);
  FullAdder U319 (w1050, w1041, IN55[4], w1051, w1052);
  FullAdder U320 (w1052, w1043, IN56[3], w1053, w1054);
  FullAdder U321 (w1054, w1045, IN57[2], w1055, w1056);
  FullAdder U322 (w1056, w1047, IN58[1], w1057, w1058);
  FullAdder U323 (w1058, w1048, IN59[0], w1059, w1060);
  HalfAdder U324 (w1051, IN55[5], Out1[55], w1062);
  FullAdder U325 (w1062, w1053, IN56[4], w1063, w1064);
  FullAdder U326 (w1064, w1055, IN57[3], w1065, w1066);
  FullAdder U327 (w1066, w1057, IN58[2], w1067, w1068);
  FullAdder U328 (w1068, w1059, IN59[1], w1069, w1070);
  FullAdder U329 (w1070, w1060, IN60[0], w1071, w1072);
  HalfAdder U330 (w1063, IN56[5], Out1[56], w1074);
  FullAdder U331 (w1074, w1065, IN57[4], w1075, w1076);
  FullAdder U332 (w1076, w1067, IN58[3], w1077, w1078);
  FullAdder U333 (w1078, w1069, IN59[2], w1079, w1080);
  FullAdder U334 (w1080, w1071, IN60[1], w1081, w1082);
  FullAdder U335 (w1082, w1072, IN61[0], w1083, w1084);
  HalfAdder U336 (w1075, IN57[5], Out1[57], w1086);
  FullAdder U337 (w1086, w1077, IN58[4], w1087, w1088);
  FullAdder U338 (w1088, w1079, IN59[3], w1089, w1090);
  FullAdder U339 (w1090, w1081, IN60[2], w1091, w1092);
  FullAdder U340 (w1092, w1083, IN61[1], w1093, w1094);
  FullAdder U341 (w1094, w1084, IN62[0], w1095, w1096);
  HalfAdder U342 (w1087, IN58[5], Out1[58], w1098);
  FullAdder U343 (w1098, w1089, IN59[4], Out1[59], w1100);
  FullAdder U344 (w1100, w1091, IN60[3], Out1[60], w1102);
  FullAdder U345 (w1102, w1093, IN61[2], Out1[61], w1104);
  FullAdder U346 (w1104, w1095, IN62[1], Out1[62], w1106);
  FullAdder U347 (w1106, w1096, IN63[0], Out1[63], Out1[64]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN7[6];
  assign Out2[1] = IN8[6];
  assign Out2[2] = IN9[6];
  assign Out2[3] = IN10[6];
  assign Out2[4] = IN11[6];
  assign Out2[5] = IN12[6];
  assign Out2[6] = IN13[6];
  assign Out2[7] = IN14[6];
  assign Out2[8] = IN15[6];
  assign Out2[9] = IN16[6];
  assign Out2[10] = IN17[6];
  assign Out2[11] = IN18[6];
  assign Out2[12] = IN19[6];
  assign Out2[13] = IN20[6];
  assign Out2[14] = IN21[6];
  assign Out2[15] = IN22[6];
  assign Out2[16] = IN23[6];
  assign Out2[17] = IN24[6];
  assign Out2[18] = IN25[6];
  assign Out2[19] = IN26[6];
  assign Out2[20] = IN27[6];
  assign Out2[21] = IN28[6];
  assign Out2[22] = IN29[6];
  assign Out2[23] = IN30[6];
  assign Out2[24] = IN31[6];
  assign Out2[25] = IN32[6];
  assign Out2[26] = IN33[6];
  assign Out2[27] = IN34[6];
  assign Out2[28] = IN35[6];
  assign Out2[29] = IN36[6];
  assign Out2[30] = IN37[6];
  assign Out2[31] = IN38[6];
  assign Out2[32] = IN39[6];
  assign Out2[33] = IN40[6];
  assign Out2[34] = IN41[6];
  assign Out2[35] = IN42[6];
  assign Out2[36] = IN43[6];
  assign Out2[37] = IN44[6];
  assign Out2[38] = IN45[6];
  assign Out2[39] = IN46[6];
  assign Out2[40] = IN47[6];
  assign Out2[41] = IN48[6];
  assign Out2[42] = IN49[6];
  assign Out2[43] = IN50[6];
  assign Out2[44] = IN51[6];
  assign Out2[45] = IN52[6];
  assign Out2[46] = IN53[6];
  assign Out2[47] = IN54[6];
  assign Out2[48] = IN55[6];
  assign Out2[49] = IN56[6];
  assign Out2[50] = IN57[6];
  assign Out2[51] = IN58[6];
  assign Out2[52] = IN59[5];
  assign Out2[53] = IN60[4];
  assign Out2[54] = IN61[3];
  assign Out2[55] = IN62[2];
  assign Out2[56] = IN63[1];
  assign Out2[57] = IN64[0];

endmodule
module RC_58_58(IN1, IN2, Out);
  input [57:0] IN1;
  input [57:0] IN2;
  output [58:0] Out;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w117);
  FullAdder U1 (IN1[1], IN2[1], w117, Out[1], w119);
  FullAdder U2 (IN1[2], IN2[2], w119, Out[2], w121);
  FullAdder U3 (IN1[3], IN2[3], w121, Out[3], w123);
  FullAdder U4 (IN1[4], IN2[4], w123, Out[4], w125);
  FullAdder U5 (IN1[5], IN2[5], w125, Out[5], w127);
  FullAdder U6 (IN1[6], IN2[6], w127, Out[6], w129);
  FullAdder U7 (IN1[7], IN2[7], w129, Out[7], w131);
  FullAdder U8 (IN1[8], IN2[8], w131, Out[8], w133);
  FullAdder U9 (IN1[9], IN2[9], w133, Out[9], w135);
  FullAdder U10 (IN1[10], IN2[10], w135, Out[10], w137);
  FullAdder U11 (IN1[11], IN2[11], w137, Out[11], w139);
  FullAdder U12 (IN1[12], IN2[12], w139, Out[12], w141);
  FullAdder U13 (IN1[13], IN2[13], w141, Out[13], w143);
  FullAdder U14 (IN1[14], IN2[14], w143, Out[14], w145);
  FullAdder U15 (IN1[15], IN2[15], w145, Out[15], w147);
  FullAdder U16 (IN1[16], IN2[16], w147, Out[16], w149);
  FullAdder U17 (IN1[17], IN2[17], w149, Out[17], w151);
  FullAdder U18 (IN1[18], IN2[18], w151, Out[18], w153);
  FullAdder U19 (IN1[19], IN2[19], w153, Out[19], w155);
  FullAdder U20 (IN1[20], IN2[20], w155, Out[20], w157);
  FullAdder U21 (IN1[21], IN2[21], w157, Out[21], w159);
  FullAdder U22 (IN1[22], IN2[22], w159, Out[22], w161);
  FullAdder U23 (IN1[23], IN2[23], w161, Out[23], w163);
  FullAdder U24 (IN1[24], IN2[24], w163, Out[24], w165);
  FullAdder U25 (IN1[25], IN2[25], w165, Out[25], w167);
  FullAdder U26 (IN1[26], IN2[26], w167, Out[26], w169);
  FullAdder U27 (IN1[27], IN2[27], w169, Out[27], w171);
  FullAdder U28 (IN1[28], IN2[28], w171, Out[28], w173);
  FullAdder U29 (IN1[29], IN2[29], w173, Out[29], w175);
  FullAdder U30 (IN1[30], IN2[30], w175, Out[30], w177);
  FullAdder U31 (IN1[31], IN2[31], w177, Out[31], w179);
  FullAdder U32 (IN1[32], IN2[32], w179, Out[32], w181);
  FullAdder U33 (IN1[33], IN2[33], w181, Out[33], w183);
  FullAdder U34 (IN1[34], IN2[34], w183, Out[34], w185);
  FullAdder U35 (IN1[35], IN2[35], w185, Out[35], w187);
  FullAdder U36 (IN1[36], IN2[36], w187, Out[36], w189);
  FullAdder U37 (IN1[37], IN2[37], w189, Out[37], w191);
  FullAdder U38 (IN1[38], IN2[38], w191, Out[38], w193);
  FullAdder U39 (IN1[39], IN2[39], w193, Out[39], w195);
  FullAdder U40 (IN1[40], IN2[40], w195, Out[40], w197);
  FullAdder U41 (IN1[41], IN2[41], w197, Out[41], w199);
  FullAdder U42 (IN1[42], IN2[42], w199, Out[42], w201);
  FullAdder U43 (IN1[43], IN2[43], w201, Out[43], w203);
  FullAdder U44 (IN1[44], IN2[44], w203, Out[44], w205);
  FullAdder U45 (IN1[45], IN2[45], w205, Out[45], w207);
  FullAdder U46 (IN1[46], IN2[46], w207, Out[46], w209);
  FullAdder U47 (IN1[47], IN2[47], w209, Out[47], w211);
  FullAdder U48 (IN1[48], IN2[48], w211, Out[48], w213);
  FullAdder U49 (IN1[49], IN2[49], w213, Out[49], w215);
  FullAdder U50 (IN1[50], IN2[50], w215, Out[50], w217);
  FullAdder U51 (IN1[51], IN2[51], w217, Out[51], w219);
  FullAdder U52 (IN1[52], IN2[52], w219, Out[52], w221);
  FullAdder U53 (IN1[53], IN2[53], w221, Out[53], w223);
  FullAdder U54 (IN1[54], IN2[54], w223, Out[54], w225);
  FullAdder U55 (IN1[55], IN2[55], w225, Out[55], w227);
  FullAdder U56 (IN1[56], IN2[56], w227, Out[56], w229);
  FullAdder U57 (IN1[57], IN2[57], w229, Out[57], Out[58]);

endmodule
module NR_7_59(IN1, IN2, Out);
  input [6:0] IN1;
  input [58:0] IN2;
  output [65:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [6:0] P37;
  wire [6:0] P38;
  wire [6:0] P39;
  wire [6:0] P40;
  wire [6:0] P41;
  wire [6:0] P42;
  wire [6:0] P43;
  wire [6:0] P44;
  wire [6:0] P45;
  wire [6:0] P46;
  wire [6:0] P47;
  wire [6:0] P48;
  wire [6:0] P49;
  wire [6:0] P50;
  wire [6:0] P51;
  wire [6:0] P52;
  wire [6:0] P53;
  wire [6:0] P54;
  wire [6:0] P55;
  wire [6:0] P56;
  wire [6:0] P57;
  wire [6:0] P58;
  wire [5:0] P59;
  wire [4:0] P60;
  wire [3:0] P61;
  wire [2:0] P62;
  wire [1:0] P63;
  wire [0:0] P64;
  wire [64:0] R1;
  wire [57:0] R2;
  wire [65:0] aOut;
  U_SP_7_59 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, R1, R2);
  RC_58_58 S2 (R1[64:7], R2, aOut[65:7]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign Out = aOut[65:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
