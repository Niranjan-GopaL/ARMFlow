
module customAdder43_0(
    input [42 : 0] A,
    input [42 : 0] B,
    output [43 : 0] Sum
);

    assign Sum = A+B;

endmodule
