
module NR_1_52(
    input [0:0]IN1,
    input [51:0]IN2,
    output [51:0]Out
);
    assign Out = IN2;
endmodule
