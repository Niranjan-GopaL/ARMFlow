
module NR_39_1(
    input [38:0]IN1,
    input [0:0]IN2,
    output [38:0]Out
);
    assign Out = IN2;
endmodule
