//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 59
  second input length: 21
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_59_21(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78);
  input [58:0] IN1;
  input [20:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [20:0] P21;
  output [20:0] P22;
  output [20:0] P23;
  output [20:0] P24;
  output [20:0] P25;
  output [20:0] P26;
  output [20:0] P27;
  output [20:0] P28;
  output [20:0] P29;
  output [20:0] P30;
  output [20:0] P31;
  output [20:0] P32;
  output [20:0] P33;
  output [20:0] P34;
  output [20:0] P35;
  output [20:0] P36;
  output [20:0] P37;
  output [20:0] P38;
  output [20:0] P39;
  output [20:0] P40;
  output [20:0] P41;
  output [20:0] P42;
  output [20:0] P43;
  output [20:0] P44;
  output [20:0] P45;
  output [20:0] P46;
  output [20:0] P47;
  output [20:0] P48;
  output [20:0] P49;
  output [20:0] P50;
  output [20:0] P51;
  output [20:0] P52;
  output [20:0] P53;
  output [20:0] P54;
  output [20:0] P55;
  output [20:0] P56;
  output [20:0] P57;
  output [20:0] P58;
  output [19:0] P59;
  output [18:0] P60;
  output [17:0] P61;
  output [16:0] P62;
  output [15:0] P63;
  output [14:0] P64;
  output [13:0] P65;
  output [12:0] P66;
  output [11:0] P67;
  output [10:0] P68;
  output [9:0] P69;
  output [8:0] P70;
  output [7:0] P71;
  output [6:0] P72;
  output [5:0] P73;
  output [4:0] P74;
  output [3:0] P75;
  output [2:0] P76;
  output [1:0] P77;
  output [0:0] P78;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[0] = IN1[1]&IN2[20];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[1] = IN1[2]&IN2[19];
  assign P22[0] = IN1[2]&IN2[20];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[2] = IN1[3]&IN2[18];
  assign P22[1] = IN1[3]&IN2[19];
  assign P23[0] = IN1[3]&IN2[20];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[3] = IN1[4]&IN2[17];
  assign P22[2] = IN1[4]&IN2[18];
  assign P23[1] = IN1[4]&IN2[19];
  assign P24[0] = IN1[4]&IN2[20];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[4] = IN1[5]&IN2[16];
  assign P22[3] = IN1[5]&IN2[17];
  assign P23[2] = IN1[5]&IN2[18];
  assign P24[1] = IN1[5]&IN2[19];
  assign P25[0] = IN1[5]&IN2[20];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[5] = IN1[6]&IN2[15];
  assign P22[4] = IN1[6]&IN2[16];
  assign P23[3] = IN1[6]&IN2[17];
  assign P24[2] = IN1[6]&IN2[18];
  assign P25[1] = IN1[6]&IN2[19];
  assign P26[0] = IN1[6]&IN2[20];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[6] = IN1[7]&IN2[14];
  assign P22[5] = IN1[7]&IN2[15];
  assign P23[4] = IN1[7]&IN2[16];
  assign P24[3] = IN1[7]&IN2[17];
  assign P25[2] = IN1[7]&IN2[18];
  assign P26[1] = IN1[7]&IN2[19];
  assign P27[0] = IN1[7]&IN2[20];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[7] = IN1[8]&IN2[13];
  assign P22[6] = IN1[8]&IN2[14];
  assign P23[5] = IN1[8]&IN2[15];
  assign P24[4] = IN1[8]&IN2[16];
  assign P25[3] = IN1[8]&IN2[17];
  assign P26[2] = IN1[8]&IN2[18];
  assign P27[1] = IN1[8]&IN2[19];
  assign P28[0] = IN1[8]&IN2[20];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[8] = IN1[9]&IN2[12];
  assign P22[7] = IN1[9]&IN2[13];
  assign P23[6] = IN1[9]&IN2[14];
  assign P24[5] = IN1[9]&IN2[15];
  assign P25[4] = IN1[9]&IN2[16];
  assign P26[3] = IN1[9]&IN2[17];
  assign P27[2] = IN1[9]&IN2[18];
  assign P28[1] = IN1[9]&IN2[19];
  assign P29[0] = IN1[9]&IN2[20];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[9] = IN1[10]&IN2[11];
  assign P22[8] = IN1[10]&IN2[12];
  assign P23[7] = IN1[10]&IN2[13];
  assign P24[6] = IN1[10]&IN2[14];
  assign P25[5] = IN1[10]&IN2[15];
  assign P26[4] = IN1[10]&IN2[16];
  assign P27[3] = IN1[10]&IN2[17];
  assign P28[2] = IN1[10]&IN2[18];
  assign P29[1] = IN1[10]&IN2[19];
  assign P30[0] = IN1[10]&IN2[20];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[10] = IN1[11]&IN2[10];
  assign P22[9] = IN1[11]&IN2[11];
  assign P23[8] = IN1[11]&IN2[12];
  assign P24[7] = IN1[11]&IN2[13];
  assign P25[6] = IN1[11]&IN2[14];
  assign P26[5] = IN1[11]&IN2[15];
  assign P27[4] = IN1[11]&IN2[16];
  assign P28[3] = IN1[11]&IN2[17];
  assign P29[2] = IN1[11]&IN2[18];
  assign P30[1] = IN1[11]&IN2[19];
  assign P31[0] = IN1[11]&IN2[20];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[11] = IN1[12]&IN2[9];
  assign P22[10] = IN1[12]&IN2[10];
  assign P23[9] = IN1[12]&IN2[11];
  assign P24[8] = IN1[12]&IN2[12];
  assign P25[7] = IN1[12]&IN2[13];
  assign P26[6] = IN1[12]&IN2[14];
  assign P27[5] = IN1[12]&IN2[15];
  assign P28[4] = IN1[12]&IN2[16];
  assign P29[3] = IN1[12]&IN2[17];
  assign P30[2] = IN1[12]&IN2[18];
  assign P31[1] = IN1[12]&IN2[19];
  assign P32[0] = IN1[12]&IN2[20];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[12] = IN1[13]&IN2[8];
  assign P22[11] = IN1[13]&IN2[9];
  assign P23[10] = IN1[13]&IN2[10];
  assign P24[9] = IN1[13]&IN2[11];
  assign P25[8] = IN1[13]&IN2[12];
  assign P26[7] = IN1[13]&IN2[13];
  assign P27[6] = IN1[13]&IN2[14];
  assign P28[5] = IN1[13]&IN2[15];
  assign P29[4] = IN1[13]&IN2[16];
  assign P30[3] = IN1[13]&IN2[17];
  assign P31[2] = IN1[13]&IN2[18];
  assign P32[1] = IN1[13]&IN2[19];
  assign P33[0] = IN1[13]&IN2[20];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[13] = IN1[14]&IN2[7];
  assign P22[12] = IN1[14]&IN2[8];
  assign P23[11] = IN1[14]&IN2[9];
  assign P24[10] = IN1[14]&IN2[10];
  assign P25[9] = IN1[14]&IN2[11];
  assign P26[8] = IN1[14]&IN2[12];
  assign P27[7] = IN1[14]&IN2[13];
  assign P28[6] = IN1[14]&IN2[14];
  assign P29[5] = IN1[14]&IN2[15];
  assign P30[4] = IN1[14]&IN2[16];
  assign P31[3] = IN1[14]&IN2[17];
  assign P32[2] = IN1[14]&IN2[18];
  assign P33[1] = IN1[14]&IN2[19];
  assign P34[0] = IN1[14]&IN2[20];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[14] = IN1[15]&IN2[6];
  assign P22[13] = IN1[15]&IN2[7];
  assign P23[12] = IN1[15]&IN2[8];
  assign P24[11] = IN1[15]&IN2[9];
  assign P25[10] = IN1[15]&IN2[10];
  assign P26[9] = IN1[15]&IN2[11];
  assign P27[8] = IN1[15]&IN2[12];
  assign P28[7] = IN1[15]&IN2[13];
  assign P29[6] = IN1[15]&IN2[14];
  assign P30[5] = IN1[15]&IN2[15];
  assign P31[4] = IN1[15]&IN2[16];
  assign P32[3] = IN1[15]&IN2[17];
  assign P33[2] = IN1[15]&IN2[18];
  assign P34[1] = IN1[15]&IN2[19];
  assign P35[0] = IN1[15]&IN2[20];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[15] = IN1[16]&IN2[5];
  assign P22[14] = IN1[16]&IN2[6];
  assign P23[13] = IN1[16]&IN2[7];
  assign P24[12] = IN1[16]&IN2[8];
  assign P25[11] = IN1[16]&IN2[9];
  assign P26[10] = IN1[16]&IN2[10];
  assign P27[9] = IN1[16]&IN2[11];
  assign P28[8] = IN1[16]&IN2[12];
  assign P29[7] = IN1[16]&IN2[13];
  assign P30[6] = IN1[16]&IN2[14];
  assign P31[5] = IN1[16]&IN2[15];
  assign P32[4] = IN1[16]&IN2[16];
  assign P33[3] = IN1[16]&IN2[17];
  assign P34[2] = IN1[16]&IN2[18];
  assign P35[1] = IN1[16]&IN2[19];
  assign P36[0] = IN1[16]&IN2[20];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[16] = IN1[17]&IN2[4];
  assign P22[15] = IN1[17]&IN2[5];
  assign P23[14] = IN1[17]&IN2[6];
  assign P24[13] = IN1[17]&IN2[7];
  assign P25[12] = IN1[17]&IN2[8];
  assign P26[11] = IN1[17]&IN2[9];
  assign P27[10] = IN1[17]&IN2[10];
  assign P28[9] = IN1[17]&IN2[11];
  assign P29[8] = IN1[17]&IN2[12];
  assign P30[7] = IN1[17]&IN2[13];
  assign P31[6] = IN1[17]&IN2[14];
  assign P32[5] = IN1[17]&IN2[15];
  assign P33[4] = IN1[17]&IN2[16];
  assign P34[3] = IN1[17]&IN2[17];
  assign P35[2] = IN1[17]&IN2[18];
  assign P36[1] = IN1[17]&IN2[19];
  assign P37[0] = IN1[17]&IN2[20];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[17] = IN1[18]&IN2[3];
  assign P22[16] = IN1[18]&IN2[4];
  assign P23[15] = IN1[18]&IN2[5];
  assign P24[14] = IN1[18]&IN2[6];
  assign P25[13] = IN1[18]&IN2[7];
  assign P26[12] = IN1[18]&IN2[8];
  assign P27[11] = IN1[18]&IN2[9];
  assign P28[10] = IN1[18]&IN2[10];
  assign P29[9] = IN1[18]&IN2[11];
  assign P30[8] = IN1[18]&IN2[12];
  assign P31[7] = IN1[18]&IN2[13];
  assign P32[6] = IN1[18]&IN2[14];
  assign P33[5] = IN1[18]&IN2[15];
  assign P34[4] = IN1[18]&IN2[16];
  assign P35[3] = IN1[18]&IN2[17];
  assign P36[2] = IN1[18]&IN2[18];
  assign P37[1] = IN1[18]&IN2[19];
  assign P38[0] = IN1[18]&IN2[20];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[18] = IN1[19]&IN2[2];
  assign P22[17] = IN1[19]&IN2[3];
  assign P23[16] = IN1[19]&IN2[4];
  assign P24[15] = IN1[19]&IN2[5];
  assign P25[14] = IN1[19]&IN2[6];
  assign P26[13] = IN1[19]&IN2[7];
  assign P27[12] = IN1[19]&IN2[8];
  assign P28[11] = IN1[19]&IN2[9];
  assign P29[10] = IN1[19]&IN2[10];
  assign P30[9] = IN1[19]&IN2[11];
  assign P31[8] = IN1[19]&IN2[12];
  assign P32[7] = IN1[19]&IN2[13];
  assign P33[6] = IN1[19]&IN2[14];
  assign P34[5] = IN1[19]&IN2[15];
  assign P35[4] = IN1[19]&IN2[16];
  assign P36[3] = IN1[19]&IN2[17];
  assign P37[2] = IN1[19]&IN2[18];
  assign P38[1] = IN1[19]&IN2[19];
  assign P39[0] = IN1[19]&IN2[20];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[19] = IN1[20]&IN2[1];
  assign P22[18] = IN1[20]&IN2[2];
  assign P23[17] = IN1[20]&IN2[3];
  assign P24[16] = IN1[20]&IN2[4];
  assign P25[15] = IN1[20]&IN2[5];
  assign P26[14] = IN1[20]&IN2[6];
  assign P27[13] = IN1[20]&IN2[7];
  assign P28[12] = IN1[20]&IN2[8];
  assign P29[11] = IN1[20]&IN2[9];
  assign P30[10] = IN1[20]&IN2[10];
  assign P31[9] = IN1[20]&IN2[11];
  assign P32[8] = IN1[20]&IN2[12];
  assign P33[7] = IN1[20]&IN2[13];
  assign P34[6] = IN1[20]&IN2[14];
  assign P35[5] = IN1[20]&IN2[15];
  assign P36[4] = IN1[20]&IN2[16];
  assign P37[3] = IN1[20]&IN2[17];
  assign P38[2] = IN1[20]&IN2[18];
  assign P39[1] = IN1[20]&IN2[19];
  assign P40[0] = IN1[20]&IN2[20];
  assign P21[20] = IN1[21]&IN2[0];
  assign P22[19] = IN1[21]&IN2[1];
  assign P23[18] = IN1[21]&IN2[2];
  assign P24[17] = IN1[21]&IN2[3];
  assign P25[16] = IN1[21]&IN2[4];
  assign P26[15] = IN1[21]&IN2[5];
  assign P27[14] = IN1[21]&IN2[6];
  assign P28[13] = IN1[21]&IN2[7];
  assign P29[12] = IN1[21]&IN2[8];
  assign P30[11] = IN1[21]&IN2[9];
  assign P31[10] = IN1[21]&IN2[10];
  assign P32[9] = IN1[21]&IN2[11];
  assign P33[8] = IN1[21]&IN2[12];
  assign P34[7] = IN1[21]&IN2[13];
  assign P35[6] = IN1[21]&IN2[14];
  assign P36[5] = IN1[21]&IN2[15];
  assign P37[4] = IN1[21]&IN2[16];
  assign P38[3] = IN1[21]&IN2[17];
  assign P39[2] = IN1[21]&IN2[18];
  assign P40[1] = IN1[21]&IN2[19];
  assign P41[0] = IN1[21]&IN2[20];
  assign P22[20] = IN1[22]&IN2[0];
  assign P23[19] = IN1[22]&IN2[1];
  assign P24[18] = IN1[22]&IN2[2];
  assign P25[17] = IN1[22]&IN2[3];
  assign P26[16] = IN1[22]&IN2[4];
  assign P27[15] = IN1[22]&IN2[5];
  assign P28[14] = IN1[22]&IN2[6];
  assign P29[13] = IN1[22]&IN2[7];
  assign P30[12] = IN1[22]&IN2[8];
  assign P31[11] = IN1[22]&IN2[9];
  assign P32[10] = IN1[22]&IN2[10];
  assign P33[9] = IN1[22]&IN2[11];
  assign P34[8] = IN1[22]&IN2[12];
  assign P35[7] = IN1[22]&IN2[13];
  assign P36[6] = IN1[22]&IN2[14];
  assign P37[5] = IN1[22]&IN2[15];
  assign P38[4] = IN1[22]&IN2[16];
  assign P39[3] = IN1[22]&IN2[17];
  assign P40[2] = IN1[22]&IN2[18];
  assign P41[1] = IN1[22]&IN2[19];
  assign P42[0] = IN1[22]&IN2[20];
  assign P23[20] = IN1[23]&IN2[0];
  assign P24[19] = IN1[23]&IN2[1];
  assign P25[18] = IN1[23]&IN2[2];
  assign P26[17] = IN1[23]&IN2[3];
  assign P27[16] = IN1[23]&IN2[4];
  assign P28[15] = IN1[23]&IN2[5];
  assign P29[14] = IN1[23]&IN2[6];
  assign P30[13] = IN1[23]&IN2[7];
  assign P31[12] = IN1[23]&IN2[8];
  assign P32[11] = IN1[23]&IN2[9];
  assign P33[10] = IN1[23]&IN2[10];
  assign P34[9] = IN1[23]&IN2[11];
  assign P35[8] = IN1[23]&IN2[12];
  assign P36[7] = IN1[23]&IN2[13];
  assign P37[6] = IN1[23]&IN2[14];
  assign P38[5] = IN1[23]&IN2[15];
  assign P39[4] = IN1[23]&IN2[16];
  assign P40[3] = IN1[23]&IN2[17];
  assign P41[2] = IN1[23]&IN2[18];
  assign P42[1] = IN1[23]&IN2[19];
  assign P43[0] = IN1[23]&IN2[20];
  assign P24[20] = IN1[24]&IN2[0];
  assign P25[19] = IN1[24]&IN2[1];
  assign P26[18] = IN1[24]&IN2[2];
  assign P27[17] = IN1[24]&IN2[3];
  assign P28[16] = IN1[24]&IN2[4];
  assign P29[15] = IN1[24]&IN2[5];
  assign P30[14] = IN1[24]&IN2[6];
  assign P31[13] = IN1[24]&IN2[7];
  assign P32[12] = IN1[24]&IN2[8];
  assign P33[11] = IN1[24]&IN2[9];
  assign P34[10] = IN1[24]&IN2[10];
  assign P35[9] = IN1[24]&IN2[11];
  assign P36[8] = IN1[24]&IN2[12];
  assign P37[7] = IN1[24]&IN2[13];
  assign P38[6] = IN1[24]&IN2[14];
  assign P39[5] = IN1[24]&IN2[15];
  assign P40[4] = IN1[24]&IN2[16];
  assign P41[3] = IN1[24]&IN2[17];
  assign P42[2] = IN1[24]&IN2[18];
  assign P43[1] = IN1[24]&IN2[19];
  assign P44[0] = IN1[24]&IN2[20];
  assign P25[20] = IN1[25]&IN2[0];
  assign P26[19] = IN1[25]&IN2[1];
  assign P27[18] = IN1[25]&IN2[2];
  assign P28[17] = IN1[25]&IN2[3];
  assign P29[16] = IN1[25]&IN2[4];
  assign P30[15] = IN1[25]&IN2[5];
  assign P31[14] = IN1[25]&IN2[6];
  assign P32[13] = IN1[25]&IN2[7];
  assign P33[12] = IN1[25]&IN2[8];
  assign P34[11] = IN1[25]&IN2[9];
  assign P35[10] = IN1[25]&IN2[10];
  assign P36[9] = IN1[25]&IN2[11];
  assign P37[8] = IN1[25]&IN2[12];
  assign P38[7] = IN1[25]&IN2[13];
  assign P39[6] = IN1[25]&IN2[14];
  assign P40[5] = IN1[25]&IN2[15];
  assign P41[4] = IN1[25]&IN2[16];
  assign P42[3] = IN1[25]&IN2[17];
  assign P43[2] = IN1[25]&IN2[18];
  assign P44[1] = IN1[25]&IN2[19];
  assign P45[0] = IN1[25]&IN2[20];
  assign P26[20] = IN1[26]&IN2[0];
  assign P27[19] = IN1[26]&IN2[1];
  assign P28[18] = IN1[26]&IN2[2];
  assign P29[17] = IN1[26]&IN2[3];
  assign P30[16] = IN1[26]&IN2[4];
  assign P31[15] = IN1[26]&IN2[5];
  assign P32[14] = IN1[26]&IN2[6];
  assign P33[13] = IN1[26]&IN2[7];
  assign P34[12] = IN1[26]&IN2[8];
  assign P35[11] = IN1[26]&IN2[9];
  assign P36[10] = IN1[26]&IN2[10];
  assign P37[9] = IN1[26]&IN2[11];
  assign P38[8] = IN1[26]&IN2[12];
  assign P39[7] = IN1[26]&IN2[13];
  assign P40[6] = IN1[26]&IN2[14];
  assign P41[5] = IN1[26]&IN2[15];
  assign P42[4] = IN1[26]&IN2[16];
  assign P43[3] = IN1[26]&IN2[17];
  assign P44[2] = IN1[26]&IN2[18];
  assign P45[1] = IN1[26]&IN2[19];
  assign P46[0] = IN1[26]&IN2[20];
  assign P27[20] = IN1[27]&IN2[0];
  assign P28[19] = IN1[27]&IN2[1];
  assign P29[18] = IN1[27]&IN2[2];
  assign P30[17] = IN1[27]&IN2[3];
  assign P31[16] = IN1[27]&IN2[4];
  assign P32[15] = IN1[27]&IN2[5];
  assign P33[14] = IN1[27]&IN2[6];
  assign P34[13] = IN1[27]&IN2[7];
  assign P35[12] = IN1[27]&IN2[8];
  assign P36[11] = IN1[27]&IN2[9];
  assign P37[10] = IN1[27]&IN2[10];
  assign P38[9] = IN1[27]&IN2[11];
  assign P39[8] = IN1[27]&IN2[12];
  assign P40[7] = IN1[27]&IN2[13];
  assign P41[6] = IN1[27]&IN2[14];
  assign P42[5] = IN1[27]&IN2[15];
  assign P43[4] = IN1[27]&IN2[16];
  assign P44[3] = IN1[27]&IN2[17];
  assign P45[2] = IN1[27]&IN2[18];
  assign P46[1] = IN1[27]&IN2[19];
  assign P47[0] = IN1[27]&IN2[20];
  assign P28[20] = IN1[28]&IN2[0];
  assign P29[19] = IN1[28]&IN2[1];
  assign P30[18] = IN1[28]&IN2[2];
  assign P31[17] = IN1[28]&IN2[3];
  assign P32[16] = IN1[28]&IN2[4];
  assign P33[15] = IN1[28]&IN2[5];
  assign P34[14] = IN1[28]&IN2[6];
  assign P35[13] = IN1[28]&IN2[7];
  assign P36[12] = IN1[28]&IN2[8];
  assign P37[11] = IN1[28]&IN2[9];
  assign P38[10] = IN1[28]&IN2[10];
  assign P39[9] = IN1[28]&IN2[11];
  assign P40[8] = IN1[28]&IN2[12];
  assign P41[7] = IN1[28]&IN2[13];
  assign P42[6] = IN1[28]&IN2[14];
  assign P43[5] = IN1[28]&IN2[15];
  assign P44[4] = IN1[28]&IN2[16];
  assign P45[3] = IN1[28]&IN2[17];
  assign P46[2] = IN1[28]&IN2[18];
  assign P47[1] = IN1[28]&IN2[19];
  assign P48[0] = IN1[28]&IN2[20];
  assign P29[20] = IN1[29]&IN2[0];
  assign P30[19] = IN1[29]&IN2[1];
  assign P31[18] = IN1[29]&IN2[2];
  assign P32[17] = IN1[29]&IN2[3];
  assign P33[16] = IN1[29]&IN2[4];
  assign P34[15] = IN1[29]&IN2[5];
  assign P35[14] = IN1[29]&IN2[6];
  assign P36[13] = IN1[29]&IN2[7];
  assign P37[12] = IN1[29]&IN2[8];
  assign P38[11] = IN1[29]&IN2[9];
  assign P39[10] = IN1[29]&IN2[10];
  assign P40[9] = IN1[29]&IN2[11];
  assign P41[8] = IN1[29]&IN2[12];
  assign P42[7] = IN1[29]&IN2[13];
  assign P43[6] = IN1[29]&IN2[14];
  assign P44[5] = IN1[29]&IN2[15];
  assign P45[4] = IN1[29]&IN2[16];
  assign P46[3] = IN1[29]&IN2[17];
  assign P47[2] = IN1[29]&IN2[18];
  assign P48[1] = IN1[29]&IN2[19];
  assign P49[0] = IN1[29]&IN2[20];
  assign P30[20] = IN1[30]&IN2[0];
  assign P31[19] = IN1[30]&IN2[1];
  assign P32[18] = IN1[30]&IN2[2];
  assign P33[17] = IN1[30]&IN2[3];
  assign P34[16] = IN1[30]&IN2[4];
  assign P35[15] = IN1[30]&IN2[5];
  assign P36[14] = IN1[30]&IN2[6];
  assign P37[13] = IN1[30]&IN2[7];
  assign P38[12] = IN1[30]&IN2[8];
  assign P39[11] = IN1[30]&IN2[9];
  assign P40[10] = IN1[30]&IN2[10];
  assign P41[9] = IN1[30]&IN2[11];
  assign P42[8] = IN1[30]&IN2[12];
  assign P43[7] = IN1[30]&IN2[13];
  assign P44[6] = IN1[30]&IN2[14];
  assign P45[5] = IN1[30]&IN2[15];
  assign P46[4] = IN1[30]&IN2[16];
  assign P47[3] = IN1[30]&IN2[17];
  assign P48[2] = IN1[30]&IN2[18];
  assign P49[1] = IN1[30]&IN2[19];
  assign P50[0] = IN1[30]&IN2[20];
  assign P31[20] = IN1[31]&IN2[0];
  assign P32[19] = IN1[31]&IN2[1];
  assign P33[18] = IN1[31]&IN2[2];
  assign P34[17] = IN1[31]&IN2[3];
  assign P35[16] = IN1[31]&IN2[4];
  assign P36[15] = IN1[31]&IN2[5];
  assign P37[14] = IN1[31]&IN2[6];
  assign P38[13] = IN1[31]&IN2[7];
  assign P39[12] = IN1[31]&IN2[8];
  assign P40[11] = IN1[31]&IN2[9];
  assign P41[10] = IN1[31]&IN2[10];
  assign P42[9] = IN1[31]&IN2[11];
  assign P43[8] = IN1[31]&IN2[12];
  assign P44[7] = IN1[31]&IN2[13];
  assign P45[6] = IN1[31]&IN2[14];
  assign P46[5] = IN1[31]&IN2[15];
  assign P47[4] = IN1[31]&IN2[16];
  assign P48[3] = IN1[31]&IN2[17];
  assign P49[2] = IN1[31]&IN2[18];
  assign P50[1] = IN1[31]&IN2[19];
  assign P51[0] = IN1[31]&IN2[20];
  assign P32[20] = IN1[32]&IN2[0];
  assign P33[19] = IN1[32]&IN2[1];
  assign P34[18] = IN1[32]&IN2[2];
  assign P35[17] = IN1[32]&IN2[3];
  assign P36[16] = IN1[32]&IN2[4];
  assign P37[15] = IN1[32]&IN2[5];
  assign P38[14] = IN1[32]&IN2[6];
  assign P39[13] = IN1[32]&IN2[7];
  assign P40[12] = IN1[32]&IN2[8];
  assign P41[11] = IN1[32]&IN2[9];
  assign P42[10] = IN1[32]&IN2[10];
  assign P43[9] = IN1[32]&IN2[11];
  assign P44[8] = IN1[32]&IN2[12];
  assign P45[7] = IN1[32]&IN2[13];
  assign P46[6] = IN1[32]&IN2[14];
  assign P47[5] = IN1[32]&IN2[15];
  assign P48[4] = IN1[32]&IN2[16];
  assign P49[3] = IN1[32]&IN2[17];
  assign P50[2] = IN1[32]&IN2[18];
  assign P51[1] = IN1[32]&IN2[19];
  assign P52[0] = IN1[32]&IN2[20];
  assign P33[20] = IN1[33]&IN2[0];
  assign P34[19] = IN1[33]&IN2[1];
  assign P35[18] = IN1[33]&IN2[2];
  assign P36[17] = IN1[33]&IN2[3];
  assign P37[16] = IN1[33]&IN2[4];
  assign P38[15] = IN1[33]&IN2[5];
  assign P39[14] = IN1[33]&IN2[6];
  assign P40[13] = IN1[33]&IN2[7];
  assign P41[12] = IN1[33]&IN2[8];
  assign P42[11] = IN1[33]&IN2[9];
  assign P43[10] = IN1[33]&IN2[10];
  assign P44[9] = IN1[33]&IN2[11];
  assign P45[8] = IN1[33]&IN2[12];
  assign P46[7] = IN1[33]&IN2[13];
  assign P47[6] = IN1[33]&IN2[14];
  assign P48[5] = IN1[33]&IN2[15];
  assign P49[4] = IN1[33]&IN2[16];
  assign P50[3] = IN1[33]&IN2[17];
  assign P51[2] = IN1[33]&IN2[18];
  assign P52[1] = IN1[33]&IN2[19];
  assign P53[0] = IN1[33]&IN2[20];
  assign P34[20] = IN1[34]&IN2[0];
  assign P35[19] = IN1[34]&IN2[1];
  assign P36[18] = IN1[34]&IN2[2];
  assign P37[17] = IN1[34]&IN2[3];
  assign P38[16] = IN1[34]&IN2[4];
  assign P39[15] = IN1[34]&IN2[5];
  assign P40[14] = IN1[34]&IN2[6];
  assign P41[13] = IN1[34]&IN2[7];
  assign P42[12] = IN1[34]&IN2[8];
  assign P43[11] = IN1[34]&IN2[9];
  assign P44[10] = IN1[34]&IN2[10];
  assign P45[9] = IN1[34]&IN2[11];
  assign P46[8] = IN1[34]&IN2[12];
  assign P47[7] = IN1[34]&IN2[13];
  assign P48[6] = IN1[34]&IN2[14];
  assign P49[5] = IN1[34]&IN2[15];
  assign P50[4] = IN1[34]&IN2[16];
  assign P51[3] = IN1[34]&IN2[17];
  assign P52[2] = IN1[34]&IN2[18];
  assign P53[1] = IN1[34]&IN2[19];
  assign P54[0] = IN1[34]&IN2[20];
  assign P35[20] = IN1[35]&IN2[0];
  assign P36[19] = IN1[35]&IN2[1];
  assign P37[18] = IN1[35]&IN2[2];
  assign P38[17] = IN1[35]&IN2[3];
  assign P39[16] = IN1[35]&IN2[4];
  assign P40[15] = IN1[35]&IN2[5];
  assign P41[14] = IN1[35]&IN2[6];
  assign P42[13] = IN1[35]&IN2[7];
  assign P43[12] = IN1[35]&IN2[8];
  assign P44[11] = IN1[35]&IN2[9];
  assign P45[10] = IN1[35]&IN2[10];
  assign P46[9] = IN1[35]&IN2[11];
  assign P47[8] = IN1[35]&IN2[12];
  assign P48[7] = IN1[35]&IN2[13];
  assign P49[6] = IN1[35]&IN2[14];
  assign P50[5] = IN1[35]&IN2[15];
  assign P51[4] = IN1[35]&IN2[16];
  assign P52[3] = IN1[35]&IN2[17];
  assign P53[2] = IN1[35]&IN2[18];
  assign P54[1] = IN1[35]&IN2[19];
  assign P55[0] = IN1[35]&IN2[20];
  assign P36[20] = IN1[36]&IN2[0];
  assign P37[19] = IN1[36]&IN2[1];
  assign P38[18] = IN1[36]&IN2[2];
  assign P39[17] = IN1[36]&IN2[3];
  assign P40[16] = IN1[36]&IN2[4];
  assign P41[15] = IN1[36]&IN2[5];
  assign P42[14] = IN1[36]&IN2[6];
  assign P43[13] = IN1[36]&IN2[7];
  assign P44[12] = IN1[36]&IN2[8];
  assign P45[11] = IN1[36]&IN2[9];
  assign P46[10] = IN1[36]&IN2[10];
  assign P47[9] = IN1[36]&IN2[11];
  assign P48[8] = IN1[36]&IN2[12];
  assign P49[7] = IN1[36]&IN2[13];
  assign P50[6] = IN1[36]&IN2[14];
  assign P51[5] = IN1[36]&IN2[15];
  assign P52[4] = IN1[36]&IN2[16];
  assign P53[3] = IN1[36]&IN2[17];
  assign P54[2] = IN1[36]&IN2[18];
  assign P55[1] = IN1[36]&IN2[19];
  assign P56[0] = IN1[36]&IN2[20];
  assign P37[20] = IN1[37]&IN2[0];
  assign P38[19] = IN1[37]&IN2[1];
  assign P39[18] = IN1[37]&IN2[2];
  assign P40[17] = IN1[37]&IN2[3];
  assign P41[16] = IN1[37]&IN2[4];
  assign P42[15] = IN1[37]&IN2[5];
  assign P43[14] = IN1[37]&IN2[6];
  assign P44[13] = IN1[37]&IN2[7];
  assign P45[12] = IN1[37]&IN2[8];
  assign P46[11] = IN1[37]&IN2[9];
  assign P47[10] = IN1[37]&IN2[10];
  assign P48[9] = IN1[37]&IN2[11];
  assign P49[8] = IN1[37]&IN2[12];
  assign P50[7] = IN1[37]&IN2[13];
  assign P51[6] = IN1[37]&IN2[14];
  assign P52[5] = IN1[37]&IN2[15];
  assign P53[4] = IN1[37]&IN2[16];
  assign P54[3] = IN1[37]&IN2[17];
  assign P55[2] = IN1[37]&IN2[18];
  assign P56[1] = IN1[37]&IN2[19];
  assign P57[0] = IN1[37]&IN2[20];
  assign P38[20] = IN1[38]&IN2[0];
  assign P39[19] = IN1[38]&IN2[1];
  assign P40[18] = IN1[38]&IN2[2];
  assign P41[17] = IN1[38]&IN2[3];
  assign P42[16] = IN1[38]&IN2[4];
  assign P43[15] = IN1[38]&IN2[5];
  assign P44[14] = IN1[38]&IN2[6];
  assign P45[13] = IN1[38]&IN2[7];
  assign P46[12] = IN1[38]&IN2[8];
  assign P47[11] = IN1[38]&IN2[9];
  assign P48[10] = IN1[38]&IN2[10];
  assign P49[9] = IN1[38]&IN2[11];
  assign P50[8] = IN1[38]&IN2[12];
  assign P51[7] = IN1[38]&IN2[13];
  assign P52[6] = IN1[38]&IN2[14];
  assign P53[5] = IN1[38]&IN2[15];
  assign P54[4] = IN1[38]&IN2[16];
  assign P55[3] = IN1[38]&IN2[17];
  assign P56[2] = IN1[38]&IN2[18];
  assign P57[1] = IN1[38]&IN2[19];
  assign P58[0] = IN1[38]&IN2[20];
  assign P39[20] = IN1[39]&IN2[0];
  assign P40[19] = IN1[39]&IN2[1];
  assign P41[18] = IN1[39]&IN2[2];
  assign P42[17] = IN1[39]&IN2[3];
  assign P43[16] = IN1[39]&IN2[4];
  assign P44[15] = IN1[39]&IN2[5];
  assign P45[14] = IN1[39]&IN2[6];
  assign P46[13] = IN1[39]&IN2[7];
  assign P47[12] = IN1[39]&IN2[8];
  assign P48[11] = IN1[39]&IN2[9];
  assign P49[10] = IN1[39]&IN2[10];
  assign P50[9] = IN1[39]&IN2[11];
  assign P51[8] = IN1[39]&IN2[12];
  assign P52[7] = IN1[39]&IN2[13];
  assign P53[6] = IN1[39]&IN2[14];
  assign P54[5] = IN1[39]&IN2[15];
  assign P55[4] = IN1[39]&IN2[16];
  assign P56[3] = IN1[39]&IN2[17];
  assign P57[2] = IN1[39]&IN2[18];
  assign P58[1] = IN1[39]&IN2[19];
  assign P59[0] = IN1[39]&IN2[20];
  assign P40[20] = IN1[40]&IN2[0];
  assign P41[19] = IN1[40]&IN2[1];
  assign P42[18] = IN1[40]&IN2[2];
  assign P43[17] = IN1[40]&IN2[3];
  assign P44[16] = IN1[40]&IN2[4];
  assign P45[15] = IN1[40]&IN2[5];
  assign P46[14] = IN1[40]&IN2[6];
  assign P47[13] = IN1[40]&IN2[7];
  assign P48[12] = IN1[40]&IN2[8];
  assign P49[11] = IN1[40]&IN2[9];
  assign P50[10] = IN1[40]&IN2[10];
  assign P51[9] = IN1[40]&IN2[11];
  assign P52[8] = IN1[40]&IN2[12];
  assign P53[7] = IN1[40]&IN2[13];
  assign P54[6] = IN1[40]&IN2[14];
  assign P55[5] = IN1[40]&IN2[15];
  assign P56[4] = IN1[40]&IN2[16];
  assign P57[3] = IN1[40]&IN2[17];
  assign P58[2] = IN1[40]&IN2[18];
  assign P59[1] = IN1[40]&IN2[19];
  assign P60[0] = IN1[40]&IN2[20];
  assign P41[20] = IN1[41]&IN2[0];
  assign P42[19] = IN1[41]&IN2[1];
  assign P43[18] = IN1[41]&IN2[2];
  assign P44[17] = IN1[41]&IN2[3];
  assign P45[16] = IN1[41]&IN2[4];
  assign P46[15] = IN1[41]&IN2[5];
  assign P47[14] = IN1[41]&IN2[6];
  assign P48[13] = IN1[41]&IN2[7];
  assign P49[12] = IN1[41]&IN2[8];
  assign P50[11] = IN1[41]&IN2[9];
  assign P51[10] = IN1[41]&IN2[10];
  assign P52[9] = IN1[41]&IN2[11];
  assign P53[8] = IN1[41]&IN2[12];
  assign P54[7] = IN1[41]&IN2[13];
  assign P55[6] = IN1[41]&IN2[14];
  assign P56[5] = IN1[41]&IN2[15];
  assign P57[4] = IN1[41]&IN2[16];
  assign P58[3] = IN1[41]&IN2[17];
  assign P59[2] = IN1[41]&IN2[18];
  assign P60[1] = IN1[41]&IN2[19];
  assign P61[0] = IN1[41]&IN2[20];
  assign P42[20] = IN1[42]&IN2[0];
  assign P43[19] = IN1[42]&IN2[1];
  assign P44[18] = IN1[42]&IN2[2];
  assign P45[17] = IN1[42]&IN2[3];
  assign P46[16] = IN1[42]&IN2[4];
  assign P47[15] = IN1[42]&IN2[5];
  assign P48[14] = IN1[42]&IN2[6];
  assign P49[13] = IN1[42]&IN2[7];
  assign P50[12] = IN1[42]&IN2[8];
  assign P51[11] = IN1[42]&IN2[9];
  assign P52[10] = IN1[42]&IN2[10];
  assign P53[9] = IN1[42]&IN2[11];
  assign P54[8] = IN1[42]&IN2[12];
  assign P55[7] = IN1[42]&IN2[13];
  assign P56[6] = IN1[42]&IN2[14];
  assign P57[5] = IN1[42]&IN2[15];
  assign P58[4] = IN1[42]&IN2[16];
  assign P59[3] = IN1[42]&IN2[17];
  assign P60[2] = IN1[42]&IN2[18];
  assign P61[1] = IN1[42]&IN2[19];
  assign P62[0] = IN1[42]&IN2[20];
  assign P43[20] = IN1[43]&IN2[0];
  assign P44[19] = IN1[43]&IN2[1];
  assign P45[18] = IN1[43]&IN2[2];
  assign P46[17] = IN1[43]&IN2[3];
  assign P47[16] = IN1[43]&IN2[4];
  assign P48[15] = IN1[43]&IN2[5];
  assign P49[14] = IN1[43]&IN2[6];
  assign P50[13] = IN1[43]&IN2[7];
  assign P51[12] = IN1[43]&IN2[8];
  assign P52[11] = IN1[43]&IN2[9];
  assign P53[10] = IN1[43]&IN2[10];
  assign P54[9] = IN1[43]&IN2[11];
  assign P55[8] = IN1[43]&IN2[12];
  assign P56[7] = IN1[43]&IN2[13];
  assign P57[6] = IN1[43]&IN2[14];
  assign P58[5] = IN1[43]&IN2[15];
  assign P59[4] = IN1[43]&IN2[16];
  assign P60[3] = IN1[43]&IN2[17];
  assign P61[2] = IN1[43]&IN2[18];
  assign P62[1] = IN1[43]&IN2[19];
  assign P63[0] = IN1[43]&IN2[20];
  assign P44[20] = IN1[44]&IN2[0];
  assign P45[19] = IN1[44]&IN2[1];
  assign P46[18] = IN1[44]&IN2[2];
  assign P47[17] = IN1[44]&IN2[3];
  assign P48[16] = IN1[44]&IN2[4];
  assign P49[15] = IN1[44]&IN2[5];
  assign P50[14] = IN1[44]&IN2[6];
  assign P51[13] = IN1[44]&IN2[7];
  assign P52[12] = IN1[44]&IN2[8];
  assign P53[11] = IN1[44]&IN2[9];
  assign P54[10] = IN1[44]&IN2[10];
  assign P55[9] = IN1[44]&IN2[11];
  assign P56[8] = IN1[44]&IN2[12];
  assign P57[7] = IN1[44]&IN2[13];
  assign P58[6] = IN1[44]&IN2[14];
  assign P59[5] = IN1[44]&IN2[15];
  assign P60[4] = IN1[44]&IN2[16];
  assign P61[3] = IN1[44]&IN2[17];
  assign P62[2] = IN1[44]&IN2[18];
  assign P63[1] = IN1[44]&IN2[19];
  assign P64[0] = IN1[44]&IN2[20];
  assign P45[20] = IN1[45]&IN2[0];
  assign P46[19] = IN1[45]&IN2[1];
  assign P47[18] = IN1[45]&IN2[2];
  assign P48[17] = IN1[45]&IN2[3];
  assign P49[16] = IN1[45]&IN2[4];
  assign P50[15] = IN1[45]&IN2[5];
  assign P51[14] = IN1[45]&IN2[6];
  assign P52[13] = IN1[45]&IN2[7];
  assign P53[12] = IN1[45]&IN2[8];
  assign P54[11] = IN1[45]&IN2[9];
  assign P55[10] = IN1[45]&IN2[10];
  assign P56[9] = IN1[45]&IN2[11];
  assign P57[8] = IN1[45]&IN2[12];
  assign P58[7] = IN1[45]&IN2[13];
  assign P59[6] = IN1[45]&IN2[14];
  assign P60[5] = IN1[45]&IN2[15];
  assign P61[4] = IN1[45]&IN2[16];
  assign P62[3] = IN1[45]&IN2[17];
  assign P63[2] = IN1[45]&IN2[18];
  assign P64[1] = IN1[45]&IN2[19];
  assign P65[0] = IN1[45]&IN2[20];
  assign P46[20] = IN1[46]&IN2[0];
  assign P47[19] = IN1[46]&IN2[1];
  assign P48[18] = IN1[46]&IN2[2];
  assign P49[17] = IN1[46]&IN2[3];
  assign P50[16] = IN1[46]&IN2[4];
  assign P51[15] = IN1[46]&IN2[5];
  assign P52[14] = IN1[46]&IN2[6];
  assign P53[13] = IN1[46]&IN2[7];
  assign P54[12] = IN1[46]&IN2[8];
  assign P55[11] = IN1[46]&IN2[9];
  assign P56[10] = IN1[46]&IN2[10];
  assign P57[9] = IN1[46]&IN2[11];
  assign P58[8] = IN1[46]&IN2[12];
  assign P59[7] = IN1[46]&IN2[13];
  assign P60[6] = IN1[46]&IN2[14];
  assign P61[5] = IN1[46]&IN2[15];
  assign P62[4] = IN1[46]&IN2[16];
  assign P63[3] = IN1[46]&IN2[17];
  assign P64[2] = IN1[46]&IN2[18];
  assign P65[1] = IN1[46]&IN2[19];
  assign P66[0] = IN1[46]&IN2[20];
  assign P47[20] = IN1[47]&IN2[0];
  assign P48[19] = IN1[47]&IN2[1];
  assign P49[18] = IN1[47]&IN2[2];
  assign P50[17] = IN1[47]&IN2[3];
  assign P51[16] = IN1[47]&IN2[4];
  assign P52[15] = IN1[47]&IN2[5];
  assign P53[14] = IN1[47]&IN2[6];
  assign P54[13] = IN1[47]&IN2[7];
  assign P55[12] = IN1[47]&IN2[8];
  assign P56[11] = IN1[47]&IN2[9];
  assign P57[10] = IN1[47]&IN2[10];
  assign P58[9] = IN1[47]&IN2[11];
  assign P59[8] = IN1[47]&IN2[12];
  assign P60[7] = IN1[47]&IN2[13];
  assign P61[6] = IN1[47]&IN2[14];
  assign P62[5] = IN1[47]&IN2[15];
  assign P63[4] = IN1[47]&IN2[16];
  assign P64[3] = IN1[47]&IN2[17];
  assign P65[2] = IN1[47]&IN2[18];
  assign P66[1] = IN1[47]&IN2[19];
  assign P67[0] = IN1[47]&IN2[20];
  assign P48[20] = IN1[48]&IN2[0];
  assign P49[19] = IN1[48]&IN2[1];
  assign P50[18] = IN1[48]&IN2[2];
  assign P51[17] = IN1[48]&IN2[3];
  assign P52[16] = IN1[48]&IN2[4];
  assign P53[15] = IN1[48]&IN2[5];
  assign P54[14] = IN1[48]&IN2[6];
  assign P55[13] = IN1[48]&IN2[7];
  assign P56[12] = IN1[48]&IN2[8];
  assign P57[11] = IN1[48]&IN2[9];
  assign P58[10] = IN1[48]&IN2[10];
  assign P59[9] = IN1[48]&IN2[11];
  assign P60[8] = IN1[48]&IN2[12];
  assign P61[7] = IN1[48]&IN2[13];
  assign P62[6] = IN1[48]&IN2[14];
  assign P63[5] = IN1[48]&IN2[15];
  assign P64[4] = IN1[48]&IN2[16];
  assign P65[3] = IN1[48]&IN2[17];
  assign P66[2] = IN1[48]&IN2[18];
  assign P67[1] = IN1[48]&IN2[19];
  assign P68[0] = IN1[48]&IN2[20];
  assign P49[20] = IN1[49]&IN2[0];
  assign P50[19] = IN1[49]&IN2[1];
  assign P51[18] = IN1[49]&IN2[2];
  assign P52[17] = IN1[49]&IN2[3];
  assign P53[16] = IN1[49]&IN2[4];
  assign P54[15] = IN1[49]&IN2[5];
  assign P55[14] = IN1[49]&IN2[6];
  assign P56[13] = IN1[49]&IN2[7];
  assign P57[12] = IN1[49]&IN2[8];
  assign P58[11] = IN1[49]&IN2[9];
  assign P59[10] = IN1[49]&IN2[10];
  assign P60[9] = IN1[49]&IN2[11];
  assign P61[8] = IN1[49]&IN2[12];
  assign P62[7] = IN1[49]&IN2[13];
  assign P63[6] = IN1[49]&IN2[14];
  assign P64[5] = IN1[49]&IN2[15];
  assign P65[4] = IN1[49]&IN2[16];
  assign P66[3] = IN1[49]&IN2[17];
  assign P67[2] = IN1[49]&IN2[18];
  assign P68[1] = IN1[49]&IN2[19];
  assign P69[0] = IN1[49]&IN2[20];
  assign P50[20] = IN1[50]&IN2[0];
  assign P51[19] = IN1[50]&IN2[1];
  assign P52[18] = IN1[50]&IN2[2];
  assign P53[17] = IN1[50]&IN2[3];
  assign P54[16] = IN1[50]&IN2[4];
  assign P55[15] = IN1[50]&IN2[5];
  assign P56[14] = IN1[50]&IN2[6];
  assign P57[13] = IN1[50]&IN2[7];
  assign P58[12] = IN1[50]&IN2[8];
  assign P59[11] = IN1[50]&IN2[9];
  assign P60[10] = IN1[50]&IN2[10];
  assign P61[9] = IN1[50]&IN2[11];
  assign P62[8] = IN1[50]&IN2[12];
  assign P63[7] = IN1[50]&IN2[13];
  assign P64[6] = IN1[50]&IN2[14];
  assign P65[5] = IN1[50]&IN2[15];
  assign P66[4] = IN1[50]&IN2[16];
  assign P67[3] = IN1[50]&IN2[17];
  assign P68[2] = IN1[50]&IN2[18];
  assign P69[1] = IN1[50]&IN2[19];
  assign P70[0] = IN1[50]&IN2[20];
  assign P51[20] = IN1[51]&IN2[0];
  assign P52[19] = IN1[51]&IN2[1];
  assign P53[18] = IN1[51]&IN2[2];
  assign P54[17] = IN1[51]&IN2[3];
  assign P55[16] = IN1[51]&IN2[4];
  assign P56[15] = IN1[51]&IN2[5];
  assign P57[14] = IN1[51]&IN2[6];
  assign P58[13] = IN1[51]&IN2[7];
  assign P59[12] = IN1[51]&IN2[8];
  assign P60[11] = IN1[51]&IN2[9];
  assign P61[10] = IN1[51]&IN2[10];
  assign P62[9] = IN1[51]&IN2[11];
  assign P63[8] = IN1[51]&IN2[12];
  assign P64[7] = IN1[51]&IN2[13];
  assign P65[6] = IN1[51]&IN2[14];
  assign P66[5] = IN1[51]&IN2[15];
  assign P67[4] = IN1[51]&IN2[16];
  assign P68[3] = IN1[51]&IN2[17];
  assign P69[2] = IN1[51]&IN2[18];
  assign P70[1] = IN1[51]&IN2[19];
  assign P71[0] = IN1[51]&IN2[20];
  assign P52[20] = IN1[52]&IN2[0];
  assign P53[19] = IN1[52]&IN2[1];
  assign P54[18] = IN1[52]&IN2[2];
  assign P55[17] = IN1[52]&IN2[3];
  assign P56[16] = IN1[52]&IN2[4];
  assign P57[15] = IN1[52]&IN2[5];
  assign P58[14] = IN1[52]&IN2[6];
  assign P59[13] = IN1[52]&IN2[7];
  assign P60[12] = IN1[52]&IN2[8];
  assign P61[11] = IN1[52]&IN2[9];
  assign P62[10] = IN1[52]&IN2[10];
  assign P63[9] = IN1[52]&IN2[11];
  assign P64[8] = IN1[52]&IN2[12];
  assign P65[7] = IN1[52]&IN2[13];
  assign P66[6] = IN1[52]&IN2[14];
  assign P67[5] = IN1[52]&IN2[15];
  assign P68[4] = IN1[52]&IN2[16];
  assign P69[3] = IN1[52]&IN2[17];
  assign P70[2] = IN1[52]&IN2[18];
  assign P71[1] = IN1[52]&IN2[19];
  assign P72[0] = IN1[52]&IN2[20];
  assign P53[20] = IN1[53]&IN2[0];
  assign P54[19] = IN1[53]&IN2[1];
  assign P55[18] = IN1[53]&IN2[2];
  assign P56[17] = IN1[53]&IN2[3];
  assign P57[16] = IN1[53]&IN2[4];
  assign P58[15] = IN1[53]&IN2[5];
  assign P59[14] = IN1[53]&IN2[6];
  assign P60[13] = IN1[53]&IN2[7];
  assign P61[12] = IN1[53]&IN2[8];
  assign P62[11] = IN1[53]&IN2[9];
  assign P63[10] = IN1[53]&IN2[10];
  assign P64[9] = IN1[53]&IN2[11];
  assign P65[8] = IN1[53]&IN2[12];
  assign P66[7] = IN1[53]&IN2[13];
  assign P67[6] = IN1[53]&IN2[14];
  assign P68[5] = IN1[53]&IN2[15];
  assign P69[4] = IN1[53]&IN2[16];
  assign P70[3] = IN1[53]&IN2[17];
  assign P71[2] = IN1[53]&IN2[18];
  assign P72[1] = IN1[53]&IN2[19];
  assign P73[0] = IN1[53]&IN2[20];
  assign P54[20] = IN1[54]&IN2[0];
  assign P55[19] = IN1[54]&IN2[1];
  assign P56[18] = IN1[54]&IN2[2];
  assign P57[17] = IN1[54]&IN2[3];
  assign P58[16] = IN1[54]&IN2[4];
  assign P59[15] = IN1[54]&IN2[5];
  assign P60[14] = IN1[54]&IN2[6];
  assign P61[13] = IN1[54]&IN2[7];
  assign P62[12] = IN1[54]&IN2[8];
  assign P63[11] = IN1[54]&IN2[9];
  assign P64[10] = IN1[54]&IN2[10];
  assign P65[9] = IN1[54]&IN2[11];
  assign P66[8] = IN1[54]&IN2[12];
  assign P67[7] = IN1[54]&IN2[13];
  assign P68[6] = IN1[54]&IN2[14];
  assign P69[5] = IN1[54]&IN2[15];
  assign P70[4] = IN1[54]&IN2[16];
  assign P71[3] = IN1[54]&IN2[17];
  assign P72[2] = IN1[54]&IN2[18];
  assign P73[1] = IN1[54]&IN2[19];
  assign P74[0] = IN1[54]&IN2[20];
  assign P55[20] = IN1[55]&IN2[0];
  assign P56[19] = IN1[55]&IN2[1];
  assign P57[18] = IN1[55]&IN2[2];
  assign P58[17] = IN1[55]&IN2[3];
  assign P59[16] = IN1[55]&IN2[4];
  assign P60[15] = IN1[55]&IN2[5];
  assign P61[14] = IN1[55]&IN2[6];
  assign P62[13] = IN1[55]&IN2[7];
  assign P63[12] = IN1[55]&IN2[8];
  assign P64[11] = IN1[55]&IN2[9];
  assign P65[10] = IN1[55]&IN2[10];
  assign P66[9] = IN1[55]&IN2[11];
  assign P67[8] = IN1[55]&IN2[12];
  assign P68[7] = IN1[55]&IN2[13];
  assign P69[6] = IN1[55]&IN2[14];
  assign P70[5] = IN1[55]&IN2[15];
  assign P71[4] = IN1[55]&IN2[16];
  assign P72[3] = IN1[55]&IN2[17];
  assign P73[2] = IN1[55]&IN2[18];
  assign P74[1] = IN1[55]&IN2[19];
  assign P75[0] = IN1[55]&IN2[20];
  assign P56[20] = IN1[56]&IN2[0];
  assign P57[19] = IN1[56]&IN2[1];
  assign P58[18] = IN1[56]&IN2[2];
  assign P59[17] = IN1[56]&IN2[3];
  assign P60[16] = IN1[56]&IN2[4];
  assign P61[15] = IN1[56]&IN2[5];
  assign P62[14] = IN1[56]&IN2[6];
  assign P63[13] = IN1[56]&IN2[7];
  assign P64[12] = IN1[56]&IN2[8];
  assign P65[11] = IN1[56]&IN2[9];
  assign P66[10] = IN1[56]&IN2[10];
  assign P67[9] = IN1[56]&IN2[11];
  assign P68[8] = IN1[56]&IN2[12];
  assign P69[7] = IN1[56]&IN2[13];
  assign P70[6] = IN1[56]&IN2[14];
  assign P71[5] = IN1[56]&IN2[15];
  assign P72[4] = IN1[56]&IN2[16];
  assign P73[3] = IN1[56]&IN2[17];
  assign P74[2] = IN1[56]&IN2[18];
  assign P75[1] = IN1[56]&IN2[19];
  assign P76[0] = IN1[56]&IN2[20];
  assign P57[20] = IN1[57]&IN2[0];
  assign P58[19] = IN1[57]&IN2[1];
  assign P59[18] = IN1[57]&IN2[2];
  assign P60[17] = IN1[57]&IN2[3];
  assign P61[16] = IN1[57]&IN2[4];
  assign P62[15] = IN1[57]&IN2[5];
  assign P63[14] = IN1[57]&IN2[6];
  assign P64[13] = IN1[57]&IN2[7];
  assign P65[12] = IN1[57]&IN2[8];
  assign P66[11] = IN1[57]&IN2[9];
  assign P67[10] = IN1[57]&IN2[10];
  assign P68[9] = IN1[57]&IN2[11];
  assign P69[8] = IN1[57]&IN2[12];
  assign P70[7] = IN1[57]&IN2[13];
  assign P71[6] = IN1[57]&IN2[14];
  assign P72[5] = IN1[57]&IN2[15];
  assign P73[4] = IN1[57]&IN2[16];
  assign P74[3] = IN1[57]&IN2[17];
  assign P75[2] = IN1[57]&IN2[18];
  assign P76[1] = IN1[57]&IN2[19];
  assign P77[0] = IN1[57]&IN2[20];
  assign P58[20] = IN1[58]&IN2[0];
  assign P59[19] = IN1[58]&IN2[1];
  assign P60[18] = IN1[58]&IN2[2];
  assign P61[17] = IN1[58]&IN2[3];
  assign P62[16] = IN1[58]&IN2[4];
  assign P63[15] = IN1[58]&IN2[5];
  assign P64[14] = IN1[58]&IN2[6];
  assign P65[13] = IN1[58]&IN2[7];
  assign P66[12] = IN1[58]&IN2[8];
  assign P67[11] = IN1[58]&IN2[9];
  assign P68[10] = IN1[58]&IN2[10];
  assign P69[9] = IN1[58]&IN2[11];
  assign P70[8] = IN1[58]&IN2[12];
  assign P71[7] = IN1[58]&IN2[13];
  assign P72[6] = IN1[58]&IN2[14];
  assign P73[5] = IN1[58]&IN2[15];
  assign P74[4] = IN1[58]&IN2[16];
  assign P75[3] = IN1[58]&IN2[17];
  assign P76[2] = IN1[58]&IN2[18];
  assign P77[1] = IN1[58]&IN2[19];
  assign P78[0] = IN1[58]&IN2[20];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [20:0] IN21;
  input [20:0] IN22;
  input [20:0] IN23;
  input [20:0] IN24;
  input [20:0] IN25;
  input [20:0] IN26;
  input [20:0] IN27;
  input [20:0] IN28;
  input [20:0] IN29;
  input [20:0] IN30;
  input [20:0] IN31;
  input [20:0] IN32;
  input [20:0] IN33;
  input [20:0] IN34;
  input [20:0] IN35;
  input [20:0] IN36;
  input [20:0] IN37;
  input [20:0] IN38;
  input [20:0] IN39;
  input [20:0] IN40;
  input [20:0] IN41;
  input [20:0] IN42;
  input [20:0] IN43;
  input [20:0] IN44;
  input [20:0] IN45;
  input [20:0] IN46;
  input [20:0] IN47;
  input [20:0] IN48;
  input [20:0] IN49;
  input [20:0] IN50;
  input [20:0] IN51;
  input [20:0] IN52;
  input [20:0] IN53;
  input [20:0] IN54;
  input [20:0] IN55;
  input [20:0] IN56;
  input [20:0] IN57;
  input [20:0] IN58;
  input [19:0] IN59;
  input [18:0] IN60;
  input [17:0] IN61;
  input [16:0] IN62;
  input [15:0] IN63;
  input [14:0] IN64;
  input [13:0] IN65;
  input [12:0] IN66;
  input [11:0] IN67;
  input [10:0] IN68;
  input [9:0] IN69;
  input [8:0] IN70;
  input [7:0] IN71;
  input [6:0] IN72;
  input [5:0] IN73;
  input [4:0] IN74;
  input [3:0] IN75;
  input [2:0] IN76;
  input [1:0] IN77;
  input [0:0] IN78;
  output [78:0] Out1;
  output [19:0] Out2;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1932;
  wire w1933;
  wire w1934;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1958;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1984;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2010;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2036;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2050;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2062;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2088;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2114;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2140;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2166;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2192;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2374;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2454;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2534;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2585;
  wire w2586;
  wire w2587;
  wire w2588;
  wire w2589;
  wire w2590;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2614;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2638;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2680;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2685;
  wire w2686;
  wire w2687;
  wire w2688;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2694;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2708;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2738;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2770;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2774;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2785;
  wire w2786;
  wire w2787;
  wire w2788;
  wire w2789;
  wire w2790;
  wire w2791;
  wire w2792;
  wire w2793;
  wire w2794;
  wire w2795;
  wire w2796;
  wire w2797;
  wire w2798;
  wire w2799;
  wire w2800;
  wire w2801;
  wire w2802;
  wire w2803;
  wire w2804;
  wire w2805;
  wire w2806;
  wire w2807;
  wire w2808;
  wire w2809;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2854;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2860;
  wire w2861;
  wire w2862;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2885;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2896;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2913;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2934;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2950;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2985;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2990;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3014;
  wire w3015;
  wire w3016;
  wire w3017;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3040;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3084;
  wire w3085;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3094;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3121;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3130;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3174;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3225;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3254;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3262;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3272;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3285;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3328;
  wire w3329;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3334;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3362;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3366;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3385;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3414;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3433;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3444;
  wire w3446;
  wire w3448;
  wire w3450;
  wire w3452;
  wire w3454;
  wire w3456;
  wire w3458;
  wire w3460;
  wire w3462;
  wire w3464;
  wire w3466;
  wire w3468;
  wire w3470;
  wire w3472;
  wire w3474;
  wire w3476;
  wire w3478;
  wire w3480;
  wire w3482;
  wire w3484;
  wire w3486;
  wire w3488;
  wire w3490;
  wire w3492;
  wire w3494;
  wire w3496;
  wire w3498;
  wire w3500;
  wire w3502;
  wire w3504;
  wire w3506;
  wire w3508;
  wire w3510;
  wire w3512;
  wire w3514;
  wire w3516;
  wire w3518;
  wire w3520;
  wire w3522;
  wire w3524;
  wire w3526;
  wire w3528;
  wire w3530;
  wire w3532;
  wire w3534;
  wire w3536;
  wire w3538;
  wire w3540;
  wire w3542;
  wire w3544;
  wire w3546;
  wire w3548;
  wire w3550;
  wire w3552;
  wire w3554;
  wire w3556;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w1240);
  FullAdder U1 (w1240, IN2[0], IN2[1], w1241, w1242);
  FullAdder U2 (w1242, IN3[0], IN3[1], w1243, w1244);
  FullAdder U3 (w1244, IN4[0], IN4[1], w1245, w1246);
  FullAdder U4 (w1246, IN5[0], IN5[1], w1247, w1248);
  FullAdder U5 (w1248, IN6[0], IN6[1], w1249, w1250);
  FullAdder U6 (w1250, IN7[0], IN7[1], w1251, w1252);
  FullAdder U7 (w1252, IN8[0], IN8[1], w1253, w1254);
  FullAdder U8 (w1254, IN9[0], IN9[1], w1255, w1256);
  FullAdder U9 (w1256, IN10[0], IN10[1], w1257, w1258);
  FullAdder U10 (w1258, IN11[0], IN11[1], w1259, w1260);
  FullAdder U11 (w1260, IN12[0], IN12[1], w1261, w1262);
  FullAdder U12 (w1262, IN13[0], IN13[1], w1263, w1264);
  FullAdder U13 (w1264, IN14[0], IN14[1], w1265, w1266);
  FullAdder U14 (w1266, IN15[0], IN15[1], w1267, w1268);
  FullAdder U15 (w1268, IN16[0], IN16[1], w1269, w1270);
  FullAdder U16 (w1270, IN17[0], IN17[1], w1271, w1272);
  FullAdder U17 (w1272, IN18[0], IN18[1], w1273, w1274);
  FullAdder U18 (w1274, IN19[0], IN19[1], w1275, w1276);
  FullAdder U19 (w1276, IN20[0], IN20[1], w1277, w1278);
  FullAdder U20 (w1278, IN21[0], IN21[1], w1279, w1280);
  FullAdder U21 (w1280, IN22[0], IN22[1], w1281, w1282);
  FullAdder U22 (w1282, IN23[0], IN23[1], w1283, w1284);
  FullAdder U23 (w1284, IN24[0], IN24[1], w1285, w1286);
  FullAdder U24 (w1286, IN25[0], IN25[1], w1287, w1288);
  FullAdder U25 (w1288, IN26[0], IN26[1], w1289, w1290);
  FullAdder U26 (w1290, IN27[0], IN27[1], w1291, w1292);
  FullAdder U27 (w1292, IN28[0], IN28[1], w1293, w1294);
  FullAdder U28 (w1294, IN29[0], IN29[1], w1295, w1296);
  FullAdder U29 (w1296, IN30[0], IN30[1], w1297, w1298);
  FullAdder U30 (w1298, IN31[0], IN31[1], w1299, w1300);
  FullAdder U31 (w1300, IN32[0], IN32[1], w1301, w1302);
  FullAdder U32 (w1302, IN33[0], IN33[1], w1303, w1304);
  FullAdder U33 (w1304, IN34[0], IN34[1], w1305, w1306);
  FullAdder U34 (w1306, IN35[0], IN35[1], w1307, w1308);
  FullAdder U35 (w1308, IN36[0], IN36[1], w1309, w1310);
  FullAdder U36 (w1310, IN37[0], IN37[1], w1311, w1312);
  FullAdder U37 (w1312, IN38[0], IN38[1], w1313, w1314);
  FullAdder U38 (w1314, IN39[0], IN39[1], w1315, w1316);
  FullAdder U39 (w1316, IN40[0], IN40[1], w1317, w1318);
  FullAdder U40 (w1318, IN41[0], IN41[1], w1319, w1320);
  FullAdder U41 (w1320, IN42[0], IN42[1], w1321, w1322);
  FullAdder U42 (w1322, IN43[0], IN43[1], w1323, w1324);
  FullAdder U43 (w1324, IN44[0], IN44[1], w1325, w1326);
  FullAdder U44 (w1326, IN45[0], IN45[1], w1327, w1328);
  FullAdder U45 (w1328, IN46[0], IN46[1], w1329, w1330);
  FullAdder U46 (w1330, IN47[0], IN47[1], w1331, w1332);
  FullAdder U47 (w1332, IN48[0], IN48[1], w1333, w1334);
  FullAdder U48 (w1334, IN49[0], IN49[1], w1335, w1336);
  FullAdder U49 (w1336, IN50[0], IN50[1], w1337, w1338);
  FullAdder U50 (w1338, IN51[0], IN51[1], w1339, w1340);
  FullAdder U51 (w1340, IN52[0], IN52[1], w1341, w1342);
  FullAdder U52 (w1342, IN53[0], IN53[1], w1343, w1344);
  FullAdder U53 (w1344, IN54[0], IN54[1], w1345, w1346);
  FullAdder U54 (w1346, IN55[0], IN55[1], w1347, w1348);
  FullAdder U55 (w1348, IN56[0], IN56[1], w1349, w1350);
  FullAdder U56 (w1350, IN57[0], IN57[1], w1351, w1352);
  FullAdder U57 (w1352, IN58[0], IN58[1], w1353, w1354);
  HalfAdder U58 (w1241, IN2[2], Out1[2], w1356);
  FullAdder U59 (w1356, w1243, IN3[2], w1357, w1358);
  FullAdder U60 (w1358, w1245, IN4[2], w1359, w1360);
  FullAdder U61 (w1360, w1247, IN5[2], w1361, w1362);
  FullAdder U62 (w1362, w1249, IN6[2], w1363, w1364);
  FullAdder U63 (w1364, w1251, IN7[2], w1365, w1366);
  FullAdder U64 (w1366, w1253, IN8[2], w1367, w1368);
  FullAdder U65 (w1368, w1255, IN9[2], w1369, w1370);
  FullAdder U66 (w1370, w1257, IN10[2], w1371, w1372);
  FullAdder U67 (w1372, w1259, IN11[2], w1373, w1374);
  FullAdder U68 (w1374, w1261, IN12[2], w1375, w1376);
  FullAdder U69 (w1376, w1263, IN13[2], w1377, w1378);
  FullAdder U70 (w1378, w1265, IN14[2], w1379, w1380);
  FullAdder U71 (w1380, w1267, IN15[2], w1381, w1382);
  FullAdder U72 (w1382, w1269, IN16[2], w1383, w1384);
  FullAdder U73 (w1384, w1271, IN17[2], w1385, w1386);
  FullAdder U74 (w1386, w1273, IN18[2], w1387, w1388);
  FullAdder U75 (w1388, w1275, IN19[2], w1389, w1390);
  FullAdder U76 (w1390, w1277, IN20[2], w1391, w1392);
  FullAdder U77 (w1392, w1279, IN21[2], w1393, w1394);
  FullAdder U78 (w1394, w1281, IN22[2], w1395, w1396);
  FullAdder U79 (w1396, w1283, IN23[2], w1397, w1398);
  FullAdder U80 (w1398, w1285, IN24[2], w1399, w1400);
  FullAdder U81 (w1400, w1287, IN25[2], w1401, w1402);
  FullAdder U82 (w1402, w1289, IN26[2], w1403, w1404);
  FullAdder U83 (w1404, w1291, IN27[2], w1405, w1406);
  FullAdder U84 (w1406, w1293, IN28[2], w1407, w1408);
  FullAdder U85 (w1408, w1295, IN29[2], w1409, w1410);
  FullAdder U86 (w1410, w1297, IN30[2], w1411, w1412);
  FullAdder U87 (w1412, w1299, IN31[2], w1413, w1414);
  FullAdder U88 (w1414, w1301, IN32[2], w1415, w1416);
  FullAdder U89 (w1416, w1303, IN33[2], w1417, w1418);
  FullAdder U90 (w1418, w1305, IN34[2], w1419, w1420);
  FullAdder U91 (w1420, w1307, IN35[2], w1421, w1422);
  FullAdder U92 (w1422, w1309, IN36[2], w1423, w1424);
  FullAdder U93 (w1424, w1311, IN37[2], w1425, w1426);
  FullAdder U94 (w1426, w1313, IN38[2], w1427, w1428);
  FullAdder U95 (w1428, w1315, IN39[2], w1429, w1430);
  FullAdder U96 (w1430, w1317, IN40[2], w1431, w1432);
  FullAdder U97 (w1432, w1319, IN41[2], w1433, w1434);
  FullAdder U98 (w1434, w1321, IN42[2], w1435, w1436);
  FullAdder U99 (w1436, w1323, IN43[2], w1437, w1438);
  FullAdder U100 (w1438, w1325, IN44[2], w1439, w1440);
  FullAdder U101 (w1440, w1327, IN45[2], w1441, w1442);
  FullAdder U102 (w1442, w1329, IN46[2], w1443, w1444);
  FullAdder U103 (w1444, w1331, IN47[2], w1445, w1446);
  FullAdder U104 (w1446, w1333, IN48[2], w1447, w1448);
  FullAdder U105 (w1448, w1335, IN49[2], w1449, w1450);
  FullAdder U106 (w1450, w1337, IN50[2], w1451, w1452);
  FullAdder U107 (w1452, w1339, IN51[2], w1453, w1454);
  FullAdder U108 (w1454, w1341, IN52[2], w1455, w1456);
  FullAdder U109 (w1456, w1343, IN53[2], w1457, w1458);
  FullAdder U110 (w1458, w1345, IN54[2], w1459, w1460);
  FullAdder U111 (w1460, w1347, IN55[2], w1461, w1462);
  FullAdder U112 (w1462, w1349, IN56[2], w1463, w1464);
  FullAdder U113 (w1464, w1351, IN57[2], w1465, w1466);
  FullAdder U114 (w1466, w1353, IN58[2], w1467, w1468);
  FullAdder U115 (w1468, w1354, IN59[0], w1469, w1470);
  HalfAdder U116 (w1357, IN3[3], Out1[3], w1472);
  FullAdder U117 (w1472, w1359, IN4[3], w1473, w1474);
  FullAdder U118 (w1474, w1361, IN5[3], w1475, w1476);
  FullAdder U119 (w1476, w1363, IN6[3], w1477, w1478);
  FullAdder U120 (w1478, w1365, IN7[3], w1479, w1480);
  FullAdder U121 (w1480, w1367, IN8[3], w1481, w1482);
  FullAdder U122 (w1482, w1369, IN9[3], w1483, w1484);
  FullAdder U123 (w1484, w1371, IN10[3], w1485, w1486);
  FullAdder U124 (w1486, w1373, IN11[3], w1487, w1488);
  FullAdder U125 (w1488, w1375, IN12[3], w1489, w1490);
  FullAdder U126 (w1490, w1377, IN13[3], w1491, w1492);
  FullAdder U127 (w1492, w1379, IN14[3], w1493, w1494);
  FullAdder U128 (w1494, w1381, IN15[3], w1495, w1496);
  FullAdder U129 (w1496, w1383, IN16[3], w1497, w1498);
  FullAdder U130 (w1498, w1385, IN17[3], w1499, w1500);
  FullAdder U131 (w1500, w1387, IN18[3], w1501, w1502);
  FullAdder U132 (w1502, w1389, IN19[3], w1503, w1504);
  FullAdder U133 (w1504, w1391, IN20[3], w1505, w1506);
  FullAdder U134 (w1506, w1393, IN21[3], w1507, w1508);
  FullAdder U135 (w1508, w1395, IN22[3], w1509, w1510);
  FullAdder U136 (w1510, w1397, IN23[3], w1511, w1512);
  FullAdder U137 (w1512, w1399, IN24[3], w1513, w1514);
  FullAdder U138 (w1514, w1401, IN25[3], w1515, w1516);
  FullAdder U139 (w1516, w1403, IN26[3], w1517, w1518);
  FullAdder U140 (w1518, w1405, IN27[3], w1519, w1520);
  FullAdder U141 (w1520, w1407, IN28[3], w1521, w1522);
  FullAdder U142 (w1522, w1409, IN29[3], w1523, w1524);
  FullAdder U143 (w1524, w1411, IN30[3], w1525, w1526);
  FullAdder U144 (w1526, w1413, IN31[3], w1527, w1528);
  FullAdder U145 (w1528, w1415, IN32[3], w1529, w1530);
  FullAdder U146 (w1530, w1417, IN33[3], w1531, w1532);
  FullAdder U147 (w1532, w1419, IN34[3], w1533, w1534);
  FullAdder U148 (w1534, w1421, IN35[3], w1535, w1536);
  FullAdder U149 (w1536, w1423, IN36[3], w1537, w1538);
  FullAdder U150 (w1538, w1425, IN37[3], w1539, w1540);
  FullAdder U151 (w1540, w1427, IN38[3], w1541, w1542);
  FullAdder U152 (w1542, w1429, IN39[3], w1543, w1544);
  FullAdder U153 (w1544, w1431, IN40[3], w1545, w1546);
  FullAdder U154 (w1546, w1433, IN41[3], w1547, w1548);
  FullAdder U155 (w1548, w1435, IN42[3], w1549, w1550);
  FullAdder U156 (w1550, w1437, IN43[3], w1551, w1552);
  FullAdder U157 (w1552, w1439, IN44[3], w1553, w1554);
  FullAdder U158 (w1554, w1441, IN45[3], w1555, w1556);
  FullAdder U159 (w1556, w1443, IN46[3], w1557, w1558);
  FullAdder U160 (w1558, w1445, IN47[3], w1559, w1560);
  FullAdder U161 (w1560, w1447, IN48[3], w1561, w1562);
  FullAdder U162 (w1562, w1449, IN49[3], w1563, w1564);
  FullAdder U163 (w1564, w1451, IN50[3], w1565, w1566);
  FullAdder U164 (w1566, w1453, IN51[3], w1567, w1568);
  FullAdder U165 (w1568, w1455, IN52[3], w1569, w1570);
  FullAdder U166 (w1570, w1457, IN53[3], w1571, w1572);
  FullAdder U167 (w1572, w1459, IN54[3], w1573, w1574);
  FullAdder U168 (w1574, w1461, IN55[3], w1575, w1576);
  FullAdder U169 (w1576, w1463, IN56[3], w1577, w1578);
  FullAdder U170 (w1578, w1465, IN57[3], w1579, w1580);
  FullAdder U171 (w1580, w1467, IN58[3], w1581, w1582);
  FullAdder U172 (w1582, w1469, IN59[1], w1583, w1584);
  FullAdder U173 (w1584, w1470, IN60[0], w1585, w1586);
  HalfAdder U174 (w1473, IN4[4], Out1[4], w1588);
  FullAdder U175 (w1588, w1475, IN5[4], w1589, w1590);
  FullAdder U176 (w1590, w1477, IN6[4], w1591, w1592);
  FullAdder U177 (w1592, w1479, IN7[4], w1593, w1594);
  FullAdder U178 (w1594, w1481, IN8[4], w1595, w1596);
  FullAdder U179 (w1596, w1483, IN9[4], w1597, w1598);
  FullAdder U180 (w1598, w1485, IN10[4], w1599, w1600);
  FullAdder U181 (w1600, w1487, IN11[4], w1601, w1602);
  FullAdder U182 (w1602, w1489, IN12[4], w1603, w1604);
  FullAdder U183 (w1604, w1491, IN13[4], w1605, w1606);
  FullAdder U184 (w1606, w1493, IN14[4], w1607, w1608);
  FullAdder U185 (w1608, w1495, IN15[4], w1609, w1610);
  FullAdder U186 (w1610, w1497, IN16[4], w1611, w1612);
  FullAdder U187 (w1612, w1499, IN17[4], w1613, w1614);
  FullAdder U188 (w1614, w1501, IN18[4], w1615, w1616);
  FullAdder U189 (w1616, w1503, IN19[4], w1617, w1618);
  FullAdder U190 (w1618, w1505, IN20[4], w1619, w1620);
  FullAdder U191 (w1620, w1507, IN21[4], w1621, w1622);
  FullAdder U192 (w1622, w1509, IN22[4], w1623, w1624);
  FullAdder U193 (w1624, w1511, IN23[4], w1625, w1626);
  FullAdder U194 (w1626, w1513, IN24[4], w1627, w1628);
  FullAdder U195 (w1628, w1515, IN25[4], w1629, w1630);
  FullAdder U196 (w1630, w1517, IN26[4], w1631, w1632);
  FullAdder U197 (w1632, w1519, IN27[4], w1633, w1634);
  FullAdder U198 (w1634, w1521, IN28[4], w1635, w1636);
  FullAdder U199 (w1636, w1523, IN29[4], w1637, w1638);
  FullAdder U200 (w1638, w1525, IN30[4], w1639, w1640);
  FullAdder U201 (w1640, w1527, IN31[4], w1641, w1642);
  FullAdder U202 (w1642, w1529, IN32[4], w1643, w1644);
  FullAdder U203 (w1644, w1531, IN33[4], w1645, w1646);
  FullAdder U204 (w1646, w1533, IN34[4], w1647, w1648);
  FullAdder U205 (w1648, w1535, IN35[4], w1649, w1650);
  FullAdder U206 (w1650, w1537, IN36[4], w1651, w1652);
  FullAdder U207 (w1652, w1539, IN37[4], w1653, w1654);
  FullAdder U208 (w1654, w1541, IN38[4], w1655, w1656);
  FullAdder U209 (w1656, w1543, IN39[4], w1657, w1658);
  FullAdder U210 (w1658, w1545, IN40[4], w1659, w1660);
  FullAdder U211 (w1660, w1547, IN41[4], w1661, w1662);
  FullAdder U212 (w1662, w1549, IN42[4], w1663, w1664);
  FullAdder U213 (w1664, w1551, IN43[4], w1665, w1666);
  FullAdder U214 (w1666, w1553, IN44[4], w1667, w1668);
  FullAdder U215 (w1668, w1555, IN45[4], w1669, w1670);
  FullAdder U216 (w1670, w1557, IN46[4], w1671, w1672);
  FullAdder U217 (w1672, w1559, IN47[4], w1673, w1674);
  FullAdder U218 (w1674, w1561, IN48[4], w1675, w1676);
  FullAdder U219 (w1676, w1563, IN49[4], w1677, w1678);
  FullAdder U220 (w1678, w1565, IN50[4], w1679, w1680);
  FullAdder U221 (w1680, w1567, IN51[4], w1681, w1682);
  FullAdder U222 (w1682, w1569, IN52[4], w1683, w1684);
  FullAdder U223 (w1684, w1571, IN53[4], w1685, w1686);
  FullAdder U224 (w1686, w1573, IN54[4], w1687, w1688);
  FullAdder U225 (w1688, w1575, IN55[4], w1689, w1690);
  FullAdder U226 (w1690, w1577, IN56[4], w1691, w1692);
  FullAdder U227 (w1692, w1579, IN57[4], w1693, w1694);
  FullAdder U228 (w1694, w1581, IN58[4], w1695, w1696);
  FullAdder U229 (w1696, w1583, IN59[2], w1697, w1698);
  FullAdder U230 (w1698, w1585, IN60[1], w1699, w1700);
  FullAdder U231 (w1700, w1586, IN61[0], w1701, w1702);
  HalfAdder U232 (w1589, IN5[5], Out1[5], w1704);
  FullAdder U233 (w1704, w1591, IN6[5], w1705, w1706);
  FullAdder U234 (w1706, w1593, IN7[5], w1707, w1708);
  FullAdder U235 (w1708, w1595, IN8[5], w1709, w1710);
  FullAdder U236 (w1710, w1597, IN9[5], w1711, w1712);
  FullAdder U237 (w1712, w1599, IN10[5], w1713, w1714);
  FullAdder U238 (w1714, w1601, IN11[5], w1715, w1716);
  FullAdder U239 (w1716, w1603, IN12[5], w1717, w1718);
  FullAdder U240 (w1718, w1605, IN13[5], w1719, w1720);
  FullAdder U241 (w1720, w1607, IN14[5], w1721, w1722);
  FullAdder U242 (w1722, w1609, IN15[5], w1723, w1724);
  FullAdder U243 (w1724, w1611, IN16[5], w1725, w1726);
  FullAdder U244 (w1726, w1613, IN17[5], w1727, w1728);
  FullAdder U245 (w1728, w1615, IN18[5], w1729, w1730);
  FullAdder U246 (w1730, w1617, IN19[5], w1731, w1732);
  FullAdder U247 (w1732, w1619, IN20[5], w1733, w1734);
  FullAdder U248 (w1734, w1621, IN21[5], w1735, w1736);
  FullAdder U249 (w1736, w1623, IN22[5], w1737, w1738);
  FullAdder U250 (w1738, w1625, IN23[5], w1739, w1740);
  FullAdder U251 (w1740, w1627, IN24[5], w1741, w1742);
  FullAdder U252 (w1742, w1629, IN25[5], w1743, w1744);
  FullAdder U253 (w1744, w1631, IN26[5], w1745, w1746);
  FullAdder U254 (w1746, w1633, IN27[5], w1747, w1748);
  FullAdder U255 (w1748, w1635, IN28[5], w1749, w1750);
  FullAdder U256 (w1750, w1637, IN29[5], w1751, w1752);
  FullAdder U257 (w1752, w1639, IN30[5], w1753, w1754);
  FullAdder U258 (w1754, w1641, IN31[5], w1755, w1756);
  FullAdder U259 (w1756, w1643, IN32[5], w1757, w1758);
  FullAdder U260 (w1758, w1645, IN33[5], w1759, w1760);
  FullAdder U261 (w1760, w1647, IN34[5], w1761, w1762);
  FullAdder U262 (w1762, w1649, IN35[5], w1763, w1764);
  FullAdder U263 (w1764, w1651, IN36[5], w1765, w1766);
  FullAdder U264 (w1766, w1653, IN37[5], w1767, w1768);
  FullAdder U265 (w1768, w1655, IN38[5], w1769, w1770);
  FullAdder U266 (w1770, w1657, IN39[5], w1771, w1772);
  FullAdder U267 (w1772, w1659, IN40[5], w1773, w1774);
  FullAdder U268 (w1774, w1661, IN41[5], w1775, w1776);
  FullAdder U269 (w1776, w1663, IN42[5], w1777, w1778);
  FullAdder U270 (w1778, w1665, IN43[5], w1779, w1780);
  FullAdder U271 (w1780, w1667, IN44[5], w1781, w1782);
  FullAdder U272 (w1782, w1669, IN45[5], w1783, w1784);
  FullAdder U273 (w1784, w1671, IN46[5], w1785, w1786);
  FullAdder U274 (w1786, w1673, IN47[5], w1787, w1788);
  FullAdder U275 (w1788, w1675, IN48[5], w1789, w1790);
  FullAdder U276 (w1790, w1677, IN49[5], w1791, w1792);
  FullAdder U277 (w1792, w1679, IN50[5], w1793, w1794);
  FullAdder U278 (w1794, w1681, IN51[5], w1795, w1796);
  FullAdder U279 (w1796, w1683, IN52[5], w1797, w1798);
  FullAdder U280 (w1798, w1685, IN53[5], w1799, w1800);
  FullAdder U281 (w1800, w1687, IN54[5], w1801, w1802);
  FullAdder U282 (w1802, w1689, IN55[5], w1803, w1804);
  FullAdder U283 (w1804, w1691, IN56[5], w1805, w1806);
  FullAdder U284 (w1806, w1693, IN57[5], w1807, w1808);
  FullAdder U285 (w1808, w1695, IN58[5], w1809, w1810);
  FullAdder U286 (w1810, w1697, IN59[3], w1811, w1812);
  FullAdder U287 (w1812, w1699, IN60[2], w1813, w1814);
  FullAdder U288 (w1814, w1701, IN61[1], w1815, w1816);
  FullAdder U289 (w1816, w1702, IN62[0], w1817, w1818);
  HalfAdder U290 (w1705, IN6[6], Out1[6], w1820);
  FullAdder U291 (w1820, w1707, IN7[6], w1821, w1822);
  FullAdder U292 (w1822, w1709, IN8[6], w1823, w1824);
  FullAdder U293 (w1824, w1711, IN9[6], w1825, w1826);
  FullAdder U294 (w1826, w1713, IN10[6], w1827, w1828);
  FullAdder U295 (w1828, w1715, IN11[6], w1829, w1830);
  FullAdder U296 (w1830, w1717, IN12[6], w1831, w1832);
  FullAdder U297 (w1832, w1719, IN13[6], w1833, w1834);
  FullAdder U298 (w1834, w1721, IN14[6], w1835, w1836);
  FullAdder U299 (w1836, w1723, IN15[6], w1837, w1838);
  FullAdder U300 (w1838, w1725, IN16[6], w1839, w1840);
  FullAdder U301 (w1840, w1727, IN17[6], w1841, w1842);
  FullAdder U302 (w1842, w1729, IN18[6], w1843, w1844);
  FullAdder U303 (w1844, w1731, IN19[6], w1845, w1846);
  FullAdder U304 (w1846, w1733, IN20[6], w1847, w1848);
  FullAdder U305 (w1848, w1735, IN21[6], w1849, w1850);
  FullAdder U306 (w1850, w1737, IN22[6], w1851, w1852);
  FullAdder U307 (w1852, w1739, IN23[6], w1853, w1854);
  FullAdder U308 (w1854, w1741, IN24[6], w1855, w1856);
  FullAdder U309 (w1856, w1743, IN25[6], w1857, w1858);
  FullAdder U310 (w1858, w1745, IN26[6], w1859, w1860);
  FullAdder U311 (w1860, w1747, IN27[6], w1861, w1862);
  FullAdder U312 (w1862, w1749, IN28[6], w1863, w1864);
  FullAdder U313 (w1864, w1751, IN29[6], w1865, w1866);
  FullAdder U314 (w1866, w1753, IN30[6], w1867, w1868);
  FullAdder U315 (w1868, w1755, IN31[6], w1869, w1870);
  FullAdder U316 (w1870, w1757, IN32[6], w1871, w1872);
  FullAdder U317 (w1872, w1759, IN33[6], w1873, w1874);
  FullAdder U318 (w1874, w1761, IN34[6], w1875, w1876);
  FullAdder U319 (w1876, w1763, IN35[6], w1877, w1878);
  FullAdder U320 (w1878, w1765, IN36[6], w1879, w1880);
  FullAdder U321 (w1880, w1767, IN37[6], w1881, w1882);
  FullAdder U322 (w1882, w1769, IN38[6], w1883, w1884);
  FullAdder U323 (w1884, w1771, IN39[6], w1885, w1886);
  FullAdder U324 (w1886, w1773, IN40[6], w1887, w1888);
  FullAdder U325 (w1888, w1775, IN41[6], w1889, w1890);
  FullAdder U326 (w1890, w1777, IN42[6], w1891, w1892);
  FullAdder U327 (w1892, w1779, IN43[6], w1893, w1894);
  FullAdder U328 (w1894, w1781, IN44[6], w1895, w1896);
  FullAdder U329 (w1896, w1783, IN45[6], w1897, w1898);
  FullAdder U330 (w1898, w1785, IN46[6], w1899, w1900);
  FullAdder U331 (w1900, w1787, IN47[6], w1901, w1902);
  FullAdder U332 (w1902, w1789, IN48[6], w1903, w1904);
  FullAdder U333 (w1904, w1791, IN49[6], w1905, w1906);
  FullAdder U334 (w1906, w1793, IN50[6], w1907, w1908);
  FullAdder U335 (w1908, w1795, IN51[6], w1909, w1910);
  FullAdder U336 (w1910, w1797, IN52[6], w1911, w1912);
  FullAdder U337 (w1912, w1799, IN53[6], w1913, w1914);
  FullAdder U338 (w1914, w1801, IN54[6], w1915, w1916);
  FullAdder U339 (w1916, w1803, IN55[6], w1917, w1918);
  FullAdder U340 (w1918, w1805, IN56[6], w1919, w1920);
  FullAdder U341 (w1920, w1807, IN57[6], w1921, w1922);
  FullAdder U342 (w1922, w1809, IN58[6], w1923, w1924);
  FullAdder U343 (w1924, w1811, IN59[4], w1925, w1926);
  FullAdder U344 (w1926, w1813, IN60[3], w1927, w1928);
  FullAdder U345 (w1928, w1815, IN61[2], w1929, w1930);
  FullAdder U346 (w1930, w1817, IN62[1], w1931, w1932);
  FullAdder U347 (w1932, w1818, IN63[0], w1933, w1934);
  HalfAdder U348 (w1821, IN7[7], Out1[7], w1936);
  FullAdder U349 (w1936, w1823, IN8[7], w1937, w1938);
  FullAdder U350 (w1938, w1825, IN9[7], w1939, w1940);
  FullAdder U351 (w1940, w1827, IN10[7], w1941, w1942);
  FullAdder U352 (w1942, w1829, IN11[7], w1943, w1944);
  FullAdder U353 (w1944, w1831, IN12[7], w1945, w1946);
  FullAdder U354 (w1946, w1833, IN13[7], w1947, w1948);
  FullAdder U355 (w1948, w1835, IN14[7], w1949, w1950);
  FullAdder U356 (w1950, w1837, IN15[7], w1951, w1952);
  FullAdder U357 (w1952, w1839, IN16[7], w1953, w1954);
  FullAdder U358 (w1954, w1841, IN17[7], w1955, w1956);
  FullAdder U359 (w1956, w1843, IN18[7], w1957, w1958);
  FullAdder U360 (w1958, w1845, IN19[7], w1959, w1960);
  FullAdder U361 (w1960, w1847, IN20[7], w1961, w1962);
  FullAdder U362 (w1962, w1849, IN21[7], w1963, w1964);
  FullAdder U363 (w1964, w1851, IN22[7], w1965, w1966);
  FullAdder U364 (w1966, w1853, IN23[7], w1967, w1968);
  FullAdder U365 (w1968, w1855, IN24[7], w1969, w1970);
  FullAdder U366 (w1970, w1857, IN25[7], w1971, w1972);
  FullAdder U367 (w1972, w1859, IN26[7], w1973, w1974);
  FullAdder U368 (w1974, w1861, IN27[7], w1975, w1976);
  FullAdder U369 (w1976, w1863, IN28[7], w1977, w1978);
  FullAdder U370 (w1978, w1865, IN29[7], w1979, w1980);
  FullAdder U371 (w1980, w1867, IN30[7], w1981, w1982);
  FullAdder U372 (w1982, w1869, IN31[7], w1983, w1984);
  FullAdder U373 (w1984, w1871, IN32[7], w1985, w1986);
  FullAdder U374 (w1986, w1873, IN33[7], w1987, w1988);
  FullAdder U375 (w1988, w1875, IN34[7], w1989, w1990);
  FullAdder U376 (w1990, w1877, IN35[7], w1991, w1992);
  FullAdder U377 (w1992, w1879, IN36[7], w1993, w1994);
  FullAdder U378 (w1994, w1881, IN37[7], w1995, w1996);
  FullAdder U379 (w1996, w1883, IN38[7], w1997, w1998);
  FullAdder U380 (w1998, w1885, IN39[7], w1999, w2000);
  FullAdder U381 (w2000, w1887, IN40[7], w2001, w2002);
  FullAdder U382 (w2002, w1889, IN41[7], w2003, w2004);
  FullAdder U383 (w2004, w1891, IN42[7], w2005, w2006);
  FullAdder U384 (w2006, w1893, IN43[7], w2007, w2008);
  FullAdder U385 (w2008, w1895, IN44[7], w2009, w2010);
  FullAdder U386 (w2010, w1897, IN45[7], w2011, w2012);
  FullAdder U387 (w2012, w1899, IN46[7], w2013, w2014);
  FullAdder U388 (w2014, w1901, IN47[7], w2015, w2016);
  FullAdder U389 (w2016, w1903, IN48[7], w2017, w2018);
  FullAdder U390 (w2018, w1905, IN49[7], w2019, w2020);
  FullAdder U391 (w2020, w1907, IN50[7], w2021, w2022);
  FullAdder U392 (w2022, w1909, IN51[7], w2023, w2024);
  FullAdder U393 (w2024, w1911, IN52[7], w2025, w2026);
  FullAdder U394 (w2026, w1913, IN53[7], w2027, w2028);
  FullAdder U395 (w2028, w1915, IN54[7], w2029, w2030);
  FullAdder U396 (w2030, w1917, IN55[7], w2031, w2032);
  FullAdder U397 (w2032, w1919, IN56[7], w2033, w2034);
  FullAdder U398 (w2034, w1921, IN57[7], w2035, w2036);
  FullAdder U399 (w2036, w1923, IN58[7], w2037, w2038);
  FullAdder U400 (w2038, w1925, IN59[5], w2039, w2040);
  FullAdder U401 (w2040, w1927, IN60[4], w2041, w2042);
  FullAdder U402 (w2042, w1929, IN61[3], w2043, w2044);
  FullAdder U403 (w2044, w1931, IN62[2], w2045, w2046);
  FullAdder U404 (w2046, w1933, IN63[1], w2047, w2048);
  FullAdder U405 (w2048, w1934, IN64[0], w2049, w2050);
  HalfAdder U406 (w1937, IN8[8], Out1[8], w2052);
  FullAdder U407 (w2052, w1939, IN9[8], w2053, w2054);
  FullAdder U408 (w2054, w1941, IN10[8], w2055, w2056);
  FullAdder U409 (w2056, w1943, IN11[8], w2057, w2058);
  FullAdder U410 (w2058, w1945, IN12[8], w2059, w2060);
  FullAdder U411 (w2060, w1947, IN13[8], w2061, w2062);
  FullAdder U412 (w2062, w1949, IN14[8], w2063, w2064);
  FullAdder U413 (w2064, w1951, IN15[8], w2065, w2066);
  FullAdder U414 (w2066, w1953, IN16[8], w2067, w2068);
  FullAdder U415 (w2068, w1955, IN17[8], w2069, w2070);
  FullAdder U416 (w2070, w1957, IN18[8], w2071, w2072);
  FullAdder U417 (w2072, w1959, IN19[8], w2073, w2074);
  FullAdder U418 (w2074, w1961, IN20[8], w2075, w2076);
  FullAdder U419 (w2076, w1963, IN21[8], w2077, w2078);
  FullAdder U420 (w2078, w1965, IN22[8], w2079, w2080);
  FullAdder U421 (w2080, w1967, IN23[8], w2081, w2082);
  FullAdder U422 (w2082, w1969, IN24[8], w2083, w2084);
  FullAdder U423 (w2084, w1971, IN25[8], w2085, w2086);
  FullAdder U424 (w2086, w1973, IN26[8], w2087, w2088);
  FullAdder U425 (w2088, w1975, IN27[8], w2089, w2090);
  FullAdder U426 (w2090, w1977, IN28[8], w2091, w2092);
  FullAdder U427 (w2092, w1979, IN29[8], w2093, w2094);
  FullAdder U428 (w2094, w1981, IN30[8], w2095, w2096);
  FullAdder U429 (w2096, w1983, IN31[8], w2097, w2098);
  FullAdder U430 (w2098, w1985, IN32[8], w2099, w2100);
  FullAdder U431 (w2100, w1987, IN33[8], w2101, w2102);
  FullAdder U432 (w2102, w1989, IN34[8], w2103, w2104);
  FullAdder U433 (w2104, w1991, IN35[8], w2105, w2106);
  FullAdder U434 (w2106, w1993, IN36[8], w2107, w2108);
  FullAdder U435 (w2108, w1995, IN37[8], w2109, w2110);
  FullAdder U436 (w2110, w1997, IN38[8], w2111, w2112);
  FullAdder U437 (w2112, w1999, IN39[8], w2113, w2114);
  FullAdder U438 (w2114, w2001, IN40[8], w2115, w2116);
  FullAdder U439 (w2116, w2003, IN41[8], w2117, w2118);
  FullAdder U440 (w2118, w2005, IN42[8], w2119, w2120);
  FullAdder U441 (w2120, w2007, IN43[8], w2121, w2122);
  FullAdder U442 (w2122, w2009, IN44[8], w2123, w2124);
  FullAdder U443 (w2124, w2011, IN45[8], w2125, w2126);
  FullAdder U444 (w2126, w2013, IN46[8], w2127, w2128);
  FullAdder U445 (w2128, w2015, IN47[8], w2129, w2130);
  FullAdder U446 (w2130, w2017, IN48[8], w2131, w2132);
  FullAdder U447 (w2132, w2019, IN49[8], w2133, w2134);
  FullAdder U448 (w2134, w2021, IN50[8], w2135, w2136);
  FullAdder U449 (w2136, w2023, IN51[8], w2137, w2138);
  FullAdder U450 (w2138, w2025, IN52[8], w2139, w2140);
  FullAdder U451 (w2140, w2027, IN53[8], w2141, w2142);
  FullAdder U452 (w2142, w2029, IN54[8], w2143, w2144);
  FullAdder U453 (w2144, w2031, IN55[8], w2145, w2146);
  FullAdder U454 (w2146, w2033, IN56[8], w2147, w2148);
  FullAdder U455 (w2148, w2035, IN57[8], w2149, w2150);
  FullAdder U456 (w2150, w2037, IN58[8], w2151, w2152);
  FullAdder U457 (w2152, w2039, IN59[6], w2153, w2154);
  FullAdder U458 (w2154, w2041, IN60[5], w2155, w2156);
  FullAdder U459 (w2156, w2043, IN61[4], w2157, w2158);
  FullAdder U460 (w2158, w2045, IN62[3], w2159, w2160);
  FullAdder U461 (w2160, w2047, IN63[2], w2161, w2162);
  FullAdder U462 (w2162, w2049, IN64[1], w2163, w2164);
  FullAdder U463 (w2164, w2050, IN65[0], w2165, w2166);
  HalfAdder U464 (w2053, IN9[9], Out1[9], w2168);
  FullAdder U465 (w2168, w2055, IN10[9], w2169, w2170);
  FullAdder U466 (w2170, w2057, IN11[9], w2171, w2172);
  FullAdder U467 (w2172, w2059, IN12[9], w2173, w2174);
  FullAdder U468 (w2174, w2061, IN13[9], w2175, w2176);
  FullAdder U469 (w2176, w2063, IN14[9], w2177, w2178);
  FullAdder U470 (w2178, w2065, IN15[9], w2179, w2180);
  FullAdder U471 (w2180, w2067, IN16[9], w2181, w2182);
  FullAdder U472 (w2182, w2069, IN17[9], w2183, w2184);
  FullAdder U473 (w2184, w2071, IN18[9], w2185, w2186);
  FullAdder U474 (w2186, w2073, IN19[9], w2187, w2188);
  FullAdder U475 (w2188, w2075, IN20[9], w2189, w2190);
  FullAdder U476 (w2190, w2077, IN21[9], w2191, w2192);
  FullAdder U477 (w2192, w2079, IN22[9], w2193, w2194);
  FullAdder U478 (w2194, w2081, IN23[9], w2195, w2196);
  FullAdder U479 (w2196, w2083, IN24[9], w2197, w2198);
  FullAdder U480 (w2198, w2085, IN25[9], w2199, w2200);
  FullAdder U481 (w2200, w2087, IN26[9], w2201, w2202);
  FullAdder U482 (w2202, w2089, IN27[9], w2203, w2204);
  FullAdder U483 (w2204, w2091, IN28[9], w2205, w2206);
  FullAdder U484 (w2206, w2093, IN29[9], w2207, w2208);
  FullAdder U485 (w2208, w2095, IN30[9], w2209, w2210);
  FullAdder U486 (w2210, w2097, IN31[9], w2211, w2212);
  FullAdder U487 (w2212, w2099, IN32[9], w2213, w2214);
  FullAdder U488 (w2214, w2101, IN33[9], w2215, w2216);
  FullAdder U489 (w2216, w2103, IN34[9], w2217, w2218);
  FullAdder U490 (w2218, w2105, IN35[9], w2219, w2220);
  FullAdder U491 (w2220, w2107, IN36[9], w2221, w2222);
  FullAdder U492 (w2222, w2109, IN37[9], w2223, w2224);
  FullAdder U493 (w2224, w2111, IN38[9], w2225, w2226);
  FullAdder U494 (w2226, w2113, IN39[9], w2227, w2228);
  FullAdder U495 (w2228, w2115, IN40[9], w2229, w2230);
  FullAdder U496 (w2230, w2117, IN41[9], w2231, w2232);
  FullAdder U497 (w2232, w2119, IN42[9], w2233, w2234);
  FullAdder U498 (w2234, w2121, IN43[9], w2235, w2236);
  FullAdder U499 (w2236, w2123, IN44[9], w2237, w2238);
  FullAdder U500 (w2238, w2125, IN45[9], w2239, w2240);
  FullAdder U501 (w2240, w2127, IN46[9], w2241, w2242);
  FullAdder U502 (w2242, w2129, IN47[9], w2243, w2244);
  FullAdder U503 (w2244, w2131, IN48[9], w2245, w2246);
  FullAdder U504 (w2246, w2133, IN49[9], w2247, w2248);
  FullAdder U505 (w2248, w2135, IN50[9], w2249, w2250);
  FullAdder U506 (w2250, w2137, IN51[9], w2251, w2252);
  FullAdder U507 (w2252, w2139, IN52[9], w2253, w2254);
  FullAdder U508 (w2254, w2141, IN53[9], w2255, w2256);
  FullAdder U509 (w2256, w2143, IN54[9], w2257, w2258);
  FullAdder U510 (w2258, w2145, IN55[9], w2259, w2260);
  FullAdder U511 (w2260, w2147, IN56[9], w2261, w2262);
  FullAdder U512 (w2262, w2149, IN57[9], w2263, w2264);
  FullAdder U513 (w2264, w2151, IN58[9], w2265, w2266);
  FullAdder U514 (w2266, w2153, IN59[7], w2267, w2268);
  FullAdder U515 (w2268, w2155, IN60[6], w2269, w2270);
  FullAdder U516 (w2270, w2157, IN61[5], w2271, w2272);
  FullAdder U517 (w2272, w2159, IN62[4], w2273, w2274);
  FullAdder U518 (w2274, w2161, IN63[3], w2275, w2276);
  FullAdder U519 (w2276, w2163, IN64[2], w2277, w2278);
  FullAdder U520 (w2278, w2165, IN65[1], w2279, w2280);
  FullAdder U521 (w2280, w2166, IN66[0], w2281, w2282);
  HalfAdder U522 (w2169, IN10[10], Out1[10], w2284);
  FullAdder U523 (w2284, w2171, IN11[10], w2285, w2286);
  FullAdder U524 (w2286, w2173, IN12[10], w2287, w2288);
  FullAdder U525 (w2288, w2175, IN13[10], w2289, w2290);
  FullAdder U526 (w2290, w2177, IN14[10], w2291, w2292);
  FullAdder U527 (w2292, w2179, IN15[10], w2293, w2294);
  FullAdder U528 (w2294, w2181, IN16[10], w2295, w2296);
  FullAdder U529 (w2296, w2183, IN17[10], w2297, w2298);
  FullAdder U530 (w2298, w2185, IN18[10], w2299, w2300);
  FullAdder U531 (w2300, w2187, IN19[10], w2301, w2302);
  FullAdder U532 (w2302, w2189, IN20[10], w2303, w2304);
  FullAdder U533 (w2304, w2191, IN21[10], w2305, w2306);
  FullAdder U534 (w2306, w2193, IN22[10], w2307, w2308);
  FullAdder U535 (w2308, w2195, IN23[10], w2309, w2310);
  FullAdder U536 (w2310, w2197, IN24[10], w2311, w2312);
  FullAdder U537 (w2312, w2199, IN25[10], w2313, w2314);
  FullAdder U538 (w2314, w2201, IN26[10], w2315, w2316);
  FullAdder U539 (w2316, w2203, IN27[10], w2317, w2318);
  FullAdder U540 (w2318, w2205, IN28[10], w2319, w2320);
  FullAdder U541 (w2320, w2207, IN29[10], w2321, w2322);
  FullAdder U542 (w2322, w2209, IN30[10], w2323, w2324);
  FullAdder U543 (w2324, w2211, IN31[10], w2325, w2326);
  FullAdder U544 (w2326, w2213, IN32[10], w2327, w2328);
  FullAdder U545 (w2328, w2215, IN33[10], w2329, w2330);
  FullAdder U546 (w2330, w2217, IN34[10], w2331, w2332);
  FullAdder U547 (w2332, w2219, IN35[10], w2333, w2334);
  FullAdder U548 (w2334, w2221, IN36[10], w2335, w2336);
  FullAdder U549 (w2336, w2223, IN37[10], w2337, w2338);
  FullAdder U550 (w2338, w2225, IN38[10], w2339, w2340);
  FullAdder U551 (w2340, w2227, IN39[10], w2341, w2342);
  FullAdder U552 (w2342, w2229, IN40[10], w2343, w2344);
  FullAdder U553 (w2344, w2231, IN41[10], w2345, w2346);
  FullAdder U554 (w2346, w2233, IN42[10], w2347, w2348);
  FullAdder U555 (w2348, w2235, IN43[10], w2349, w2350);
  FullAdder U556 (w2350, w2237, IN44[10], w2351, w2352);
  FullAdder U557 (w2352, w2239, IN45[10], w2353, w2354);
  FullAdder U558 (w2354, w2241, IN46[10], w2355, w2356);
  FullAdder U559 (w2356, w2243, IN47[10], w2357, w2358);
  FullAdder U560 (w2358, w2245, IN48[10], w2359, w2360);
  FullAdder U561 (w2360, w2247, IN49[10], w2361, w2362);
  FullAdder U562 (w2362, w2249, IN50[10], w2363, w2364);
  FullAdder U563 (w2364, w2251, IN51[10], w2365, w2366);
  FullAdder U564 (w2366, w2253, IN52[10], w2367, w2368);
  FullAdder U565 (w2368, w2255, IN53[10], w2369, w2370);
  FullAdder U566 (w2370, w2257, IN54[10], w2371, w2372);
  FullAdder U567 (w2372, w2259, IN55[10], w2373, w2374);
  FullAdder U568 (w2374, w2261, IN56[10], w2375, w2376);
  FullAdder U569 (w2376, w2263, IN57[10], w2377, w2378);
  FullAdder U570 (w2378, w2265, IN58[10], w2379, w2380);
  FullAdder U571 (w2380, w2267, IN59[8], w2381, w2382);
  FullAdder U572 (w2382, w2269, IN60[7], w2383, w2384);
  FullAdder U573 (w2384, w2271, IN61[6], w2385, w2386);
  FullAdder U574 (w2386, w2273, IN62[5], w2387, w2388);
  FullAdder U575 (w2388, w2275, IN63[4], w2389, w2390);
  FullAdder U576 (w2390, w2277, IN64[3], w2391, w2392);
  FullAdder U577 (w2392, w2279, IN65[2], w2393, w2394);
  FullAdder U578 (w2394, w2281, IN66[1], w2395, w2396);
  FullAdder U579 (w2396, w2282, IN67[0], w2397, w2398);
  HalfAdder U580 (w2285, IN11[11], Out1[11], w2400);
  FullAdder U581 (w2400, w2287, IN12[11], w2401, w2402);
  FullAdder U582 (w2402, w2289, IN13[11], w2403, w2404);
  FullAdder U583 (w2404, w2291, IN14[11], w2405, w2406);
  FullAdder U584 (w2406, w2293, IN15[11], w2407, w2408);
  FullAdder U585 (w2408, w2295, IN16[11], w2409, w2410);
  FullAdder U586 (w2410, w2297, IN17[11], w2411, w2412);
  FullAdder U587 (w2412, w2299, IN18[11], w2413, w2414);
  FullAdder U588 (w2414, w2301, IN19[11], w2415, w2416);
  FullAdder U589 (w2416, w2303, IN20[11], w2417, w2418);
  FullAdder U590 (w2418, w2305, IN21[11], w2419, w2420);
  FullAdder U591 (w2420, w2307, IN22[11], w2421, w2422);
  FullAdder U592 (w2422, w2309, IN23[11], w2423, w2424);
  FullAdder U593 (w2424, w2311, IN24[11], w2425, w2426);
  FullAdder U594 (w2426, w2313, IN25[11], w2427, w2428);
  FullAdder U595 (w2428, w2315, IN26[11], w2429, w2430);
  FullAdder U596 (w2430, w2317, IN27[11], w2431, w2432);
  FullAdder U597 (w2432, w2319, IN28[11], w2433, w2434);
  FullAdder U598 (w2434, w2321, IN29[11], w2435, w2436);
  FullAdder U599 (w2436, w2323, IN30[11], w2437, w2438);
  FullAdder U600 (w2438, w2325, IN31[11], w2439, w2440);
  FullAdder U601 (w2440, w2327, IN32[11], w2441, w2442);
  FullAdder U602 (w2442, w2329, IN33[11], w2443, w2444);
  FullAdder U603 (w2444, w2331, IN34[11], w2445, w2446);
  FullAdder U604 (w2446, w2333, IN35[11], w2447, w2448);
  FullAdder U605 (w2448, w2335, IN36[11], w2449, w2450);
  FullAdder U606 (w2450, w2337, IN37[11], w2451, w2452);
  FullAdder U607 (w2452, w2339, IN38[11], w2453, w2454);
  FullAdder U608 (w2454, w2341, IN39[11], w2455, w2456);
  FullAdder U609 (w2456, w2343, IN40[11], w2457, w2458);
  FullAdder U610 (w2458, w2345, IN41[11], w2459, w2460);
  FullAdder U611 (w2460, w2347, IN42[11], w2461, w2462);
  FullAdder U612 (w2462, w2349, IN43[11], w2463, w2464);
  FullAdder U613 (w2464, w2351, IN44[11], w2465, w2466);
  FullAdder U614 (w2466, w2353, IN45[11], w2467, w2468);
  FullAdder U615 (w2468, w2355, IN46[11], w2469, w2470);
  FullAdder U616 (w2470, w2357, IN47[11], w2471, w2472);
  FullAdder U617 (w2472, w2359, IN48[11], w2473, w2474);
  FullAdder U618 (w2474, w2361, IN49[11], w2475, w2476);
  FullAdder U619 (w2476, w2363, IN50[11], w2477, w2478);
  FullAdder U620 (w2478, w2365, IN51[11], w2479, w2480);
  FullAdder U621 (w2480, w2367, IN52[11], w2481, w2482);
  FullAdder U622 (w2482, w2369, IN53[11], w2483, w2484);
  FullAdder U623 (w2484, w2371, IN54[11], w2485, w2486);
  FullAdder U624 (w2486, w2373, IN55[11], w2487, w2488);
  FullAdder U625 (w2488, w2375, IN56[11], w2489, w2490);
  FullAdder U626 (w2490, w2377, IN57[11], w2491, w2492);
  FullAdder U627 (w2492, w2379, IN58[11], w2493, w2494);
  FullAdder U628 (w2494, w2381, IN59[9], w2495, w2496);
  FullAdder U629 (w2496, w2383, IN60[8], w2497, w2498);
  FullAdder U630 (w2498, w2385, IN61[7], w2499, w2500);
  FullAdder U631 (w2500, w2387, IN62[6], w2501, w2502);
  FullAdder U632 (w2502, w2389, IN63[5], w2503, w2504);
  FullAdder U633 (w2504, w2391, IN64[4], w2505, w2506);
  FullAdder U634 (w2506, w2393, IN65[3], w2507, w2508);
  FullAdder U635 (w2508, w2395, IN66[2], w2509, w2510);
  FullAdder U636 (w2510, w2397, IN67[1], w2511, w2512);
  FullAdder U637 (w2512, w2398, IN68[0], w2513, w2514);
  HalfAdder U638 (w2401, IN12[12], Out1[12], w2516);
  FullAdder U639 (w2516, w2403, IN13[12], w2517, w2518);
  FullAdder U640 (w2518, w2405, IN14[12], w2519, w2520);
  FullAdder U641 (w2520, w2407, IN15[12], w2521, w2522);
  FullAdder U642 (w2522, w2409, IN16[12], w2523, w2524);
  FullAdder U643 (w2524, w2411, IN17[12], w2525, w2526);
  FullAdder U644 (w2526, w2413, IN18[12], w2527, w2528);
  FullAdder U645 (w2528, w2415, IN19[12], w2529, w2530);
  FullAdder U646 (w2530, w2417, IN20[12], w2531, w2532);
  FullAdder U647 (w2532, w2419, IN21[12], w2533, w2534);
  FullAdder U648 (w2534, w2421, IN22[12], w2535, w2536);
  FullAdder U649 (w2536, w2423, IN23[12], w2537, w2538);
  FullAdder U650 (w2538, w2425, IN24[12], w2539, w2540);
  FullAdder U651 (w2540, w2427, IN25[12], w2541, w2542);
  FullAdder U652 (w2542, w2429, IN26[12], w2543, w2544);
  FullAdder U653 (w2544, w2431, IN27[12], w2545, w2546);
  FullAdder U654 (w2546, w2433, IN28[12], w2547, w2548);
  FullAdder U655 (w2548, w2435, IN29[12], w2549, w2550);
  FullAdder U656 (w2550, w2437, IN30[12], w2551, w2552);
  FullAdder U657 (w2552, w2439, IN31[12], w2553, w2554);
  FullAdder U658 (w2554, w2441, IN32[12], w2555, w2556);
  FullAdder U659 (w2556, w2443, IN33[12], w2557, w2558);
  FullAdder U660 (w2558, w2445, IN34[12], w2559, w2560);
  FullAdder U661 (w2560, w2447, IN35[12], w2561, w2562);
  FullAdder U662 (w2562, w2449, IN36[12], w2563, w2564);
  FullAdder U663 (w2564, w2451, IN37[12], w2565, w2566);
  FullAdder U664 (w2566, w2453, IN38[12], w2567, w2568);
  FullAdder U665 (w2568, w2455, IN39[12], w2569, w2570);
  FullAdder U666 (w2570, w2457, IN40[12], w2571, w2572);
  FullAdder U667 (w2572, w2459, IN41[12], w2573, w2574);
  FullAdder U668 (w2574, w2461, IN42[12], w2575, w2576);
  FullAdder U669 (w2576, w2463, IN43[12], w2577, w2578);
  FullAdder U670 (w2578, w2465, IN44[12], w2579, w2580);
  FullAdder U671 (w2580, w2467, IN45[12], w2581, w2582);
  FullAdder U672 (w2582, w2469, IN46[12], w2583, w2584);
  FullAdder U673 (w2584, w2471, IN47[12], w2585, w2586);
  FullAdder U674 (w2586, w2473, IN48[12], w2587, w2588);
  FullAdder U675 (w2588, w2475, IN49[12], w2589, w2590);
  FullAdder U676 (w2590, w2477, IN50[12], w2591, w2592);
  FullAdder U677 (w2592, w2479, IN51[12], w2593, w2594);
  FullAdder U678 (w2594, w2481, IN52[12], w2595, w2596);
  FullAdder U679 (w2596, w2483, IN53[12], w2597, w2598);
  FullAdder U680 (w2598, w2485, IN54[12], w2599, w2600);
  FullAdder U681 (w2600, w2487, IN55[12], w2601, w2602);
  FullAdder U682 (w2602, w2489, IN56[12], w2603, w2604);
  FullAdder U683 (w2604, w2491, IN57[12], w2605, w2606);
  FullAdder U684 (w2606, w2493, IN58[12], w2607, w2608);
  FullAdder U685 (w2608, w2495, IN59[10], w2609, w2610);
  FullAdder U686 (w2610, w2497, IN60[9], w2611, w2612);
  FullAdder U687 (w2612, w2499, IN61[8], w2613, w2614);
  FullAdder U688 (w2614, w2501, IN62[7], w2615, w2616);
  FullAdder U689 (w2616, w2503, IN63[6], w2617, w2618);
  FullAdder U690 (w2618, w2505, IN64[5], w2619, w2620);
  FullAdder U691 (w2620, w2507, IN65[4], w2621, w2622);
  FullAdder U692 (w2622, w2509, IN66[3], w2623, w2624);
  FullAdder U693 (w2624, w2511, IN67[2], w2625, w2626);
  FullAdder U694 (w2626, w2513, IN68[1], w2627, w2628);
  FullAdder U695 (w2628, w2514, IN69[0], w2629, w2630);
  HalfAdder U696 (w2517, IN13[13], Out1[13], w2632);
  FullAdder U697 (w2632, w2519, IN14[13], w2633, w2634);
  FullAdder U698 (w2634, w2521, IN15[13], w2635, w2636);
  FullAdder U699 (w2636, w2523, IN16[13], w2637, w2638);
  FullAdder U700 (w2638, w2525, IN17[13], w2639, w2640);
  FullAdder U701 (w2640, w2527, IN18[13], w2641, w2642);
  FullAdder U702 (w2642, w2529, IN19[13], w2643, w2644);
  FullAdder U703 (w2644, w2531, IN20[13], w2645, w2646);
  FullAdder U704 (w2646, w2533, IN21[13], w2647, w2648);
  FullAdder U705 (w2648, w2535, IN22[13], w2649, w2650);
  FullAdder U706 (w2650, w2537, IN23[13], w2651, w2652);
  FullAdder U707 (w2652, w2539, IN24[13], w2653, w2654);
  FullAdder U708 (w2654, w2541, IN25[13], w2655, w2656);
  FullAdder U709 (w2656, w2543, IN26[13], w2657, w2658);
  FullAdder U710 (w2658, w2545, IN27[13], w2659, w2660);
  FullAdder U711 (w2660, w2547, IN28[13], w2661, w2662);
  FullAdder U712 (w2662, w2549, IN29[13], w2663, w2664);
  FullAdder U713 (w2664, w2551, IN30[13], w2665, w2666);
  FullAdder U714 (w2666, w2553, IN31[13], w2667, w2668);
  FullAdder U715 (w2668, w2555, IN32[13], w2669, w2670);
  FullAdder U716 (w2670, w2557, IN33[13], w2671, w2672);
  FullAdder U717 (w2672, w2559, IN34[13], w2673, w2674);
  FullAdder U718 (w2674, w2561, IN35[13], w2675, w2676);
  FullAdder U719 (w2676, w2563, IN36[13], w2677, w2678);
  FullAdder U720 (w2678, w2565, IN37[13], w2679, w2680);
  FullAdder U721 (w2680, w2567, IN38[13], w2681, w2682);
  FullAdder U722 (w2682, w2569, IN39[13], w2683, w2684);
  FullAdder U723 (w2684, w2571, IN40[13], w2685, w2686);
  FullAdder U724 (w2686, w2573, IN41[13], w2687, w2688);
  FullAdder U725 (w2688, w2575, IN42[13], w2689, w2690);
  FullAdder U726 (w2690, w2577, IN43[13], w2691, w2692);
  FullAdder U727 (w2692, w2579, IN44[13], w2693, w2694);
  FullAdder U728 (w2694, w2581, IN45[13], w2695, w2696);
  FullAdder U729 (w2696, w2583, IN46[13], w2697, w2698);
  FullAdder U730 (w2698, w2585, IN47[13], w2699, w2700);
  FullAdder U731 (w2700, w2587, IN48[13], w2701, w2702);
  FullAdder U732 (w2702, w2589, IN49[13], w2703, w2704);
  FullAdder U733 (w2704, w2591, IN50[13], w2705, w2706);
  FullAdder U734 (w2706, w2593, IN51[13], w2707, w2708);
  FullAdder U735 (w2708, w2595, IN52[13], w2709, w2710);
  FullAdder U736 (w2710, w2597, IN53[13], w2711, w2712);
  FullAdder U737 (w2712, w2599, IN54[13], w2713, w2714);
  FullAdder U738 (w2714, w2601, IN55[13], w2715, w2716);
  FullAdder U739 (w2716, w2603, IN56[13], w2717, w2718);
  FullAdder U740 (w2718, w2605, IN57[13], w2719, w2720);
  FullAdder U741 (w2720, w2607, IN58[13], w2721, w2722);
  FullAdder U742 (w2722, w2609, IN59[11], w2723, w2724);
  FullAdder U743 (w2724, w2611, IN60[10], w2725, w2726);
  FullAdder U744 (w2726, w2613, IN61[9], w2727, w2728);
  FullAdder U745 (w2728, w2615, IN62[8], w2729, w2730);
  FullAdder U746 (w2730, w2617, IN63[7], w2731, w2732);
  FullAdder U747 (w2732, w2619, IN64[6], w2733, w2734);
  FullAdder U748 (w2734, w2621, IN65[5], w2735, w2736);
  FullAdder U749 (w2736, w2623, IN66[4], w2737, w2738);
  FullAdder U750 (w2738, w2625, IN67[3], w2739, w2740);
  FullAdder U751 (w2740, w2627, IN68[2], w2741, w2742);
  FullAdder U752 (w2742, w2629, IN69[1], w2743, w2744);
  FullAdder U753 (w2744, w2630, IN70[0], w2745, w2746);
  HalfAdder U754 (w2633, IN14[14], Out1[14], w2748);
  FullAdder U755 (w2748, w2635, IN15[14], w2749, w2750);
  FullAdder U756 (w2750, w2637, IN16[14], w2751, w2752);
  FullAdder U757 (w2752, w2639, IN17[14], w2753, w2754);
  FullAdder U758 (w2754, w2641, IN18[14], w2755, w2756);
  FullAdder U759 (w2756, w2643, IN19[14], w2757, w2758);
  FullAdder U760 (w2758, w2645, IN20[14], w2759, w2760);
  FullAdder U761 (w2760, w2647, IN21[14], w2761, w2762);
  FullAdder U762 (w2762, w2649, IN22[14], w2763, w2764);
  FullAdder U763 (w2764, w2651, IN23[14], w2765, w2766);
  FullAdder U764 (w2766, w2653, IN24[14], w2767, w2768);
  FullAdder U765 (w2768, w2655, IN25[14], w2769, w2770);
  FullAdder U766 (w2770, w2657, IN26[14], w2771, w2772);
  FullAdder U767 (w2772, w2659, IN27[14], w2773, w2774);
  FullAdder U768 (w2774, w2661, IN28[14], w2775, w2776);
  FullAdder U769 (w2776, w2663, IN29[14], w2777, w2778);
  FullAdder U770 (w2778, w2665, IN30[14], w2779, w2780);
  FullAdder U771 (w2780, w2667, IN31[14], w2781, w2782);
  FullAdder U772 (w2782, w2669, IN32[14], w2783, w2784);
  FullAdder U773 (w2784, w2671, IN33[14], w2785, w2786);
  FullAdder U774 (w2786, w2673, IN34[14], w2787, w2788);
  FullAdder U775 (w2788, w2675, IN35[14], w2789, w2790);
  FullAdder U776 (w2790, w2677, IN36[14], w2791, w2792);
  FullAdder U777 (w2792, w2679, IN37[14], w2793, w2794);
  FullAdder U778 (w2794, w2681, IN38[14], w2795, w2796);
  FullAdder U779 (w2796, w2683, IN39[14], w2797, w2798);
  FullAdder U780 (w2798, w2685, IN40[14], w2799, w2800);
  FullAdder U781 (w2800, w2687, IN41[14], w2801, w2802);
  FullAdder U782 (w2802, w2689, IN42[14], w2803, w2804);
  FullAdder U783 (w2804, w2691, IN43[14], w2805, w2806);
  FullAdder U784 (w2806, w2693, IN44[14], w2807, w2808);
  FullAdder U785 (w2808, w2695, IN45[14], w2809, w2810);
  FullAdder U786 (w2810, w2697, IN46[14], w2811, w2812);
  FullAdder U787 (w2812, w2699, IN47[14], w2813, w2814);
  FullAdder U788 (w2814, w2701, IN48[14], w2815, w2816);
  FullAdder U789 (w2816, w2703, IN49[14], w2817, w2818);
  FullAdder U790 (w2818, w2705, IN50[14], w2819, w2820);
  FullAdder U791 (w2820, w2707, IN51[14], w2821, w2822);
  FullAdder U792 (w2822, w2709, IN52[14], w2823, w2824);
  FullAdder U793 (w2824, w2711, IN53[14], w2825, w2826);
  FullAdder U794 (w2826, w2713, IN54[14], w2827, w2828);
  FullAdder U795 (w2828, w2715, IN55[14], w2829, w2830);
  FullAdder U796 (w2830, w2717, IN56[14], w2831, w2832);
  FullAdder U797 (w2832, w2719, IN57[14], w2833, w2834);
  FullAdder U798 (w2834, w2721, IN58[14], w2835, w2836);
  FullAdder U799 (w2836, w2723, IN59[12], w2837, w2838);
  FullAdder U800 (w2838, w2725, IN60[11], w2839, w2840);
  FullAdder U801 (w2840, w2727, IN61[10], w2841, w2842);
  FullAdder U802 (w2842, w2729, IN62[9], w2843, w2844);
  FullAdder U803 (w2844, w2731, IN63[8], w2845, w2846);
  FullAdder U804 (w2846, w2733, IN64[7], w2847, w2848);
  FullAdder U805 (w2848, w2735, IN65[6], w2849, w2850);
  FullAdder U806 (w2850, w2737, IN66[5], w2851, w2852);
  FullAdder U807 (w2852, w2739, IN67[4], w2853, w2854);
  FullAdder U808 (w2854, w2741, IN68[3], w2855, w2856);
  FullAdder U809 (w2856, w2743, IN69[2], w2857, w2858);
  FullAdder U810 (w2858, w2745, IN70[1], w2859, w2860);
  FullAdder U811 (w2860, w2746, IN71[0], w2861, w2862);
  HalfAdder U812 (w2749, IN15[15], Out1[15], w2864);
  FullAdder U813 (w2864, w2751, IN16[15], w2865, w2866);
  FullAdder U814 (w2866, w2753, IN17[15], w2867, w2868);
  FullAdder U815 (w2868, w2755, IN18[15], w2869, w2870);
  FullAdder U816 (w2870, w2757, IN19[15], w2871, w2872);
  FullAdder U817 (w2872, w2759, IN20[15], w2873, w2874);
  FullAdder U818 (w2874, w2761, IN21[15], w2875, w2876);
  FullAdder U819 (w2876, w2763, IN22[15], w2877, w2878);
  FullAdder U820 (w2878, w2765, IN23[15], w2879, w2880);
  FullAdder U821 (w2880, w2767, IN24[15], w2881, w2882);
  FullAdder U822 (w2882, w2769, IN25[15], w2883, w2884);
  FullAdder U823 (w2884, w2771, IN26[15], w2885, w2886);
  FullAdder U824 (w2886, w2773, IN27[15], w2887, w2888);
  FullAdder U825 (w2888, w2775, IN28[15], w2889, w2890);
  FullAdder U826 (w2890, w2777, IN29[15], w2891, w2892);
  FullAdder U827 (w2892, w2779, IN30[15], w2893, w2894);
  FullAdder U828 (w2894, w2781, IN31[15], w2895, w2896);
  FullAdder U829 (w2896, w2783, IN32[15], w2897, w2898);
  FullAdder U830 (w2898, w2785, IN33[15], w2899, w2900);
  FullAdder U831 (w2900, w2787, IN34[15], w2901, w2902);
  FullAdder U832 (w2902, w2789, IN35[15], w2903, w2904);
  FullAdder U833 (w2904, w2791, IN36[15], w2905, w2906);
  FullAdder U834 (w2906, w2793, IN37[15], w2907, w2908);
  FullAdder U835 (w2908, w2795, IN38[15], w2909, w2910);
  FullAdder U836 (w2910, w2797, IN39[15], w2911, w2912);
  FullAdder U837 (w2912, w2799, IN40[15], w2913, w2914);
  FullAdder U838 (w2914, w2801, IN41[15], w2915, w2916);
  FullAdder U839 (w2916, w2803, IN42[15], w2917, w2918);
  FullAdder U840 (w2918, w2805, IN43[15], w2919, w2920);
  FullAdder U841 (w2920, w2807, IN44[15], w2921, w2922);
  FullAdder U842 (w2922, w2809, IN45[15], w2923, w2924);
  FullAdder U843 (w2924, w2811, IN46[15], w2925, w2926);
  FullAdder U844 (w2926, w2813, IN47[15], w2927, w2928);
  FullAdder U845 (w2928, w2815, IN48[15], w2929, w2930);
  FullAdder U846 (w2930, w2817, IN49[15], w2931, w2932);
  FullAdder U847 (w2932, w2819, IN50[15], w2933, w2934);
  FullAdder U848 (w2934, w2821, IN51[15], w2935, w2936);
  FullAdder U849 (w2936, w2823, IN52[15], w2937, w2938);
  FullAdder U850 (w2938, w2825, IN53[15], w2939, w2940);
  FullAdder U851 (w2940, w2827, IN54[15], w2941, w2942);
  FullAdder U852 (w2942, w2829, IN55[15], w2943, w2944);
  FullAdder U853 (w2944, w2831, IN56[15], w2945, w2946);
  FullAdder U854 (w2946, w2833, IN57[15], w2947, w2948);
  FullAdder U855 (w2948, w2835, IN58[15], w2949, w2950);
  FullAdder U856 (w2950, w2837, IN59[13], w2951, w2952);
  FullAdder U857 (w2952, w2839, IN60[12], w2953, w2954);
  FullAdder U858 (w2954, w2841, IN61[11], w2955, w2956);
  FullAdder U859 (w2956, w2843, IN62[10], w2957, w2958);
  FullAdder U860 (w2958, w2845, IN63[9], w2959, w2960);
  FullAdder U861 (w2960, w2847, IN64[8], w2961, w2962);
  FullAdder U862 (w2962, w2849, IN65[7], w2963, w2964);
  FullAdder U863 (w2964, w2851, IN66[6], w2965, w2966);
  FullAdder U864 (w2966, w2853, IN67[5], w2967, w2968);
  FullAdder U865 (w2968, w2855, IN68[4], w2969, w2970);
  FullAdder U866 (w2970, w2857, IN69[3], w2971, w2972);
  FullAdder U867 (w2972, w2859, IN70[2], w2973, w2974);
  FullAdder U868 (w2974, w2861, IN71[1], w2975, w2976);
  FullAdder U869 (w2976, w2862, IN72[0], w2977, w2978);
  HalfAdder U870 (w2865, IN16[16], Out1[16], w2980);
  FullAdder U871 (w2980, w2867, IN17[16], w2981, w2982);
  FullAdder U872 (w2982, w2869, IN18[16], w2983, w2984);
  FullAdder U873 (w2984, w2871, IN19[16], w2985, w2986);
  FullAdder U874 (w2986, w2873, IN20[16], w2987, w2988);
  FullAdder U875 (w2988, w2875, IN21[16], w2989, w2990);
  FullAdder U876 (w2990, w2877, IN22[16], w2991, w2992);
  FullAdder U877 (w2992, w2879, IN23[16], w2993, w2994);
  FullAdder U878 (w2994, w2881, IN24[16], w2995, w2996);
  FullAdder U879 (w2996, w2883, IN25[16], w2997, w2998);
  FullAdder U880 (w2998, w2885, IN26[16], w2999, w3000);
  FullAdder U881 (w3000, w2887, IN27[16], w3001, w3002);
  FullAdder U882 (w3002, w2889, IN28[16], w3003, w3004);
  FullAdder U883 (w3004, w2891, IN29[16], w3005, w3006);
  FullAdder U884 (w3006, w2893, IN30[16], w3007, w3008);
  FullAdder U885 (w3008, w2895, IN31[16], w3009, w3010);
  FullAdder U886 (w3010, w2897, IN32[16], w3011, w3012);
  FullAdder U887 (w3012, w2899, IN33[16], w3013, w3014);
  FullAdder U888 (w3014, w2901, IN34[16], w3015, w3016);
  FullAdder U889 (w3016, w2903, IN35[16], w3017, w3018);
  FullAdder U890 (w3018, w2905, IN36[16], w3019, w3020);
  FullAdder U891 (w3020, w2907, IN37[16], w3021, w3022);
  FullAdder U892 (w3022, w2909, IN38[16], w3023, w3024);
  FullAdder U893 (w3024, w2911, IN39[16], w3025, w3026);
  FullAdder U894 (w3026, w2913, IN40[16], w3027, w3028);
  FullAdder U895 (w3028, w2915, IN41[16], w3029, w3030);
  FullAdder U896 (w3030, w2917, IN42[16], w3031, w3032);
  FullAdder U897 (w3032, w2919, IN43[16], w3033, w3034);
  FullAdder U898 (w3034, w2921, IN44[16], w3035, w3036);
  FullAdder U899 (w3036, w2923, IN45[16], w3037, w3038);
  FullAdder U900 (w3038, w2925, IN46[16], w3039, w3040);
  FullAdder U901 (w3040, w2927, IN47[16], w3041, w3042);
  FullAdder U902 (w3042, w2929, IN48[16], w3043, w3044);
  FullAdder U903 (w3044, w2931, IN49[16], w3045, w3046);
  FullAdder U904 (w3046, w2933, IN50[16], w3047, w3048);
  FullAdder U905 (w3048, w2935, IN51[16], w3049, w3050);
  FullAdder U906 (w3050, w2937, IN52[16], w3051, w3052);
  FullAdder U907 (w3052, w2939, IN53[16], w3053, w3054);
  FullAdder U908 (w3054, w2941, IN54[16], w3055, w3056);
  FullAdder U909 (w3056, w2943, IN55[16], w3057, w3058);
  FullAdder U910 (w3058, w2945, IN56[16], w3059, w3060);
  FullAdder U911 (w3060, w2947, IN57[16], w3061, w3062);
  FullAdder U912 (w3062, w2949, IN58[16], w3063, w3064);
  FullAdder U913 (w3064, w2951, IN59[14], w3065, w3066);
  FullAdder U914 (w3066, w2953, IN60[13], w3067, w3068);
  FullAdder U915 (w3068, w2955, IN61[12], w3069, w3070);
  FullAdder U916 (w3070, w2957, IN62[11], w3071, w3072);
  FullAdder U917 (w3072, w2959, IN63[10], w3073, w3074);
  FullAdder U918 (w3074, w2961, IN64[9], w3075, w3076);
  FullAdder U919 (w3076, w2963, IN65[8], w3077, w3078);
  FullAdder U920 (w3078, w2965, IN66[7], w3079, w3080);
  FullAdder U921 (w3080, w2967, IN67[6], w3081, w3082);
  FullAdder U922 (w3082, w2969, IN68[5], w3083, w3084);
  FullAdder U923 (w3084, w2971, IN69[4], w3085, w3086);
  FullAdder U924 (w3086, w2973, IN70[3], w3087, w3088);
  FullAdder U925 (w3088, w2975, IN71[2], w3089, w3090);
  FullAdder U926 (w3090, w2977, IN72[1], w3091, w3092);
  FullAdder U927 (w3092, w2978, IN73[0], w3093, w3094);
  HalfAdder U928 (w2981, IN17[17], Out1[17], w3096);
  FullAdder U929 (w3096, w2983, IN18[17], w3097, w3098);
  FullAdder U930 (w3098, w2985, IN19[17], w3099, w3100);
  FullAdder U931 (w3100, w2987, IN20[17], w3101, w3102);
  FullAdder U932 (w3102, w2989, IN21[17], w3103, w3104);
  FullAdder U933 (w3104, w2991, IN22[17], w3105, w3106);
  FullAdder U934 (w3106, w2993, IN23[17], w3107, w3108);
  FullAdder U935 (w3108, w2995, IN24[17], w3109, w3110);
  FullAdder U936 (w3110, w2997, IN25[17], w3111, w3112);
  FullAdder U937 (w3112, w2999, IN26[17], w3113, w3114);
  FullAdder U938 (w3114, w3001, IN27[17], w3115, w3116);
  FullAdder U939 (w3116, w3003, IN28[17], w3117, w3118);
  FullAdder U940 (w3118, w3005, IN29[17], w3119, w3120);
  FullAdder U941 (w3120, w3007, IN30[17], w3121, w3122);
  FullAdder U942 (w3122, w3009, IN31[17], w3123, w3124);
  FullAdder U943 (w3124, w3011, IN32[17], w3125, w3126);
  FullAdder U944 (w3126, w3013, IN33[17], w3127, w3128);
  FullAdder U945 (w3128, w3015, IN34[17], w3129, w3130);
  FullAdder U946 (w3130, w3017, IN35[17], w3131, w3132);
  FullAdder U947 (w3132, w3019, IN36[17], w3133, w3134);
  FullAdder U948 (w3134, w3021, IN37[17], w3135, w3136);
  FullAdder U949 (w3136, w3023, IN38[17], w3137, w3138);
  FullAdder U950 (w3138, w3025, IN39[17], w3139, w3140);
  FullAdder U951 (w3140, w3027, IN40[17], w3141, w3142);
  FullAdder U952 (w3142, w3029, IN41[17], w3143, w3144);
  FullAdder U953 (w3144, w3031, IN42[17], w3145, w3146);
  FullAdder U954 (w3146, w3033, IN43[17], w3147, w3148);
  FullAdder U955 (w3148, w3035, IN44[17], w3149, w3150);
  FullAdder U956 (w3150, w3037, IN45[17], w3151, w3152);
  FullAdder U957 (w3152, w3039, IN46[17], w3153, w3154);
  FullAdder U958 (w3154, w3041, IN47[17], w3155, w3156);
  FullAdder U959 (w3156, w3043, IN48[17], w3157, w3158);
  FullAdder U960 (w3158, w3045, IN49[17], w3159, w3160);
  FullAdder U961 (w3160, w3047, IN50[17], w3161, w3162);
  FullAdder U962 (w3162, w3049, IN51[17], w3163, w3164);
  FullAdder U963 (w3164, w3051, IN52[17], w3165, w3166);
  FullAdder U964 (w3166, w3053, IN53[17], w3167, w3168);
  FullAdder U965 (w3168, w3055, IN54[17], w3169, w3170);
  FullAdder U966 (w3170, w3057, IN55[17], w3171, w3172);
  FullAdder U967 (w3172, w3059, IN56[17], w3173, w3174);
  FullAdder U968 (w3174, w3061, IN57[17], w3175, w3176);
  FullAdder U969 (w3176, w3063, IN58[17], w3177, w3178);
  FullAdder U970 (w3178, w3065, IN59[15], w3179, w3180);
  FullAdder U971 (w3180, w3067, IN60[14], w3181, w3182);
  FullAdder U972 (w3182, w3069, IN61[13], w3183, w3184);
  FullAdder U973 (w3184, w3071, IN62[12], w3185, w3186);
  FullAdder U974 (w3186, w3073, IN63[11], w3187, w3188);
  FullAdder U975 (w3188, w3075, IN64[10], w3189, w3190);
  FullAdder U976 (w3190, w3077, IN65[9], w3191, w3192);
  FullAdder U977 (w3192, w3079, IN66[8], w3193, w3194);
  FullAdder U978 (w3194, w3081, IN67[7], w3195, w3196);
  FullAdder U979 (w3196, w3083, IN68[6], w3197, w3198);
  FullAdder U980 (w3198, w3085, IN69[5], w3199, w3200);
  FullAdder U981 (w3200, w3087, IN70[4], w3201, w3202);
  FullAdder U982 (w3202, w3089, IN71[3], w3203, w3204);
  FullAdder U983 (w3204, w3091, IN72[2], w3205, w3206);
  FullAdder U984 (w3206, w3093, IN73[1], w3207, w3208);
  FullAdder U985 (w3208, w3094, IN74[0], w3209, w3210);
  HalfAdder U986 (w3097, IN18[18], Out1[18], w3212);
  FullAdder U987 (w3212, w3099, IN19[18], w3213, w3214);
  FullAdder U988 (w3214, w3101, IN20[18], w3215, w3216);
  FullAdder U989 (w3216, w3103, IN21[18], w3217, w3218);
  FullAdder U990 (w3218, w3105, IN22[18], w3219, w3220);
  FullAdder U991 (w3220, w3107, IN23[18], w3221, w3222);
  FullAdder U992 (w3222, w3109, IN24[18], w3223, w3224);
  FullAdder U993 (w3224, w3111, IN25[18], w3225, w3226);
  FullAdder U994 (w3226, w3113, IN26[18], w3227, w3228);
  FullAdder U995 (w3228, w3115, IN27[18], w3229, w3230);
  FullAdder U996 (w3230, w3117, IN28[18], w3231, w3232);
  FullAdder U997 (w3232, w3119, IN29[18], w3233, w3234);
  FullAdder U998 (w3234, w3121, IN30[18], w3235, w3236);
  FullAdder U999 (w3236, w3123, IN31[18], w3237, w3238);
  FullAdder U1000 (w3238, w3125, IN32[18], w3239, w3240);
  FullAdder U1001 (w3240, w3127, IN33[18], w3241, w3242);
  FullAdder U1002 (w3242, w3129, IN34[18], w3243, w3244);
  FullAdder U1003 (w3244, w3131, IN35[18], w3245, w3246);
  FullAdder U1004 (w3246, w3133, IN36[18], w3247, w3248);
  FullAdder U1005 (w3248, w3135, IN37[18], w3249, w3250);
  FullAdder U1006 (w3250, w3137, IN38[18], w3251, w3252);
  FullAdder U1007 (w3252, w3139, IN39[18], w3253, w3254);
  FullAdder U1008 (w3254, w3141, IN40[18], w3255, w3256);
  FullAdder U1009 (w3256, w3143, IN41[18], w3257, w3258);
  FullAdder U1010 (w3258, w3145, IN42[18], w3259, w3260);
  FullAdder U1011 (w3260, w3147, IN43[18], w3261, w3262);
  FullAdder U1012 (w3262, w3149, IN44[18], w3263, w3264);
  FullAdder U1013 (w3264, w3151, IN45[18], w3265, w3266);
  FullAdder U1014 (w3266, w3153, IN46[18], w3267, w3268);
  FullAdder U1015 (w3268, w3155, IN47[18], w3269, w3270);
  FullAdder U1016 (w3270, w3157, IN48[18], w3271, w3272);
  FullAdder U1017 (w3272, w3159, IN49[18], w3273, w3274);
  FullAdder U1018 (w3274, w3161, IN50[18], w3275, w3276);
  FullAdder U1019 (w3276, w3163, IN51[18], w3277, w3278);
  FullAdder U1020 (w3278, w3165, IN52[18], w3279, w3280);
  FullAdder U1021 (w3280, w3167, IN53[18], w3281, w3282);
  FullAdder U1022 (w3282, w3169, IN54[18], w3283, w3284);
  FullAdder U1023 (w3284, w3171, IN55[18], w3285, w3286);
  FullAdder U1024 (w3286, w3173, IN56[18], w3287, w3288);
  FullAdder U1025 (w3288, w3175, IN57[18], w3289, w3290);
  FullAdder U1026 (w3290, w3177, IN58[18], w3291, w3292);
  FullAdder U1027 (w3292, w3179, IN59[16], w3293, w3294);
  FullAdder U1028 (w3294, w3181, IN60[15], w3295, w3296);
  FullAdder U1029 (w3296, w3183, IN61[14], w3297, w3298);
  FullAdder U1030 (w3298, w3185, IN62[13], w3299, w3300);
  FullAdder U1031 (w3300, w3187, IN63[12], w3301, w3302);
  FullAdder U1032 (w3302, w3189, IN64[11], w3303, w3304);
  FullAdder U1033 (w3304, w3191, IN65[10], w3305, w3306);
  FullAdder U1034 (w3306, w3193, IN66[9], w3307, w3308);
  FullAdder U1035 (w3308, w3195, IN67[8], w3309, w3310);
  FullAdder U1036 (w3310, w3197, IN68[7], w3311, w3312);
  FullAdder U1037 (w3312, w3199, IN69[6], w3313, w3314);
  FullAdder U1038 (w3314, w3201, IN70[5], w3315, w3316);
  FullAdder U1039 (w3316, w3203, IN71[4], w3317, w3318);
  FullAdder U1040 (w3318, w3205, IN72[3], w3319, w3320);
  FullAdder U1041 (w3320, w3207, IN73[2], w3321, w3322);
  FullAdder U1042 (w3322, w3209, IN74[1], w3323, w3324);
  FullAdder U1043 (w3324, w3210, IN75[0], w3325, w3326);
  HalfAdder U1044 (w3213, IN19[19], Out1[19], w3328);
  FullAdder U1045 (w3328, w3215, IN20[19], w3329, w3330);
  FullAdder U1046 (w3330, w3217, IN21[19], w3331, w3332);
  FullAdder U1047 (w3332, w3219, IN22[19], w3333, w3334);
  FullAdder U1048 (w3334, w3221, IN23[19], w3335, w3336);
  FullAdder U1049 (w3336, w3223, IN24[19], w3337, w3338);
  FullAdder U1050 (w3338, w3225, IN25[19], w3339, w3340);
  FullAdder U1051 (w3340, w3227, IN26[19], w3341, w3342);
  FullAdder U1052 (w3342, w3229, IN27[19], w3343, w3344);
  FullAdder U1053 (w3344, w3231, IN28[19], w3345, w3346);
  FullAdder U1054 (w3346, w3233, IN29[19], w3347, w3348);
  FullAdder U1055 (w3348, w3235, IN30[19], w3349, w3350);
  FullAdder U1056 (w3350, w3237, IN31[19], w3351, w3352);
  FullAdder U1057 (w3352, w3239, IN32[19], w3353, w3354);
  FullAdder U1058 (w3354, w3241, IN33[19], w3355, w3356);
  FullAdder U1059 (w3356, w3243, IN34[19], w3357, w3358);
  FullAdder U1060 (w3358, w3245, IN35[19], w3359, w3360);
  FullAdder U1061 (w3360, w3247, IN36[19], w3361, w3362);
  FullAdder U1062 (w3362, w3249, IN37[19], w3363, w3364);
  FullAdder U1063 (w3364, w3251, IN38[19], w3365, w3366);
  FullAdder U1064 (w3366, w3253, IN39[19], w3367, w3368);
  FullAdder U1065 (w3368, w3255, IN40[19], w3369, w3370);
  FullAdder U1066 (w3370, w3257, IN41[19], w3371, w3372);
  FullAdder U1067 (w3372, w3259, IN42[19], w3373, w3374);
  FullAdder U1068 (w3374, w3261, IN43[19], w3375, w3376);
  FullAdder U1069 (w3376, w3263, IN44[19], w3377, w3378);
  FullAdder U1070 (w3378, w3265, IN45[19], w3379, w3380);
  FullAdder U1071 (w3380, w3267, IN46[19], w3381, w3382);
  FullAdder U1072 (w3382, w3269, IN47[19], w3383, w3384);
  FullAdder U1073 (w3384, w3271, IN48[19], w3385, w3386);
  FullAdder U1074 (w3386, w3273, IN49[19], w3387, w3388);
  FullAdder U1075 (w3388, w3275, IN50[19], w3389, w3390);
  FullAdder U1076 (w3390, w3277, IN51[19], w3391, w3392);
  FullAdder U1077 (w3392, w3279, IN52[19], w3393, w3394);
  FullAdder U1078 (w3394, w3281, IN53[19], w3395, w3396);
  FullAdder U1079 (w3396, w3283, IN54[19], w3397, w3398);
  FullAdder U1080 (w3398, w3285, IN55[19], w3399, w3400);
  FullAdder U1081 (w3400, w3287, IN56[19], w3401, w3402);
  FullAdder U1082 (w3402, w3289, IN57[19], w3403, w3404);
  FullAdder U1083 (w3404, w3291, IN58[19], w3405, w3406);
  FullAdder U1084 (w3406, w3293, IN59[17], w3407, w3408);
  FullAdder U1085 (w3408, w3295, IN60[16], w3409, w3410);
  FullAdder U1086 (w3410, w3297, IN61[15], w3411, w3412);
  FullAdder U1087 (w3412, w3299, IN62[14], w3413, w3414);
  FullAdder U1088 (w3414, w3301, IN63[13], w3415, w3416);
  FullAdder U1089 (w3416, w3303, IN64[12], w3417, w3418);
  FullAdder U1090 (w3418, w3305, IN65[11], w3419, w3420);
  FullAdder U1091 (w3420, w3307, IN66[10], w3421, w3422);
  FullAdder U1092 (w3422, w3309, IN67[9], w3423, w3424);
  FullAdder U1093 (w3424, w3311, IN68[8], w3425, w3426);
  FullAdder U1094 (w3426, w3313, IN69[7], w3427, w3428);
  FullAdder U1095 (w3428, w3315, IN70[6], w3429, w3430);
  FullAdder U1096 (w3430, w3317, IN71[5], w3431, w3432);
  FullAdder U1097 (w3432, w3319, IN72[4], w3433, w3434);
  FullAdder U1098 (w3434, w3321, IN73[3], w3435, w3436);
  FullAdder U1099 (w3436, w3323, IN74[2], w3437, w3438);
  FullAdder U1100 (w3438, w3325, IN75[1], w3439, w3440);
  FullAdder U1101 (w3440, w3326, IN76[0], w3441, w3442);
  HalfAdder U1102 (w3329, IN20[20], Out1[20], w3444);
  FullAdder U1103 (w3444, w3331, IN21[20], Out1[21], w3446);
  FullAdder U1104 (w3446, w3333, IN22[20], Out1[22], w3448);
  FullAdder U1105 (w3448, w3335, IN23[20], Out1[23], w3450);
  FullAdder U1106 (w3450, w3337, IN24[20], Out1[24], w3452);
  FullAdder U1107 (w3452, w3339, IN25[20], Out1[25], w3454);
  FullAdder U1108 (w3454, w3341, IN26[20], Out1[26], w3456);
  FullAdder U1109 (w3456, w3343, IN27[20], Out1[27], w3458);
  FullAdder U1110 (w3458, w3345, IN28[20], Out1[28], w3460);
  FullAdder U1111 (w3460, w3347, IN29[20], Out1[29], w3462);
  FullAdder U1112 (w3462, w3349, IN30[20], Out1[30], w3464);
  FullAdder U1113 (w3464, w3351, IN31[20], Out1[31], w3466);
  FullAdder U1114 (w3466, w3353, IN32[20], Out1[32], w3468);
  FullAdder U1115 (w3468, w3355, IN33[20], Out1[33], w3470);
  FullAdder U1116 (w3470, w3357, IN34[20], Out1[34], w3472);
  FullAdder U1117 (w3472, w3359, IN35[20], Out1[35], w3474);
  FullAdder U1118 (w3474, w3361, IN36[20], Out1[36], w3476);
  FullAdder U1119 (w3476, w3363, IN37[20], Out1[37], w3478);
  FullAdder U1120 (w3478, w3365, IN38[20], Out1[38], w3480);
  FullAdder U1121 (w3480, w3367, IN39[20], Out1[39], w3482);
  FullAdder U1122 (w3482, w3369, IN40[20], Out1[40], w3484);
  FullAdder U1123 (w3484, w3371, IN41[20], Out1[41], w3486);
  FullAdder U1124 (w3486, w3373, IN42[20], Out1[42], w3488);
  FullAdder U1125 (w3488, w3375, IN43[20], Out1[43], w3490);
  FullAdder U1126 (w3490, w3377, IN44[20], Out1[44], w3492);
  FullAdder U1127 (w3492, w3379, IN45[20], Out1[45], w3494);
  FullAdder U1128 (w3494, w3381, IN46[20], Out1[46], w3496);
  FullAdder U1129 (w3496, w3383, IN47[20], Out1[47], w3498);
  FullAdder U1130 (w3498, w3385, IN48[20], Out1[48], w3500);
  FullAdder U1131 (w3500, w3387, IN49[20], Out1[49], w3502);
  FullAdder U1132 (w3502, w3389, IN50[20], Out1[50], w3504);
  FullAdder U1133 (w3504, w3391, IN51[20], Out1[51], w3506);
  FullAdder U1134 (w3506, w3393, IN52[20], Out1[52], w3508);
  FullAdder U1135 (w3508, w3395, IN53[20], Out1[53], w3510);
  FullAdder U1136 (w3510, w3397, IN54[20], Out1[54], w3512);
  FullAdder U1137 (w3512, w3399, IN55[20], Out1[55], w3514);
  FullAdder U1138 (w3514, w3401, IN56[20], Out1[56], w3516);
  FullAdder U1139 (w3516, w3403, IN57[20], Out1[57], w3518);
  FullAdder U1140 (w3518, w3405, IN58[20], Out1[58], w3520);
  FullAdder U1141 (w3520, w3407, IN59[18], Out1[59], w3522);
  FullAdder U1142 (w3522, w3409, IN60[17], Out1[60], w3524);
  FullAdder U1143 (w3524, w3411, IN61[16], Out1[61], w3526);
  FullAdder U1144 (w3526, w3413, IN62[15], Out1[62], w3528);
  FullAdder U1145 (w3528, w3415, IN63[14], Out1[63], w3530);
  FullAdder U1146 (w3530, w3417, IN64[13], Out1[64], w3532);
  FullAdder U1147 (w3532, w3419, IN65[12], Out1[65], w3534);
  FullAdder U1148 (w3534, w3421, IN66[11], Out1[66], w3536);
  FullAdder U1149 (w3536, w3423, IN67[10], Out1[67], w3538);
  FullAdder U1150 (w3538, w3425, IN68[9], Out1[68], w3540);
  FullAdder U1151 (w3540, w3427, IN69[8], Out1[69], w3542);
  FullAdder U1152 (w3542, w3429, IN70[7], Out1[70], w3544);
  FullAdder U1153 (w3544, w3431, IN71[6], Out1[71], w3546);
  FullAdder U1154 (w3546, w3433, IN72[5], Out1[72], w3548);
  FullAdder U1155 (w3548, w3435, IN73[4], Out1[73], w3550);
  FullAdder U1156 (w3550, w3437, IN74[3], Out1[74], w3552);
  FullAdder U1157 (w3552, w3439, IN75[2], Out1[75], w3554);
  FullAdder U1158 (w3554, w3441, IN76[1], Out1[76], w3556);
  FullAdder U1159 (w3556, w3442, IN77[0], Out1[77], Out1[78]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN59[19];
  assign Out2[1] = IN60[18];
  assign Out2[2] = IN61[17];
  assign Out2[3] = IN62[16];
  assign Out2[4] = IN63[15];
  assign Out2[5] = IN64[14];
  assign Out2[6] = IN65[13];
  assign Out2[7] = IN66[12];
  assign Out2[8] = IN67[11];
  assign Out2[9] = IN68[10];
  assign Out2[10] = IN69[9];
  assign Out2[11] = IN70[8];
  assign Out2[12] = IN71[7];
  assign Out2[13] = IN72[6];
  assign Out2[14] = IN73[5];
  assign Out2[15] = IN74[4];
  assign Out2[16] = IN75[3];
  assign Out2[17] = IN76[2];
  assign Out2[18] = IN77[1];
  assign Out2[19] = IN78[0];

endmodule
module RC_20_20(IN1, IN2, Out);
  input [19:0] IN1;
  input [19:0] IN2;
  output [20:0] Out;
  wire w41;
  wire w43;
  wire w45;
  wire w47;
  wire w49;
  wire w51;
  wire w53;
  wire w55;
  wire w57;
  wire w59;
  wire w61;
  wire w63;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w41);
  FullAdder U1 (IN1[1], IN2[1], w41, Out[1], w43);
  FullAdder U2 (IN1[2], IN2[2], w43, Out[2], w45);
  FullAdder U3 (IN1[3], IN2[3], w45, Out[3], w47);
  FullAdder U4 (IN1[4], IN2[4], w47, Out[4], w49);
  FullAdder U5 (IN1[5], IN2[5], w49, Out[5], w51);
  FullAdder U6 (IN1[6], IN2[6], w51, Out[6], w53);
  FullAdder U7 (IN1[7], IN2[7], w53, Out[7], w55);
  FullAdder U8 (IN1[8], IN2[8], w55, Out[8], w57);
  FullAdder U9 (IN1[9], IN2[9], w57, Out[9], w59);
  FullAdder U10 (IN1[10], IN2[10], w59, Out[10], w61);
  FullAdder U11 (IN1[11], IN2[11], w61, Out[11], w63);
  FullAdder U12 (IN1[12], IN2[12], w63, Out[12], w65);
  FullAdder U13 (IN1[13], IN2[13], w65, Out[13], w67);
  FullAdder U14 (IN1[14], IN2[14], w67, Out[14], w69);
  FullAdder U15 (IN1[15], IN2[15], w69, Out[15], w71);
  FullAdder U16 (IN1[16], IN2[16], w71, Out[16], w73);
  FullAdder U17 (IN1[17], IN2[17], w73, Out[17], w75);
  FullAdder U18 (IN1[18], IN2[18], w75, Out[18], w77);
  FullAdder U19 (IN1[19], IN2[19], w77, Out[19], Out[20]);

endmodule
module NR_59_21(IN1, IN2, Out);
  input [58:0] IN1;
  input [20:0] IN2;
  output [79:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [20:0] P21;
  wire [20:0] P22;
  wire [20:0] P23;
  wire [20:0] P24;
  wire [20:0] P25;
  wire [20:0] P26;
  wire [20:0] P27;
  wire [20:0] P28;
  wire [20:0] P29;
  wire [20:0] P30;
  wire [20:0] P31;
  wire [20:0] P32;
  wire [20:0] P33;
  wire [20:0] P34;
  wire [20:0] P35;
  wire [20:0] P36;
  wire [20:0] P37;
  wire [20:0] P38;
  wire [20:0] P39;
  wire [20:0] P40;
  wire [20:0] P41;
  wire [20:0] P42;
  wire [20:0] P43;
  wire [20:0] P44;
  wire [20:0] P45;
  wire [20:0] P46;
  wire [20:0] P47;
  wire [20:0] P48;
  wire [20:0] P49;
  wire [20:0] P50;
  wire [20:0] P51;
  wire [20:0] P52;
  wire [20:0] P53;
  wire [20:0] P54;
  wire [20:0] P55;
  wire [20:0] P56;
  wire [20:0] P57;
  wire [20:0] P58;
  wire [19:0] P59;
  wire [18:0] P60;
  wire [17:0] P61;
  wire [16:0] P62;
  wire [15:0] P63;
  wire [14:0] P64;
  wire [13:0] P65;
  wire [12:0] P66;
  wire [11:0] P67;
  wire [10:0] P68;
  wire [9:0] P69;
  wire [8:0] P70;
  wire [7:0] P71;
  wire [6:0] P72;
  wire [5:0] P73;
  wire [4:0] P74;
  wire [3:0] P75;
  wire [2:0] P76;
  wire [1:0] P77;
  wire [0:0] P78;
  wire [78:0] R1;
  wire [19:0] R2;
  wire [79:0] aOut;
  U_SP_59_21 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, R1, R2);
  RC_20_20 S2 (R1[78:59], R2, aOut[79:59]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign aOut[57] = R1[57];
  assign aOut[58] = R1[58];
  assign Out = aOut[79:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
