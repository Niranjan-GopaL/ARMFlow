
module NR_1_38(
    input [0:0]IN1,
    input [37:0]IN2,
    output [37:0]Out
);
    assign Out = IN2;
endmodule
