//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 9
  second input length: 43
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_9_43(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50);
  input [8:0] IN1;
  input [42:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [8:0] P9;
  output [8:0] P10;
  output [8:0] P11;
  output [8:0] P12;
  output [8:0] P13;
  output [8:0] P14;
  output [8:0] P15;
  output [8:0] P16;
  output [8:0] P17;
  output [8:0] P18;
  output [8:0] P19;
  output [8:0] P20;
  output [8:0] P21;
  output [8:0] P22;
  output [8:0] P23;
  output [8:0] P24;
  output [8:0] P25;
  output [8:0] P26;
  output [8:0] P27;
  output [8:0] P28;
  output [8:0] P29;
  output [8:0] P30;
  output [8:0] P31;
  output [8:0] P32;
  output [8:0] P33;
  output [8:0] P34;
  output [8:0] P35;
  output [8:0] P36;
  output [8:0] P37;
  output [8:0] P38;
  output [8:0] P39;
  output [8:0] P40;
  output [8:0] P41;
  output [8:0] P42;
  output [7:0] P43;
  output [6:0] P44;
  output [5:0] P45;
  output [4:0] P46;
  output [3:0] P47;
  output [2:0] P48;
  output [1:0] P49;
  output [0:0] P50;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[0] = IN1[1]&IN2[42];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[1] = IN1[2]&IN2[41];
  assign P44[0] = IN1[2]&IN2[42];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[2] = IN1[3]&IN2[40];
  assign P44[1] = IN1[3]&IN2[41];
  assign P45[0] = IN1[3]&IN2[42];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[3] = IN1[4]&IN2[39];
  assign P44[2] = IN1[4]&IN2[40];
  assign P45[1] = IN1[4]&IN2[41];
  assign P46[0] = IN1[4]&IN2[42];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[4] = IN1[5]&IN2[38];
  assign P44[3] = IN1[5]&IN2[39];
  assign P45[2] = IN1[5]&IN2[40];
  assign P46[1] = IN1[5]&IN2[41];
  assign P47[0] = IN1[5]&IN2[42];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[5] = IN1[6]&IN2[37];
  assign P44[4] = IN1[6]&IN2[38];
  assign P45[3] = IN1[6]&IN2[39];
  assign P46[2] = IN1[6]&IN2[40];
  assign P47[1] = IN1[6]&IN2[41];
  assign P48[0] = IN1[6]&IN2[42];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[6] = IN1[7]&IN2[36];
  assign P44[5] = IN1[7]&IN2[37];
  assign P45[4] = IN1[7]&IN2[38];
  assign P46[3] = IN1[7]&IN2[39];
  assign P47[2] = IN1[7]&IN2[40];
  assign P48[1] = IN1[7]&IN2[41];
  assign P49[0] = IN1[7]&IN2[42];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[7] = IN1[8]&IN2[35];
  assign P44[6] = IN1[8]&IN2[36];
  assign P45[5] = IN1[8]&IN2[37];
  assign P46[4] = IN1[8]&IN2[38];
  assign P47[3] = IN1[8]&IN2[39];
  assign P48[2] = IN1[8]&IN2[40];
  assign P49[1] = IN1[8]&IN2[41];
  assign P50[0] = IN1[8]&IN2[42];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [8:0] IN9;
  input [8:0] IN10;
  input [8:0] IN11;
  input [8:0] IN12;
  input [8:0] IN13;
  input [8:0] IN14;
  input [8:0] IN15;
  input [8:0] IN16;
  input [8:0] IN17;
  input [8:0] IN18;
  input [8:0] IN19;
  input [8:0] IN20;
  input [8:0] IN21;
  input [8:0] IN22;
  input [8:0] IN23;
  input [8:0] IN24;
  input [8:0] IN25;
  input [8:0] IN26;
  input [8:0] IN27;
  input [8:0] IN28;
  input [8:0] IN29;
  input [8:0] IN30;
  input [8:0] IN31;
  input [8:0] IN32;
  input [8:0] IN33;
  input [8:0] IN34;
  input [8:0] IN35;
  input [8:0] IN36;
  input [8:0] IN37;
  input [8:0] IN38;
  input [8:0] IN39;
  input [8:0] IN40;
  input [8:0] IN41;
  input [8:0] IN42;
  input [7:0] IN43;
  input [6:0] IN44;
  input [5:0] IN45;
  input [4:0] IN46;
  input [3:0] IN47;
  input [2:0] IN48;
  input [1:0] IN49;
  input [0:0] IN50;
  output [50:0] Out1;
  output [41:0] Out2;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1044;
  wire w1046;
  wire w1048;
  wire w1050;
  wire w1052;
  wire w1054;
  wire w1056;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w388);
  FullAdder U1 (w388, IN2[0], IN2[1], w389, w390);
  FullAdder U2 (w390, IN3[0], IN3[1], w391, w392);
  FullAdder U3 (w392, IN4[0], IN4[1], w393, w394);
  FullAdder U4 (w394, IN5[0], IN5[1], w395, w396);
  FullAdder U5 (w396, IN6[0], IN6[1], w397, w398);
  FullAdder U6 (w398, IN7[0], IN7[1], w399, w400);
  FullAdder U7 (w400, IN8[0], IN8[1], w401, w402);
  HalfAdder U8 (w389, IN2[2], Out1[2], w404);
  FullAdder U9 (w404, w391, IN3[2], w405, w406);
  FullAdder U10 (w406, w393, IN4[2], w407, w408);
  FullAdder U11 (w408, w395, IN5[2], w409, w410);
  FullAdder U12 (w410, w397, IN6[2], w411, w412);
  FullAdder U13 (w412, w399, IN7[2], w413, w414);
  FullAdder U14 (w414, w401, IN8[2], w415, w416);
  FullAdder U15 (w416, w402, IN9[0], w417, w418);
  HalfAdder U16 (w405, IN3[3], Out1[3], w420);
  FullAdder U17 (w420, w407, IN4[3], w421, w422);
  FullAdder U18 (w422, w409, IN5[3], w423, w424);
  FullAdder U19 (w424, w411, IN6[3], w425, w426);
  FullAdder U20 (w426, w413, IN7[3], w427, w428);
  FullAdder U21 (w428, w415, IN8[3], w429, w430);
  FullAdder U22 (w430, w417, IN9[1], w431, w432);
  FullAdder U23 (w432, w418, IN10[0], w433, w434);
  HalfAdder U24 (w421, IN4[4], Out1[4], w436);
  FullAdder U25 (w436, w423, IN5[4], w437, w438);
  FullAdder U26 (w438, w425, IN6[4], w439, w440);
  FullAdder U27 (w440, w427, IN7[4], w441, w442);
  FullAdder U28 (w442, w429, IN8[4], w443, w444);
  FullAdder U29 (w444, w431, IN9[2], w445, w446);
  FullAdder U30 (w446, w433, IN10[1], w447, w448);
  FullAdder U31 (w448, w434, IN11[0], w449, w450);
  HalfAdder U32 (w437, IN5[5], Out1[5], w452);
  FullAdder U33 (w452, w439, IN6[5], w453, w454);
  FullAdder U34 (w454, w441, IN7[5], w455, w456);
  FullAdder U35 (w456, w443, IN8[5], w457, w458);
  FullAdder U36 (w458, w445, IN9[3], w459, w460);
  FullAdder U37 (w460, w447, IN10[2], w461, w462);
  FullAdder U38 (w462, w449, IN11[1], w463, w464);
  FullAdder U39 (w464, w450, IN12[0], w465, w466);
  HalfAdder U40 (w453, IN6[6], Out1[6], w468);
  FullAdder U41 (w468, w455, IN7[6], w469, w470);
  FullAdder U42 (w470, w457, IN8[6], w471, w472);
  FullAdder U43 (w472, w459, IN9[4], w473, w474);
  FullAdder U44 (w474, w461, IN10[3], w475, w476);
  FullAdder U45 (w476, w463, IN11[2], w477, w478);
  FullAdder U46 (w478, w465, IN12[1], w479, w480);
  FullAdder U47 (w480, w466, IN13[0], w481, w482);
  HalfAdder U48 (w469, IN7[7], Out1[7], w484);
  FullAdder U49 (w484, w471, IN8[7], w485, w486);
  FullAdder U50 (w486, w473, IN9[5], w487, w488);
  FullAdder U51 (w488, w475, IN10[4], w489, w490);
  FullAdder U52 (w490, w477, IN11[3], w491, w492);
  FullAdder U53 (w492, w479, IN12[2], w493, w494);
  FullAdder U54 (w494, w481, IN13[1], w495, w496);
  FullAdder U55 (w496, w482, IN14[0], w497, w498);
  HalfAdder U56 (w485, IN8[8], Out1[8], w500);
  FullAdder U57 (w500, w487, IN9[6], w501, w502);
  FullAdder U58 (w502, w489, IN10[5], w503, w504);
  FullAdder U59 (w504, w491, IN11[4], w505, w506);
  FullAdder U60 (w506, w493, IN12[3], w507, w508);
  FullAdder U61 (w508, w495, IN13[2], w509, w510);
  FullAdder U62 (w510, w497, IN14[1], w511, w512);
  FullAdder U63 (w512, w498, IN15[0], w513, w514);
  HalfAdder U64 (w501, IN9[7], Out1[9], w516);
  FullAdder U65 (w516, w503, IN10[6], w517, w518);
  FullAdder U66 (w518, w505, IN11[5], w519, w520);
  FullAdder U67 (w520, w507, IN12[4], w521, w522);
  FullAdder U68 (w522, w509, IN13[3], w523, w524);
  FullAdder U69 (w524, w511, IN14[2], w525, w526);
  FullAdder U70 (w526, w513, IN15[1], w527, w528);
  FullAdder U71 (w528, w514, IN16[0], w529, w530);
  HalfAdder U72 (w517, IN10[7], Out1[10], w532);
  FullAdder U73 (w532, w519, IN11[6], w533, w534);
  FullAdder U74 (w534, w521, IN12[5], w535, w536);
  FullAdder U75 (w536, w523, IN13[4], w537, w538);
  FullAdder U76 (w538, w525, IN14[3], w539, w540);
  FullAdder U77 (w540, w527, IN15[2], w541, w542);
  FullAdder U78 (w542, w529, IN16[1], w543, w544);
  FullAdder U79 (w544, w530, IN17[0], w545, w546);
  HalfAdder U80 (w533, IN11[7], Out1[11], w548);
  FullAdder U81 (w548, w535, IN12[6], w549, w550);
  FullAdder U82 (w550, w537, IN13[5], w551, w552);
  FullAdder U83 (w552, w539, IN14[4], w553, w554);
  FullAdder U84 (w554, w541, IN15[3], w555, w556);
  FullAdder U85 (w556, w543, IN16[2], w557, w558);
  FullAdder U86 (w558, w545, IN17[1], w559, w560);
  FullAdder U87 (w560, w546, IN18[0], w561, w562);
  HalfAdder U88 (w549, IN12[7], Out1[12], w564);
  FullAdder U89 (w564, w551, IN13[6], w565, w566);
  FullAdder U90 (w566, w553, IN14[5], w567, w568);
  FullAdder U91 (w568, w555, IN15[4], w569, w570);
  FullAdder U92 (w570, w557, IN16[3], w571, w572);
  FullAdder U93 (w572, w559, IN17[2], w573, w574);
  FullAdder U94 (w574, w561, IN18[1], w575, w576);
  FullAdder U95 (w576, w562, IN19[0], w577, w578);
  HalfAdder U96 (w565, IN13[7], Out1[13], w580);
  FullAdder U97 (w580, w567, IN14[6], w581, w582);
  FullAdder U98 (w582, w569, IN15[5], w583, w584);
  FullAdder U99 (w584, w571, IN16[4], w585, w586);
  FullAdder U100 (w586, w573, IN17[3], w587, w588);
  FullAdder U101 (w588, w575, IN18[2], w589, w590);
  FullAdder U102 (w590, w577, IN19[1], w591, w592);
  FullAdder U103 (w592, w578, IN20[0], w593, w594);
  HalfAdder U104 (w581, IN14[7], Out1[14], w596);
  FullAdder U105 (w596, w583, IN15[6], w597, w598);
  FullAdder U106 (w598, w585, IN16[5], w599, w600);
  FullAdder U107 (w600, w587, IN17[4], w601, w602);
  FullAdder U108 (w602, w589, IN18[3], w603, w604);
  FullAdder U109 (w604, w591, IN19[2], w605, w606);
  FullAdder U110 (w606, w593, IN20[1], w607, w608);
  FullAdder U111 (w608, w594, IN21[0], w609, w610);
  HalfAdder U112 (w597, IN15[7], Out1[15], w612);
  FullAdder U113 (w612, w599, IN16[6], w613, w614);
  FullAdder U114 (w614, w601, IN17[5], w615, w616);
  FullAdder U115 (w616, w603, IN18[4], w617, w618);
  FullAdder U116 (w618, w605, IN19[3], w619, w620);
  FullAdder U117 (w620, w607, IN20[2], w621, w622);
  FullAdder U118 (w622, w609, IN21[1], w623, w624);
  FullAdder U119 (w624, w610, IN22[0], w625, w626);
  HalfAdder U120 (w613, IN16[7], Out1[16], w628);
  FullAdder U121 (w628, w615, IN17[6], w629, w630);
  FullAdder U122 (w630, w617, IN18[5], w631, w632);
  FullAdder U123 (w632, w619, IN19[4], w633, w634);
  FullAdder U124 (w634, w621, IN20[3], w635, w636);
  FullAdder U125 (w636, w623, IN21[2], w637, w638);
  FullAdder U126 (w638, w625, IN22[1], w639, w640);
  FullAdder U127 (w640, w626, IN23[0], w641, w642);
  HalfAdder U128 (w629, IN17[7], Out1[17], w644);
  FullAdder U129 (w644, w631, IN18[6], w645, w646);
  FullAdder U130 (w646, w633, IN19[5], w647, w648);
  FullAdder U131 (w648, w635, IN20[4], w649, w650);
  FullAdder U132 (w650, w637, IN21[3], w651, w652);
  FullAdder U133 (w652, w639, IN22[2], w653, w654);
  FullAdder U134 (w654, w641, IN23[1], w655, w656);
  FullAdder U135 (w656, w642, IN24[0], w657, w658);
  HalfAdder U136 (w645, IN18[7], Out1[18], w660);
  FullAdder U137 (w660, w647, IN19[6], w661, w662);
  FullAdder U138 (w662, w649, IN20[5], w663, w664);
  FullAdder U139 (w664, w651, IN21[4], w665, w666);
  FullAdder U140 (w666, w653, IN22[3], w667, w668);
  FullAdder U141 (w668, w655, IN23[2], w669, w670);
  FullAdder U142 (w670, w657, IN24[1], w671, w672);
  FullAdder U143 (w672, w658, IN25[0], w673, w674);
  HalfAdder U144 (w661, IN19[7], Out1[19], w676);
  FullAdder U145 (w676, w663, IN20[6], w677, w678);
  FullAdder U146 (w678, w665, IN21[5], w679, w680);
  FullAdder U147 (w680, w667, IN22[4], w681, w682);
  FullAdder U148 (w682, w669, IN23[3], w683, w684);
  FullAdder U149 (w684, w671, IN24[2], w685, w686);
  FullAdder U150 (w686, w673, IN25[1], w687, w688);
  FullAdder U151 (w688, w674, IN26[0], w689, w690);
  HalfAdder U152 (w677, IN20[7], Out1[20], w692);
  FullAdder U153 (w692, w679, IN21[6], w693, w694);
  FullAdder U154 (w694, w681, IN22[5], w695, w696);
  FullAdder U155 (w696, w683, IN23[4], w697, w698);
  FullAdder U156 (w698, w685, IN24[3], w699, w700);
  FullAdder U157 (w700, w687, IN25[2], w701, w702);
  FullAdder U158 (w702, w689, IN26[1], w703, w704);
  FullAdder U159 (w704, w690, IN27[0], w705, w706);
  HalfAdder U160 (w693, IN21[7], Out1[21], w708);
  FullAdder U161 (w708, w695, IN22[6], w709, w710);
  FullAdder U162 (w710, w697, IN23[5], w711, w712);
  FullAdder U163 (w712, w699, IN24[4], w713, w714);
  FullAdder U164 (w714, w701, IN25[3], w715, w716);
  FullAdder U165 (w716, w703, IN26[2], w717, w718);
  FullAdder U166 (w718, w705, IN27[1], w719, w720);
  FullAdder U167 (w720, w706, IN28[0], w721, w722);
  HalfAdder U168 (w709, IN22[7], Out1[22], w724);
  FullAdder U169 (w724, w711, IN23[6], w725, w726);
  FullAdder U170 (w726, w713, IN24[5], w727, w728);
  FullAdder U171 (w728, w715, IN25[4], w729, w730);
  FullAdder U172 (w730, w717, IN26[3], w731, w732);
  FullAdder U173 (w732, w719, IN27[2], w733, w734);
  FullAdder U174 (w734, w721, IN28[1], w735, w736);
  FullAdder U175 (w736, w722, IN29[0], w737, w738);
  HalfAdder U176 (w725, IN23[7], Out1[23], w740);
  FullAdder U177 (w740, w727, IN24[6], w741, w742);
  FullAdder U178 (w742, w729, IN25[5], w743, w744);
  FullAdder U179 (w744, w731, IN26[4], w745, w746);
  FullAdder U180 (w746, w733, IN27[3], w747, w748);
  FullAdder U181 (w748, w735, IN28[2], w749, w750);
  FullAdder U182 (w750, w737, IN29[1], w751, w752);
  FullAdder U183 (w752, w738, IN30[0], w753, w754);
  HalfAdder U184 (w741, IN24[7], Out1[24], w756);
  FullAdder U185 (w756, w743, IN25[6], w757, w758);
  FullAdder U186 (w758, w745, IN26[5], w759, w760);
  FullAdder U187 (w760, w747, IN27[4], w761, w762);
  FullAdder U188 (w762, w749, IN28[3], w763, w764);
  FullAdder U189 (w764, w751, IN29[2], w765, w766);
  FullAdder U190 (w766, w753, IN30[1], w767, w768);
  FullAdder U191 (w768, w754, IN31[0], w769, w770);
  HalfAdder U192 (w757, IN25[7], Out1[25], w772);
  FullAdder U193 (w772, w759, IN26[6], w773, w774);
  FullAdder U194 (w774, w761, IN27[5], w775, w776);
  FullAdder U195 (w776, w763, IN28[4], w777, w778);
  FullAdder U196 (w778, w765, IN29[3], w779, w780);
  FullAdder U197 (w780, w767, IN30[2], w781, w782);
  FullAdder U198 (w782, w769, IN31[1], w783, w784);
  FullAdder U199 (w784, w770, IN32[0], w785, w786);
  HalfAdder U200 (w773, IN26[7], Out1[26], w788);
  FullAdder U201 (w788, w775, IN27[6], w789, w790);
  FullAdder U202 (w790, w777, IN28[5], w791, w792);
  FullAdder U203 (w792, w779, IN29[4], w793, w794);
  FullAdder U204 (w794, w781, IN30[3], w795, w796);
  FullAdder U205 (w796, w783, IN31[2], w797, w798);
  FullAdder U206 (w798, w785, IN32[1], w799, w800);
  FullAdder U207 (w800, w786, IN33[0], w801, w802);
  HalfAdder U208 (w789, IN27[7], Out1[27], w804);
  FullAdder U209 (w804, w791, IN28[6], w805, w806);
  FullAdder U210 (w806, w793, IN29[5], w807, w808);
  FullAdder U211 (w808, w795, IN30[4], w809, w810);
  FullAdder U212 (w810, w797, IN31[3], w811, w812);
  FullAdder U213 (w812, w799, IN32[2], w813, w814);
  FullAdder U214 (w814, w801, IN33[1], w815, w816);
  FullAdder U215 (w816, w802, IN34[0], w817, w818);
  HalfAdder U216 (w805, IN28[7], Out1[28], w820);
  FullAdder U217 (w820, w807, IN29[6], w821, w822);
  FullAdder U218 (w822, w809, IN30[5], w823, w824);
  FullAdder U219 (w824, w811, IN31[4], w825, w826);
  FullAdder U220 (w826, w813, IN32[3], w827, w828);
  FullAdder U221 (w828, w815, IN33[2], w829, w830);
  FullAdder U222 (w830, w817, IN34[1], w831, w832);
  FullAdder U223 (w832, w818, IN35[0], w833, w834);
  HalfAdder U224 (w821, IN29[7], Out1[29], w836);
  FullAdder U225 (w836, w823, IN30[6], w837, w838);
  FullAdder U226 (w838, w825, IN31[5], w839, w840);
  FullAdder U227 (w840, w827, IN32[4], w841, w842);
  FullAdder U228 (w842, w829, IN33[3], w843, w844);
  FullAdder U229 (w844, w831, IN34[2], w845, w846);
  FullAdder U230 (w846, w833, IN35[1], w847, w848);
  FullAdder U231 (w848, w834, IN36[0], w849, w850);
  HalfAdder U232 (w837, IN30[7], Out1[30], w852);
  FullAdder U233 (w852, w839, IN31[6], w853, w854);
  FullAdder U234 (w854, w841, IN32[5], w855, w856);
  FullAdder U235 (w856, w843, IN33[4], w857, w858);
  FullAdder U236 (w858, w845, IN34[3], w859, w860);
  FullAdder U237 (w860, w847, IN35[2], w861, w862);
  FullAdder U238 (w862, w849, IN36[1], w863, w864);
  FullAdder U239 (w864, w850, IN37[0], w865, w866);
  HalfAdder U240 (w853, IN31[7], Out1[31], w868);
  FullAdder U241 (w868, w855, IN32[6], w869, w870);
  FullAdder U242 (w870, w857, IN33[5], w871, w872);
  FullAdder U243 (w872, w859, IN34[4], w873, w874);
  FullAdder U244 (w874, w861, IN35[3], w875, w876);
  FullAdder U245 (w876, w863, IN36[2], w877, w878);
  FullAdder U246 (w878, w865, IN37[1], w879, w880);
  FullAdder U247 (w880, w866, IN38[0], w881, w882);
  HalfAdder U248 (w869, IN32[7], Out1[32], w884);
  FullAdder U249 (w884, w871, IN33[6], w885, w886);
  FullAdder U250 (w886, w873, IN34[5], w887, w888);
  FullAdder U251 (w888, w875, IN35[4], w889, w890);
  FullAdder U252 (w890, w877, IN36[3], w891, w892);
  FullAdder U253 (w892, w879, IN37[2], w893, w894);
  FullAdder U254 (w894, w881, IN38[1], w895, w896);
  FullAdder U255 (w896, w882, IN39[0], w897, w898);
  HalfAdder U256 (w885, IN33[7], Out1[33], w900);
  FullAdder U257 (w900, w887, IN34[6], w901, w902);
  FullAdder U258 (w902, w889, IN35[5], w903, w904);
  FullAdder U259 (w904, w891, IN36[4], w905, w906);
  FullAdder U260 (w906, w893, IN37[3], w907, w908);
  FullAdder U261 (w908, w895, IN38[2], w909, w910);
  FullAdder U262 (w910, w897, IN39[1], w911, w912);
  FullAdder U263 (w912, w898, IN40[0], w913, w914);
  HalfAdder U264 (w901, IN34[7], Out1[34], w916);
  FullAdder U265 (w916, w903, IN35[6], w917, w918);
  FullAdder U266 (w918, w905, IN36[5], w919, w920);
  FullAdder U267 (w920, w907, IN37[4], w921, w922);
  FullAdder U268 (w922, w909, IN38[3], w923, w924);
  FullAdder U269 (w924, w911, IN39[2], w925, w926);
  FullAdder U270 (w926, w913, IN40[1], w927, w928);
  FullAdder U271 (w928, w914, IN41[0], w929, w930);
  HalfAdder U272 (w917, IN35[7], Out1[35], w932);
  FullAdder U273 (w932, w919, IN36[6], w933, w934);
  FullAdder U274 (w934, w921, IN37[5], w935, w936);
  FullAdder U275 (w936, w923, IN38[4], w937, w938);
  FullAdder U276 (w938, w925, IN39[3], w939, w940);
  FullAdder U277 (w940, w927, IN40[2], w941, w942);
  FullAdder U278 (w942, w929, IN41[1], w943, w944);
  FullAdder U279 (w944, w930, IN42[0], w945, w946);
  HalfAdder U280 (w933, IN36[7], Out1[36], w948);
  FullAdder U281 (w948, w935, IN37[6], w949, w950);
  FullAdder U282 (w950, w937, IN38[5], w951, w952);
  FullAdder U283 (w952, w939, IN39[4], w953, w954);
  FullAdder U284 (w954, w941, IN40[3], w955, w956);
  FullAdder U285 (w956, w943, IN41[2], w957, w958);
  FullAdder U286 (w958, w945, IN42[1], w959, w960);
  FullAdder U287 (w960, w946, IN43[0], w961, w962);
  HalfAdder U288 (w949, IN37[7], Out1[37], w964);
  FullAdder U289 (w964, w951, IN38[6], w965, w966);
  FullAdder U290 (w966, w953, IN39[5], w967, w968);
  FullAdder U291 (w968, w955, IN40[4], w969, w970);
  FullAdder U292 (w970, w957, IN41[3], w971, w972);
  FullAdder U293 (w972, w959, IN42[2], w973, w974);
  FullAdder U294 (w974, w961, IN43[1], w975, w976);
  FullAdder U295 (w976, w962, IN44[0], w977, w978);
  HalfAdder U296 (w965, IN38[7], Out1[38], w980);
  FullAdder U297 (w980, w967, IN39[6], w981, w982);
  FullAdder U298 (w982, w969, IN40[5], w983, w984);
  FullAdder U299 (w984, w971, IN41[4], w985, w986);
  FullAdder U300 (w986, w973, IN42[3], w987, w988);
  FullAdder U301 (w988, w975, IN43[2], w989, w990);
  FullAdder U302 (w990, w977, IN44[1], w991, w992);
  FullAdder U303 (w992, w978, IN45[0], w993, w994);
  HalfAdder U304 (w981, IN39[7], Out1[39], w996);
  FullAdder U305 (w996, w983, IN40[6], w997, w998);
  FullAdder U306 (w998, w985, IN41[5], w999, w1000);
  FullAdder U307 (w1000, w987, IN42[4], w1001, w1002);
  FullAdder U308 (w1002, w989, IN43[3], w1003, w1004);
  FullAdder U309 (w1004, w991, IN44[2], w1005, w1006);
  FullAdder U310 (w1006, w993, IN45[1], w1007, w1008);
  FullAdder U311 (w1008, w994, IN46[0], w1009, w1010);
  HalfAdder U312 (w997, IN40[7], Out1[40], w1012);
  FullAdder U313 (w1012, w999, IN41[6], w1013, w1014);
  FullAdder U314 (w1014, w1001, IN42[5], w1015, w1016);
  FullAdder U315 (w1016, w1003, IN43[4], w1017, w1018);
  FullAdder U316 (w1018, w1005, IN44[3], w1019, w1020);
  FullAdder U317 (w1020, w1007, IN45[2], w1021, w1022);
  FullAdder U318 (w1022, w1009, IN46[1], w1023, w1024);
  FullAdder U319 (w1024, w1010, IN47[0], w1025, w1026);
  HalfAdder U320 (w1013, IN41[7], Out1[41], w1028);
  FullAdder U321 (w1028, w1015, IN42[6], w1029, w1030);
  FullAdder U322 (w1030, w1017, IN43[5], w1031, w1032);
  FullAdder U323 (w1032, w1019, IN44[4], w1033, w1034);
  FullAdder U324 (w1034, w1021, IN45[3], w1035, w1036);
  FullAdder U325 (w1036, w1023, IN46[2], w1037, w1038);
  FullAdder U326 (w1038, w1025, IN47[1], w1039, w1040);
  FullAdder U327 (w1040, w1026, IN48[0], w1041, w1042);
  HalfAdder U328 (w1029, IN42[7], Out1[42], w1044);
  FullAdder U329 (w1044, w1031, IN43[6], Out1[43], w1046);
  FullAdder U330 (w1046, w1033, IN44[5], Out1[44], w1048);
  FullAdder U331 (w1048, w1035, IN45[4], Out1[45], w1050);
  FullAdder U332 (w1050, w1037, IN46[3], Out1[46], w1052);
  FullAdder U333 (w1052, w1039, IN47[2], Out1[47], w1054);
  FullAdder U334 (w1054, w1041, IN48[1], Out1[48], w1056);
  FullAdder U335 (w1056, w1042, IN49[0], Out1[49], Out1[50]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN9[8];
  assign Out2[1] = IN10[8];
  assign Out2[2] = IN11[8];
  assign Out2[3] = IN12[8];
  assign Out2[4] = IN13[8];
  assign Out2[5] = IN14[8];
  assign Out2[6] = IN15[8];
  assign Out2[7] = IN16[8];
  assign Out2[8] = IN17[8];
  assign Out2[9] = IN18[8];
  assign Out2[10] = IN19[8];
  assign Out2[11] = IN20[8];
  assign Out2[12] = IN21[8];
  assign Out2[13] = IN22[8];
  assign Out2[14] = IN23[8];
  assign Out2[15] = IN24[8];
  assign Out2[16] = IN25[8];
  assign Out2[17] = IN26[8];
  assign Out2[18] = IN27[8];
  assign Out2[19] = IN28[8];
  assign Out2[20] = IN29[8];
  assign Out2[21] = IN30[8];
  assign Out2[22] = IN31[8];
  assign Out2[23] = IN32[8];
  assign Out2[24] = IN33[8];
  assign Out2[25] = IN34[8];
  assign Out2[26] = IN35[8];
  assign Out2[27] = IN36[8];
  assign Out2[28] = IN37[8];
  assign Out2[29] = IN38[8];
  assign Out2[30] = IN39[8];
  assign Out2[31] = IN40[8];
  assign Out2[32] = IN41[8];
  assign Out2[33] = IN42[8];
  assign Out2[34] = IN43[7];
  assign Out2[35] = IN44[6];
  assign Out2[36] = IN45[5];
  assign Out2[37] = IN46[4];
  assign Out2[38] = IN47[3];
  assign Out2[39] = IN48[2];
  assign Out2[40] = IN49[1];
  assign Out2[41] = IN50[0];

endmodule
module RC_42_42(IN1, IN2, Out);
  input [41:0] IN1;
  input [41:0] IN2;
  output [42:0] Out;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w85);
  FullAdder U1 (IN1[1], IN2[1], w85, Out[1], w87);
  FullAdder U2 (IN1[2], IN2[2], w87, Out[2], w89);
  FullAdder U3 (IN1[3], IN2[3], w89, Out[3], w91);
  FullAdder U4 (IN1[4], IN2[4], w91, Out[4], w93);
  FullAdder U5 (IN1[5], IN2[5], w93, Out[5], w95);
  FullAdder U6 (IN1[6], IN2[6], w95, Out[6], w97);
  FullAdder U7 (IN1[7], IN2[7], w97, Out[7], w99);
  FullAdder U8 (IN1[8], IN2[8], w99, Out[8], w101);
  FullAdder U9 (IN1[9], IN2[9], w101, Out[9], w103);
  FullAdder U10 (IN1[10], IN2[10], w103, Out[10], w105);
  FullAdder U11 (IN1[11], IN2[11], w105, Out[11], w107);
  FullAdder U12 (IN1[12], IN2[12], w107, Out[12], w109);
  FullAdder U13 (IN1[13], IN2[13], w109, Out[13], w111);
  FullAdder U14 (IN1[14], IN2[14], w111, Out[14], w113);
  FullAdder U15 (IN1[15], IN2[15], w113, Out[15], w115);
  FullAdder U16 (IN1[16], IN2[16], w115, Out[16], w117);
  FullAdder U17 (IN1[17], IN2[17], w117, Out[17], w119);
  FullAdder U18 (IN1[18], IN2[18], w119, Out[18], w121);
  FullAdder U19 (IN1[19], IN2[19], w121, Out[19], w123);
  FullAdder U20 (IN1[20], IN2[20], w123, Out[20], w125);
  FullAdder U21 (IN1[21], IN2[21], w125, Out[21], w127);
  FullAdder U22 (IN1[22], IN2[22], w127, Out[22], w129);
  FullAdder U23 (IN1[23], IN2[23], w129, Out[23], w131);
  FullAdder U24 (IN1[24], IN2[24], w131, Out[24], w133);
  FullAdder U25 (IN1[25], IN2[25], w133, Out[25], w135);
  FullAdder U26 (IN1[26], IN2[26], w135, Out[26], w137);
  FullAdder U27 (IN1[27], IN2[27], w137, Out[27], w139);
  FullAdder U28 (IN1[28], IN2[28], w139, Out[28], w141);
  FullAdder U29 (IN1[29], IN2[29], w141, Out[29], w143);
  FullAdder U30 (IN1[30], IN2[30], w143, Out[30], w145);
  FullAdder U31 (IN1[31], IN2[31], w145, Out[31], w147);
  FullAdder U32 (IN1[32], IN2[32], w147, Out[32], w149);
  FullAdder U33 (IN1[33], IN2[33], w149, Out[33], w151);
  FullAdder U34 (IN1[34], IN2[34], w151, Out[34], w153);
  FullAdder U35 (IN1[35], IN2[35], w153, Out[35], w155);
  FullAdder U36 (IN1[36], IN2[36], w155, Out[36], w157);
  FullAdder U37 (IN1[37], IN2[37], w157, Out[37], w159);
  FullAdder U38 (IN1[38], IN2[38], w159, Out[38], w161);
  FullAdder U39 (IN1[39], IN2[39], w161, Out[39], w163);
  FullAdder U40 (IN1[40], IN2[40], w163, Out[40], w165);
  FullAdder U41 (IN1[41], IN2[41], w165, Out[41], Out[42]);

endmodule
module NR_9_43(IN1, IN2, Out);
  input [8:0] IN1;
  input [42:0] IN2;
  output [51:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [8:0] P9;
  wire [8:0] P10;
  wire [8:0] P11;
  wire [8:0] P12;
  wire [8:0] P13;
  wire [8:0] P14;
  wire [8:0] P15;
  wire [8:0] P16;
  wire [8:0] P17;
  wire [8:0] P18;
  wire [8:0] P19;
  wire [8:0] P20;
  wire [8:0] P21;
  wire [8:0] P22;
  wire [8:0] P23;
  wire [8:0] P24;
  wire [8:0] P25;
  wire [8:0] P26;
  wire [8:0] P27;
  wire [8:0] P28;
  wire [8:0] P29;
  wire [8:0] P30;
  wire [8:0] P31;
  wire [8:0] P32;
  wire [8:0] P33;
  wire [8:0] P34;
  wire [8:0] P35;
  wire [8:0] P36;
  wire [8:0] P37;
  wire [8:0] P38;
  wire [8:0] P39;
  wire [8:0] P40;
  wire [8:0] P41;
  wire [8:0] P42;
  wire [7:0] P43;
  wire [6:0] P44;
  wire [5:0] P45;
  wire [4:0] P46;
  wire [3:0] P47;
  wire [2:0] P48;
  wire [1:0] P49;
  wire [0:0] P50;
  wire [50:0] R1;
  wire [41:0] R2;
  wire [51:0] aOut;
  U_SP_9_43 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, R1, R2);
  RC_42_42 S2 (R1[50:9], R2, aOut[51:9]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign Out = aOut[51:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
