//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 57
  second input length: 6
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_57_6(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61);
  input [56:0] IN1;
  input [5:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [5:0] P6;
  output [5:0] P7;
  output [5:0] P8;
  output [5:0] P9;
  output [5:0] P10;
  output [5:0] P11;
  output [5:0] P12;
  output [5:0] P13;
  output [5:0] P14;
  output [5:0] P15;
  output [5:0] P16;
  output [5:0] P17;
  output [5:0] P18;
  output [5:0] P19;
  output [5:0] P20;
  output [5:0] P21;
  output [5:0] P22;
  output [5:0] P23;
  output [5:0] P24;
  output [5:0] P25;
  output [5:0] P26;
  output [5:0] P27;
  output [5:0] P28;
  output [5:0] P29;
  output [5:0] P30;
  output [5:0] P31;
  output [5:0] P32;
  output [5:0] P33;
  output [5:0] P34;
  output [5:0] P35;
  output [5:0] P36;
  output [5:0] P37;
  output [5:0] P38;
  output [5:0] P39;
  output [5:0] P40;
  output [5:0] P41;
  output [5:0] P42;
  output [5:0] P43;
  output [5:0] P44;
  output [5:0] P45;
  output [5:0] P46;
  output [5:0] P47;
  output [5:0] P48;
  output [5:0] P49;
  output [5:0] P50;
  output [5:0] P51;
  output [5:0] P52;
  output [5:0] P53;
  output [5:0] P54;
  output [5:0] P55;
  output [5:0] P56;
  output [4:0] P57;
  output [3:0] P58;
  output [2:0] P59;
  output [1:0] P60;
  output [0:0] P61;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[0] = IN1[1]&IN2[5];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[1] = IN1[2]&IN2[4];
  assign P7[0] = IN1[2]&IN2[5];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[2] = IN1[3]&IN2[3];
  assign P7[1] = IN1[3]&IN2[4];
  assign P8[0] = IN1[3]&IN2[5];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[3] = IN1[4]&IN2[2];
  assign P7[2] = IN1[4]&IN2[3];
  assign P8[1] = IN1[4]&IN2[4];
  assign P9[0] = IN1[4]&IN2[5];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[4] = IN1[5]&IN2[1];
  assign P7[3] = IN1[5]&IN2[2];
  assign P8[2] = IN1[5]&IN2[3];
  assign P9[1] = IN1[5]&IN2[4];
  assign P10[0] = IN1[5]&IN2[5];
  assign P6[5] = IN1[6]&IN2[0];
  assign P7[4] = IN1[6]&IN2[1];
  assign P8[3] = IN1[6]&IN2[2];
  assign P9[2] = IN1[6]&IN2[3];
  assign P10[1] = IN1[6]&IN2[4];
  assign P11[0] = IN1[6]&IN2[5];
  assign P7[5] = IN1[7]&IN2[0];
  assign P8[4] = IN1[7]&IN2[1];
  assign P9[3] = IN1[7]&IN2[2];
  assign P10[2] = IN1[7]&IN2[3];
  assign P11[1] = IN1[7]&IN2[4];
  assign P12[0] = IN1[7]&IN2[5];
  assign P8[5] = IN1[8]&IN2[0];
  assign P9[4] = IN1[8]&IN2[1];
  assign P10[3] = IN1[8]&IN2[2];
  assign P11[2] = IN1[8]&IN2[3];
  assign P12[1] = IN1[8]&IN2[4];
  assign P13[0] = IN1[8]&IN2[5];
  assign P9[5] = IN1[9]&IN2[0];
  assign P10[4] = IN1[9]&IN2[1];
  assign P11[3] = IN1[9]&IN2[2];
  assign P12[2] = IN1[9]&IN2[3];
  assign P13[1] = IN1[9]&IN2[4];
  assign P14[0] = IN1[9]&IN2[5];
  assign P10[5] = IN1[10]&IN2[0];
  assign P11[4] = IN1[10]&IN2[1];
  assign P12[3] = IN1[10]&IN2[2];
  assign P13[2] = IN1[10]&IN2[3];
  assign P14[1] = IN1[10]&IN2[4];
  assign P15[0] = IN1[10]&IN2[5];
  assign P11[5] = IN1[11]&IN2[0];
  assign P12[4] = IN1[11]&IN2[1];
  assign P13[3] = IN1[11]&IN2[2];
  assign P14[2] = IN1[11]&IN2[3];
  assign P15[1] = IN1[11]&IN2[4];
  assign P16[0] = IN1[11]&IN2[5];
  assign P12[5] = IN1[12]&IN2[0];
  assign P13[4] = IN1[12]&IN2[1];
  assign P14[3] = IN1[12]&IN2[2];
  assign P15[2] = IN1[12]&IN2[3];
  assign P16[1] = IN1[12]&IN2[4];
  assign P17[0] = IN1[12]&IN2[5];
  assign P13[5] = IN1[13]&IN2[0];
  assign P14[4] = IN1[13]&IN2[1];
  assign P15[3] = IN1[13]&IN2[2];
  assign P16[2] = IN1[13]&IN2[3];
  assign P17[1] = IN1[13]&IN2[4];
  assign P18[0] = IN1[13]&IN2[5];
  assign P14[5] = IN1[14]&IN2[0];
  assign P15[4] = IN1[14]&IN2[1];
  assign P16[3] = IN1[14]&IN2[2];
  assign P17[2] = IN1[14]&IN2[3];
  assign P18[1] = IN1[14]&IN2[4];
  assign P19[0] = IN1[14]&IN2[5];
  assign P15[5] = IN1[15]&IN2[0];
  assign P16[4] = IN1[15]&IN2[1];
  assign P17[3] = IN1[15]&IN2[2];
  assign P18[2] = IN1[15]&IN2[3];
  assign P19[1] = IN1[15]&IN2[4];
  assign P20[0] = IN1[15]&IN2[5];
  assign P16[5] = IN1[16]&IN2[0];
  assign P17[4] = IN1[16]&IN2[1];
  assign P18[3] = IN1[16]&IN2[2];
  assign P19[2] = IN1[16]&IN2[3];
  assign P20[1] = IN1[16]&IN2[4];
  assign P21[0] = IN1[16]&IN2[5];
  assign P17[5] = IN1[17]&IN2[0];
  assign P18[4] = IN1[17]&IN2[1];
  assign P19[3] = IN1[17]&IN2[2];
  assign P20[2] = IN1[17]&IN2[3];
  assign P21[1] = IN1[17]&IN2[4];
  assign P22[0] = IN1[17]&IN2[5];
  assign P18[5] = IN1[18]&IN2[0];
  assign P19[4] = IN1[18]&IN2[1];
  assign P20[3] = IN1[18]&IN2[2];
  assign P21[2] = IN1[18]&IN2[3];
  assign P22[1] = IN1[18]&IN2[4];
  assign P23[0] = IN1[18]&IN2[5];
  assign P19[5] = IN1[19]&IN2[0];
  assign P20[4] = IN1[19]&IN2[1];
  assign P21[3] = IN1[19]&IN2[2];
  assign P22[2] = IN1[19]&IN2[3];
  assign P23[1] = IN1[19]&IN2[4];
  assign P24[0] = IN1[19]&IN2[5];
  assign P20[5] = IN1[20]&IN2[0];
  assign P21[4] = IN1[20]&IN2[1];
  assign P22[3] = IN1[20]&IN2[2];
  assign P23[2] = IN1[20]&IN2[3];
  assign P24[1] = IN1[20]&IN2[4];
  assign P25[0] = IN1[20]&IN2[5];
  assign P21[5] = IN1[21]&IN2[0];
  assign P22[4] = IN1[21]&IN2[1];
  assign P23[3] = IN1[21]&IN2[2];
  assign P24[2] = IN1[21]&IN2[3];
  assign P25[1] = IN1[21]&IN2[4];
  assign P26[0] = IN1[21]&IN2[5];
  assign P22[5] = IN1[22]&IN2[0];
  assign P23[4] = IN1[22]&IN2[1];
  assign P24[3] = IN1[22]&IN2[2];
  assign P25[2] = IN1[22]&IN2[3];
  assign P26[1] = IN1[22]&IN2[4];
  assign P27[0] = IN1[22]&IN2[5];
  assign P23[5] = IN1[23]&IN2[0];
  assign P24[4] = IN1[23]&IN2[1];
  assign P25[3] = IN1[23]&IN2[2];
  assign P26[2] = IN1[23]&IN2[3];
  assign P27[1] = IN1[23]&IN2[4];
  assign P28[0] = IN1[23]&IN2[5];
  assign P24[5] = IN1[24]&IN2[0];
  assign P25[4] = IN1[24]&IN2[1];
  assign P26[3] = IN1[24]&IN2[2];
  assign P27[2] = IN1[24]&IN2[3];
  assign P28[1] = IN1[24]&IN2[4];
  assign P29[0] = IN1[24]&IN2[5];
  assign P25[5] = IN1[25]&IN2[0];
  assign P26[4] = IN1[25]&IN2[1];
  assign P27[3] = IN1[25]&IN2[2];
  assign P28[2] = IN1[25]&IN2[3];
  assign P29[1] = IN1[25]&IN2[4];
  assign P30[0] = IN1[25]&IN2[5];
  assign P26[5] = IN1[26]&IN2[0];
  assign P27[4] = IN1[26]&IN2[1];
  assign P28[3] = IN1[26]&IN2[2];
  assign P29[2] = IN1[26]&IN2[3];
  assign P30[1] = IN1[26]&IN2[4];
  assign P31[0] = IN1[26]&IN2[5];
  assign P27[5] = IN1[27]&IN2[0];
  assign P28[4] = IN1[27]&IN2[1];
  assign P29[3] = IN1[27]&IN2[2];
  assign P30[2] = IN1[27]&IN2[3];
  assign P31[1] = IN1[27]&IN2[4];
  assign P32[0] = IN1[27]&IN2[5];
  assign P28[5] = IN1[28]&IN2[0];
  assign P29[4] = IN1[28]&IN2[1];
  assign P30[3] = IN1[28]&IN2[2];
  assign P31[2] = IN1[28]&IN2[3];
  assign P32[1] = IN1[28]&IN2[4];
  assign P33[0] = IN1[28]&IN2[5];
  assign P29[5] = IN1[29]&IN2[0];
  assign P30[4] = IN1[29]&IN2[1];
  assign P31[3] = IN1[29]&IN2[2];
  assign P32[2] = IN1[29]&IN2[3];
  assign P33[1] = IN1[29]&IN2[4];
  assign P34[0] = IN1[29]&IN2[5];
  assign P30[5] = IN1[30]&IN2[0];
  assign P31[4] = IN1[30]&IN2[1];
  assign P32[3] = IN1[30]&IN2[2];
  assign P33[2] = IN1[30]&IN2[3];
  assign P34[1] = IN1[30]&IN2[4];
  assign P35[0] = IN1[30]&IN2[5];
  assign P31[5] = IN1[31]&IN2[0];
  assign P32[4] = IN1[31]&IN2[1];
  assign P33[3] = IN1[31]&IN2[2];
  assign P34[2] = IN1[31]&IN2[3];
  assign P35[1] = IN1[31]&IN2[4];
  assign P36[0] = IN1[31]&IN2[5];
  assign P32[5] = IN1[32]&IN2[0];
  assign P33[4] = IN1[32]&IN2[1];
  assign P34[3] = IN1[32]&IN2[2];
  assign P35[2] = IN1[32]&IN2[3];
  assign P36[1] = IN1[32]&IN2[4];
  assign P37[0] = IN1[32]&IN2[5];
  assign P33[5] = IN1[33]&IN2[0];
  assign P34[4] = IN1[33]&IN2[1];
  assign P35[3] = IN1[33]&IN2[2];
  assign P36[2] = IN1[33]&IN2[3];
  assign P37[1] = IN1[33]&IN2[4];
  assign P38[0] = IN1[33]&IN2[5];
  assign P34[5] = IN1[34]&IN2[0];
  assign P35[4] = IN1[34]&IN2[1];
  assign P36[3] = IN1[34]&IN2[2];
  assign P37[2] = IN1[34]&IN2[3];
  assign P38[1] = IN1[34]&IN2[4];
  assign P39[0] = IN1[34]&IN2[5];
  assign P35[5] = IN1[35]&IN2[0];
  assign P36[4] = IN1[35]&IN2[1];
  assign P37[3] = IN1[35]&IN2[2];
  assign P38[2] = IN1[35]&IN2[3];
  assign P39[1] = IN1[35]&IN2[4];
  assign P40[0] = IN1[35]&IN2[5];
  assign P36[5] = IN1[36]&IN2[0];
  assign P37[4] = IN1[36]&IN2[1];
  assign P38[3] = IN1[36]&IN2[2];
  assign P39[2] = IN1[36]&IN2[3];
  assign P40[1] = IN1[36]&IN2[4];
  assign P41[0] = IN1[36]&IN2[5];
  assign P37[5] = IN1[37]&IN2[0];
  assign P38[4] = IN1[37]&IN2[1];
  assign P39[3] = IN1[37]&IN2[2];
  assign P40[2] = IN1[37]&IN2[3];
  assign P41[1] = IN1[37]&IN2[4];
  assign P42[0] = IN1[37]&IN2[5];
  assign P38[5] = IN1[38]&IN2[0];
  assign P39[4] = IN1[38]&IN2[1];
  assign P40[3] = IN1[38]&IN2[2];
  assign P41[2] = IN1[38]&IN2[3];
  assign P42[1] = IN1[38]&IN2[4];
  assign P43[0] = IN1[38]&IN2[5];
  assign P39[5] = IN1[39]&IN2[0];
  assign P40[4] = IN1[39]&IN2[1];
  assign P41[3] = IN1[39]&IN2[2];
  assign P42[2] = IN1[39]&IN2[3];
  assign P43[1] = IN1[39]&IN2[4];
  assign P44[0] = IN1[39]&IN2[5];
  assign P40[5] = IN1[40]&IN2[0];
  assign P41[4] = IN1[40]&IN2[1];
  assign P42[3] = IN1[40]&IN2[2];
  assign P43[2] = IN1[40]&IN2[3];
  assign P44[1] = IN1[40]&IN2[4];
  assign P45[0] = IN1[40]&IN2[5];
  assign P41[5] = IN1[41]&IN2[0];
  assign P42[4] = IN1[41]&IN2[1];
  assign P43[3] = IN1[41]&IN2[2];
  assign P44[2] = IN1[41]&IN2[3];
  assign P45[1] = IN1[41]&IN2[4];
  assign P46[0] = IN1[41]&IN2[5];
  assign P42[5] = IN1[42]&IN2[0];
  assign P43[4] = IN1[42]&IN2[1];
  assign P44[3] = IN1[42]&IN2[2];
  assign P45[2] = IN1[42]&IN2[3];
  assign P46[1] = IN1[42]&IN2[4];
  assign P47[0] = IN1[42]&IN2[5];
  assign P43[5] = IN1[43]&IN2[0];
  assign P44[4] = IN1[43]&IN2[1];
  assign P45[3] = IN1[43]&IN2[2];
  assign P46[2] = IN1[43]&IN2[3];
  assign P47[1] = IN1[43]&IN2[4];
  assign P48[0] = IN1[43]&IN2[5];
  assign P44[5] = IN1[44]&IN2[0];
  assign P45[4] = IN1[44]&IN2[1];
  assign P46[3] = IN1[44]&IN2[2];
  assign P47[2] = IN1[44]&IN2[3];
  assign P48[1] = IN1[44]&IN2[4];
  assign P49[0] = IN1[44]&IN2[5];
  assign P45[5] = IN1[45]&IN2[0];
  assign P46[4] = IN1[45]&IN2[1];
  assign P47[3] = IN1[45]&IN2[2];
  assign P48[2] = IN1[45]&IN2[3];
  assign P49[1] = IN1[45]&IN2[4];
  assign P50[0] = IN1[45]&IN2[5];
  assign P46[5] = IN1[46]&IN2[0];
  assign P47[4] = IN1[46]&IN2[1];
  assign P48[3] = IN1[46]&IN2[2];
  assign P49[2] = IN1[46]&IN2[3];
  assign P50[1] = IN1[46]&IN2[4];
  assign P51[0] = IN1[46]&IN2[5];
  assign P47[5] = IN1[47]&IN2[0];
  assign P48[4] = IN1[47]&IN2[1];
  assign P49[3] = IN1[47]&IN2[2];
  assign P50[2] = IN1[47]&IN2[3];
  assign P51[1] = IN1[47]&IN2[4];
  assign P52[0] = IN1[47]&IN2[5];
  assign P48[5] = IN1[48]&IN2[0];
  assign P49[4] = IN1[48]&IN2[1];
  assign P50[3] = IN1[48]&IN2[2];
  assign P51[2] = IN1[48]&IN2[3];
  assign P52[1] = IN1[48]&IN2[4];
  assign P53[0] = IN1[48]&IN2[5];
  assign P49[5] = IN1[49]&IN2[0];
  assign P50[4] = IN1[49]&IN2[1];
  assign P51[3] = IN1[49]&IN2[2];
  assign P52[2] = IN1[49]&IN2[3];
  assign P53[1] = IN1[49]&IN2[4];
  assign P54[0] = IN1[49]&IN2[5];
  assign P50[5] = IN1[50]&IN2[0];
  assign P51[4] = IN1[50]&IN2[1];
  assign P52[3] = IN1[50]&IN2[2];
  assign P53[2] = IN1[50]&IN2[3];
  assign P54[1] = IN1[50]&IN2[4];
  assign P55[0] = IN1[50]&IN2[5];
  assign P51[5] = IN1[51]&IN2[0];
  assign P52[4] = IN1[51]&IN2[1];
  assign P53[3] = IN1[51]&IN2[2];
  assign P54[2] = IN1[51]&IN2[3];
  assign P55[1] = IN1[51]&IN2[4];
  assign P56[0] = IN1[51]&IN2[5];
  assign P52[5] = IN1[52]&IN2[0];
  assign P53[4] = IN1[52]&IN2[1];
  assign P54[3] = IN1[52]&IN2[2];
  assign P55[2] = IN1[52]&IN2[3];
  assign P56[1] = IN1[52]&IN2[4];
  assign P57[0] = IN1[52]&IN2[5];
  assign P53[5] = IN1[53]&IN2[0];
  assign P54[4] = IN1[53]&IN2[1];
  assign P55[3] = IN1[53]&IN2[2];
  assign P56[2] = IN1[53]&IN2[3];
  assign P57[1] = IN1[53]&IN2[4];
  assign P58[0] = IN1[53]&IN2[5];
  assign P54[5] = IN1[54]&IN2[0];
  assign P55[4] = IN1[54]&IN2[1];
  assign P56[3] = IN1[54]&IN2[2];
  assign P57[2] = IN1[54]&IN2[3];
  assign P58[1] = IN1[54]&IN2[4];
  assign P59[0] = IN1[54]&IN2[5];
  assign P55[5] = IN1[55]&IN2[0];
  assign P56[4] = IN1[55]&IN2[1];
  assign P57[3] = IN1[55]&IN2[2];
  assign P58[2] = IN1[55]&IN2[3];
  assign P59[1] = IN1[55]&IN2[4];
  assign P60[0] = IN1[55]&IN2[5];
  assign P56[5] = IN1[56]&IN2[0];
  assign P57[4] = IN1[56]&IN2[1];
  assign P58[3] = IN1[56]&IN2[2];
  assign P59[2] = IN1[56]&IN2[3];
  assign P60[1] = IN1[56]&IN2[4];
  assign P61[0] = IN1[56]&IN2[5];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [5:0] IN6;
  input [5:0] IN7;
  input [5:0] IN8;
  input [5:0] IN9;
  input [5:0] IN10;
  input [5:0] IN11;
  input [5:0] IN12;
  input [5:0] IN13;
  input [5:0] IN14;
  input [5:0] IN15;
  input [5:0] IN16;
  input [5:0] IN17;
  input [5:0] IN18;
  input [5:0] IN19;
  input [5:0] IN20;
  input [5:0] IN21;
  input [5:0] IN22;
  input [5:0] IN23;
  input [5:0] IN24;
  input [5:0] IN25;
  input [5:0] IN26;
  input [5:0] IN27;
  input [5:0] IN28;
  input [5:0] IN29;
  input [5:0] IN30;
  input [5:0] IN31;
  input [5:0] IN32;
  input [5:0] IN33;
  input [5:0] IN34;
  input [5:0] IN35;
  input [5:0] IN36;
  input [5:0] IN37;
  input [5:0] IN38;
  input [5:0] IN39;
  input [5:0] IN40;
  input [5:0] IN41;
  input [5:0] IN42;
  input [5:0] IN43;
  input [5:0] IN44;
  input [5:0] IN45;
  input [5:0] IN46;
  input [5:0] IN47;
  input [5:0] IN48;
  input [5:0] IN49;
  input [5:0] IN50;
  input [5:0] IN51;
  input [5:0] IN52;
  input [5:0] IN53;
  input [5:0] IN54;
  input [5:0] IN55;
  input [5:0] IN56;
  input [4:0] IN57;
  input [3:0] IN58;
  input [2:0] IN59;
  input [1:0] IN60;
  input [0:0] IN61;
  output [61:0] Out1;
  output [4:0] Out2;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w791;
  wire w793;
  wire w795;
  wire w797;
  wire w799;
  wire w801;
  wire w803;
  wire w805;
  wire w807;
  wire w809;
  wire w811;
  wire w813;
  wire w815;
  wire w817;
  wire w819;
  wire w821;
  wire w823;
  wire w825;
  wire w827;
  wire w829;
  wire w831;
  wire w833;
  wire w835;
  wire w837;
  wire w839;
  wire w841;
  wire w843;
  wire w845;
  wire w847;
  wire w849;
  wire w851;
  wire w853;
  wire w855;
  wire w857;
  wire w859;
  wire w861;
  wire w863;
  wire w865;
  wire w867;
  wire w869;
  wire w871;
  wire w873;
  wire w875;
  wire w877;
  wire w879;
  wire w881;
  wire w883;
  wire w885;
  wire w887;
  wire w889;
  wire w891;
  wire w893;
  wire w895;
  wire w897;
  wire w899;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w343);
  FullAdder U1 (w343, IN2[0], IN2[1], w344, w345);
  FullAdder U2 (w345, IN3[0], IN3[1], w346, w347);
  FullAdder U3 (w347, IN4[0], IN4[1], w348, w349);
  FullAdder U4 (w349, IN5[0], IN5[1], w350, w351);
  FullAdder U5 (w351, IN6[0], IN6[1], w352, w353);
  FullAdder U6 (w353, IN7[0], IN7[1], w354, w355);
  FullAdder U7 (w355, IN8[0], IN8[1], w356, w357);
  FullAdder U8 (w357, IN9[0], IN9[1], w358, w359);
  FullAdder U9 (w359, IN10[0], IN10[1], w360, w361);
  FullAdder U10 (w361, IN11[0], IN11[1], w362, w363);
  FullAdder U11 (w363, IN12[0], IN12[1], w364, w365);
  FullAdder U12 (w365, IN13[0], IN13[1], w366, w367);
  FullAdder U13 (w367, IN14[0], IN14[1], w368, w369);
  FullAdder U14 (w369, IN15[0], IN15[1], w370, w371);
  FullAdder U15 (w371, IN16[0], IN16[1], w372, w373);
  FullAdder U16 (w373, IN17[0], IN17[1], w374, w375);
  FullAdder U17 (w375, IN18[0], IN18[1], w376, w377);
  FullAdder U18 (w377, IN19[0], IN19[1], w378, w379);
  FullAdder U19 (w379, IN20[0], IN20[1], w380, w381);
  FullAdder U20 (w381, IN21[0], IN21[1], w382, w383);
  FullAdder U21 (w383, IN22[0], IN22[1], w384, w385);
  FullAdder U22 (w385, IN23[0], IN23[1], w386, w387);
  FullAdder U23 (w387, IN24[0], IN24[1], w388, w389);
  FullAdder U24 (w389, IN25[0], IN25[1], w390, w391);
  FullAdder U25 (w391, IN26[0], IN26[1], w392, w393);
  FullAdder U26 (w393, IN27[0], IN27[1], w394, w395);
  FullAdder U27 (w395, IN28[0], IN28[1], w396, w397);
  FullAdder U28 (w397, IN29[0], IN29[1], w398, w399);
  FullAdder U29 (w399, IN30[0], IN30[1], w400, w401);
  FullAdder U30 (w401, IN31[0], IN31[1], w402, w403);
  FullAdder U31 (w403, IN32[0], IN32[1], w404, w405);
  FullAdder U32 (w405, IN33[0], IN33[1], w406, w407);
  FullAdder U33 (w407, IN34[0], IN34[1], w408, w409);
  FullAdder U34 (w409, IN35[0], IN35[1], w410, w411);
  FullAdder U35 (w411, IN36[0], IN36[1], w412, w413);
  FullAdder U36 (w413, IN37[0], IN37[1], w414, w415);
  FullAdder U37 (w415, IN38[0], IN38[1], w416, w417);
  FullAdder U38 (w417, IN39[0], IN39[1], w418, w419);
  FullAdder U39 (w419, IN40[0], IN40[1], w420, w421);
  FullAdder U40 (w421, IN41[0], IN41[1], w422, w423);
  FullAdder U41 (w423, IN42[0], IN42[1], w424, w425);
  FullAdder U42 (w425, IN43[0], IN43[1], w426, w427);
  FullAdder U43 (w427, IN44[0], IN44[1], w428, w429);
  FullAdder U44 (w429, IN45[0], IN45[1], w430, w431);
  FullAdder U45 (w431, IN46[0], IN46[1], w432, w433);
  FullAdder U46 (w433, IN47[0], IN47[1], w434, w435);
  FullAdder U47 (w435, IN48[0], IN48[1], w436, w437);
  FullAdder U48 (w437, IN49[0], IN49[1], w438, w439);
  FullAdder U49 (w439, IN50[0], IN50[1], w440, w441);
  FullAdder U50 (w441, IN51[0], IN51[1], w442, w443);
  FullAdder U51 (w443, IN52[0], IN52[1], w444, w445);
  FullAdder U52 (w445, IN53[0], IN53[1], w446, w447);
  FullAdder U53 (w447, IN54[0], IN54[1], w448, w449);
  FullAdder U54 (w449, IN55[0], IN55[1], w450, w451);
  FullAdder U55 (w451, IN56[0], IN56[1], w452, w453);
  HalfAdder U56 (w344, IN2[2], Out1[2], w455);
  FullAdder U57 (w455, w346, IN3[2], w456, w457);
  FullAdder U58 (w457, w348, IN4[2], w458, w459);
  FullAdder U59 (w459, w350, IN5[2], w460, w461);
  FullAdder U60 (w461, w352, IN6[2], w462, w463);
  FullAdder U61 (w463, w354, IN7[2], w464, w465);
  FullAdder U62 (w465, w356, IN8[2], w466, w467);
  FullAdder U63 (w467, w358, IN9[2], w468, w469);
  FullAdder U64 (w469, w360, IN10[2], w470, w471);
  FullAdder U65 (w471, w362, IN11[2], w472, w473);
  FullAdder U66 (w473, w364, IN12[2], w474, w475);
  FullAdder U67 (w475, w366, IN13[2], w476, w477);
  FullAdder U68 (w477, w368, IN14[2], w478, w479);
  FullAdder U69 (w479, w370, IN15[2], w480, w481);
  FullAdder U70 (w481, w372, IN16[2], w482, w483);
  FullAdder U71 (w483, w374, IN17[2], w484, w485);
  FullAdder U72 (w485, w376, IN18[2], w486, w487);
  FullAdder U73 (w487, w378, IN19[2], w488, w489);
  FullAdder U74 (w489, w380, IN20[2], w490, w491);
  FullAdder U75 (w491, w382, IN21[2], w492, w493);
  FullAdder U76 (w493, w384, IN22[2], w494, w495);
  FullAdder U77 (w495, w386, IN23[2], w496, w497);
  FullAdder U78 (w497, w388, IN24[2], w498, w499);
  FullAdder U79 (w499, w390, IN25[2], w500, w501);
  FullAdder U80 (w501, w392, IN26[2], w502, w503);
  FullAdder U81 (w503, w394, IN27[2], w504, w505);
  FullAdder U82 (w505, w396, IN28[2], w506, w507);
  FullAdder U83 (w507, w398, IN29[2], w508, w509);
  FullAdder U84 (w509, w400, IN30[2], w510, w511);
  FullAdder U85 (w511, w402, IN31[2], w512, w513);
  FullAdder U86 (w513, w404, IN32[2], w514, w515);
  FullAdder U87 (w515, w406, IN33[2], w516, w517);
  FullAdder U88 (w517, w408, IN34[2], w518, w519);
  FullAdder U89 (w519, w410, IN35[2], w520, w521);
  FullAdder U90 (w521, w412, IN36[2], w522, w523);
  FullAdder U91 (w523, w414, IN37[2], w524, w525);
  FullAdder U92 (w525, w416, IN38[2], w526, w527);
  FullAdder U93 (w527, w418, IN39[2], w528, w529);
  FullAdder U94 (w529, w420, IN40[2], w530, w531);
  FullAdder U95 (w531, w422, IN41[2], w532, w533);
  FullAdder U96 (w533, w424, IN42[2], w534, w535);
  FullAdder U97 (w535, w426, IN43[2], w536, w537);
  FullAdder U98 (w537, w428, IN44[2], w538, w539);
  FullAdder U99 (w539, w430, IN45[2], w540, w541);
  FullAdder U100 (w541, w432, IN46[2], w542, w543);
  FullAdder U101 (w543, w434, IN47[2], w544, w545);
  FullAdder U102 (w545, w436, IN48[2], w546, w547);
  FullAdder U103 (w547, w438, IN49[2], w548, w549);
  FullAdder U104 (w549, w440, IN50[2], w550, w551);
  FullAdder U105 (w551, w442, IN51[2], w552, w553);
  FullAdder U106 (w553, w444, IN52[2], w554, w555);
  FullAdder U107 (w555, w446, IN53[2], w556, w557);
  FullAdder U108 (w557, w448, IN54[2], w558, w559);
  FullAdder U109 (w559, w450, IN55[2], w560, w561);
  FullAdder U110 (w561, w452, IN56[2], w562, w563);
  FullAdder U111 (w563, w453, IN57[0], w564, w565);
  HalfAdder U112 (w456, IN3[3], Out1[3], w567);
  FullAdder U113 (w567, w458, IN4[3], w568, w569);
  FullAdder U114 (w569, w460, IN5[3], w570, w571);
  FullAdder U115 (w571, w462, IN6[3], w572, w573);
  FullAdder U116 (w573, w464, IN7[3], w574, w575);
  FullAdder U117 (w575, w466, IN8[3], w576, w577);
  FullAdder U118 (w577, w468, IN9[3], w578, w579);
  FullAdder U119 (w579, w470, IN10[3], w580, w581);
  FullAdder U120 (w581, w472, IN11[3], w582, w583);
  FullAdder U121 (w583, w474, IN12[3], w584, w585);
  FullAdder U122 (w585, w476, IN13[3], w586, w587);
  FullAdder U123 (w587, w478, IN14[3], w588, w589);
  FullAdder U124 (w589, w480, IN15[3], w590, w591);
  FullAdder U125 (w591, w482, IN16[3], w592, w593);
  FullAdder U126 (w593, w484, IN17[3], w594, w595);
  FullAdder U127 (w595, w486, IN18[3], w596, w597);
  FullAdder U128 (w597, w488, IN19[3], w598, w599);
  FullAdder U129 (w599, w490, IN20[3], w600, w601);
  FullAdder U130 (w601, w492, IN21[3], w602, w603);
  FullAdder U131 (w603, w494, IN22[3], w604, w605);
  FullAdder U132 (w605, w496, IN23[3], w606, w607);
  FullAdder U133 (w607, w498, IN24[3], w608, w609);
  FullAdder U134 (w609, w500, IN25[3], w610, w611);
  FullAdder U135 (w611, w502, IN26[3], w612, w613);
  FullAdder U136 (w613, w504, IN27[3], w614, w615);
  FullAdder U137 (w615, w506, IN28[3], w616, w617);
  FullAdder U138 (w617, w508, IN29[3], w618, w619);
  FullAdder U139 (w619, w510, IN30[3], w620, w621);
  FullAdder U140 (w621, w512, IN31[3], w622, w623);
  FullAdder U141 (w623, w514, IN32[3], w624, w625);
  FullAdder U142 (w625, w516, IN33[3], w626, w627);
  FullAdder U143 (w627, w518, IN34[3], w628, w629);
  FullAdder U144 (w629, w520, IN35[3], w630, w631);
  FullAdder U145 (w631, w522, IN36[3], w632, w633);
  FullAdder U146 (w633, w524, IN37[3], w634, w635);
  FullAdder U147 (w635, w526, IN38[3], w636, w637);
  FullAdder U148 (w637, w528, IN39[3], w638, w639);
  FullAdder U149 (w639, w530, IN40[3], w640, w641);
  FullAdder U150 (w641, w532, IN41[3], w642, w643);
  FullAdder U151 (w643, w534, IN42[3], w644, w645);
  FullAdder U152 (w645, w536, IN43[3], w646, w647);
  FullAdder U153 (w647, w538, IN44[3], w648, w649);
  FullAdder U154 (w649, w540, IN45[3], w650, w651);
  FullAdder U155 (w651, w542, IN46[3], w652, w653);
  FullAdder U156 (w653, w544, IN47[3], w654, w655);
  FullAdder U157 (w655, w546, IN48[3], w656, w657);
  FullAdder U158 (w657, w548, IN49[3], w658, w659);
  FullAdder U159 (w659, w550, IN50[3], w660, w661);
  FullAdder U160 (w661, w552, IN51[3], w662, w663);
  FullAdder U161 (w663, w554, IN52[3], w664, w665);
  FullAdder U162 (w665, w556, IN53[3], w666, w667);
  FullAdder U163 (w667, w558, IN54[3], w668, w669);
  FullAdder U164 (w669, w560, IN55[3], w670, w671);
  FullAdder U165 (w671, w562, IN56[3], w672, w673);
  FullAdder U166 (w673, w564, IN57[1], w674, w675);
  FullAdder U167 (w675, w565, IN58[0], w676, w677);
  HalfAdder U168 (w568, IN4[4], Out1[4], w679);
  FullAdder U169 (w679, w570, IN5[4], w680, w681);
  FullAdder U170 (w681, w572, IN6[4], w682, w683);
  FullAdder U171 (w683, w574, IN7[4], w684, w685);
  FullAdder U172 (w685, w576, IN8[4], w686, w687);
  FullAdder U173 (w687, w578, IN9[4], w688, w689);
  FullAdder U174 (w689, w580, IN10[4], w690, w691);
  FullAdder U175 (w691, w582, IN11[4], w692, w693);
  FullAdder U176 (w693, w584, IN12[4], w694, w695);
  FullAdder U177 (w695, w586, IN13[4], w696, w697);
  FullAdder U178 (w697, w588, IN14[4], w698, w699);
  FullAdder U179 (w699, w590, IN15[4], w700, w701);
  FullAdder U180 (w701, w592, IN16[4], w702, w703);
  FullAdder U181 (w703, w594, IN17[4], w704, w705);
  FullAdder U182 (w705, w596, IN18[4], w706, w707);
  FullAdder U183 (w707, w598, IN19[4], w708, w709);
  FullAdder U184 (w709, w600, IN20[4], w710, w711);
  FullAdder U185 (w711, w602, IN21[4], w712, w713);
  FullAdder U186 (w713, w604, IN22[4], w714, w715);
  FullAdder U187 (w715, w606, IN23[4], w716, w717);
  FullAdder U188 (w717, w608, IN24[4], w718, w719);
  FullAdder U189 (w719, w610, IN25[4], w720, w721);
  FullAdder U190 (w721, w612, IN26[4], w722, w723);
  FullAdder U191 (w723, w614, IN27[4], w724, w725);
  FullAdder U192 (w725, w616, IN28[4], w726, w727);
  FullAdder U193 (w727, w618, IN29[4], w728, w729);
  FullAdder U194 (w729, w620, IN30[4], w730, w731);
  FullAdder U195 (w731, w622, IN31[4], w732, w733);
  FullAdder U196 (w733, w624, IN32[4], w734, w735);
  FullAdder U197 (w735, w626, IN33[4], w736, w737);
  FullAdder U198 (w737, w628, IN34[4], w738, w739);
  FullAdder U199 (w739, w630, IN35[4], w740, w741);
  FullAdder U200 (w741, w632, IN36[4], w742, w743);
  FullAdder U201 (w743, w634, IN37[4], w744, w745);
  FullAdder U202 (w745, w636, IN38[4], w746, w747);
  FullAdder U203 (w747, w638, IN39[4], w748, w749);
  FullAdder U204 (w749, w640, IN40[4], w750, w751);
  FullAdder U205 (w751, w642, IN41[4], w752, w753);
  FullAdder U206 (w753, w644, IN42[4], w754, w755);
  FullAdder U207 (w755, w646, IN43[4], w756, w757);
  FullAdder U208 (w757, w648, IN44[4], w758, w759);
  FullAdder U209 (w759, w650, IN45[4], w760, w761);
  FullAdder U210 (w761, w652, IN46[4], w762, w763);
  FullAdder U211 (w763, w654, IN47[4], w764, w765);
  FullAdder U212 (w765, w656, IN48[4], w766, w767);
  FullAdder U213 (w767, w658, IN49[4], w768, w769);
  FullAdder U214 (w769, w660, IN50[4], w770, w771);
  FullAdder U215 (w771, w662, IN51[4], w772, w773);
  FullAdder U216 (w773, w664, IN52[4], w774, w775);
  FullAdder U217 (w775, w666, IN53[4], w776, w777);
  FullAdder U218 (w777, w668, IN54[4], w778, w779);
  FullAdder U219 (w779, w670, IN55[4], w780, w781);
  FullAdder U220 (w781, w672, IN56[4], w782, w783);
  FullAdder U221 (w783, w674, IN57[2], w784, w785);
  FullAdder U222 (w785, w676, IN58[1], w786, w787);
  FullAdder U223 (w787, w677, IN59[0], w788, w789);
  HalfAdder U224 (w680, IN5[5], Out1[5], w791);
  FullAdder U225 (w791, w682, IN6[5], Out1[6], w793);
  FullAdder U226 (w793, w684, IN7[5], Out1[7], w795);
  FullAdder U227 (w795, w686, IN8[5], Out1[8], w797);
  FullAdder U228 (w797, w688, IN9[5], Out1[9], w799);
  FullAdder U229 (w799, w690, IN10[5], Out1[10], w801);
  FullAdder U230 (w801, w692, IN11[5], Out1[11], w803);
  FullAdder U231 (w803, w694, IN12[5], Out1[12], w805);
  FullAdder U232 (w805, w696, IN13[5], Out1[13], w807);
  FullAdder U233 (w807, w698, IN14[5], Out1[14], w809);
  FullAdder U234 (w809, w700, IN15[5], Out1[15], w811);
  FullAdder U235 (w811, w702, IN16[5], Out1[16], w813);
  FullAdder U236 (w813, w704, IN17[5], Out1[17], w815);
  FullAdder U237 (w815, w706, IN18[5], Out1[18], w817);
  FullAdder U238 (w817, w708, IN19[5], Out1[19], w819);
  FullAdder U239 (w819, w710, IN20[5], Out1[20], w821);
  FullAdder U240 (w821, w712, IN21[5], Out1[21], w823);
  FullAdder U241 (w823, w714, IN22[5], Out1[22], w825);
  FullAdder U242 (w825, w716, IN23[5], Out1[23], w827);
  FullAdder U243 (w827, w718, IN24[5], Out1[24], w829);
  FullAdder U244 (w829, w720, IN25[5], Out1[25], w831);
  FullAdder U245 (w831, w722, IN26[5], Out1[26], w833);
  FullAdder U246 (w833, w724, IN27[5], Out1[27], w835);
  FullAdder U247 (w835, w726, IN28[5], Out1[28], w837);
  FullAdder U248 (w837, w728, IN29[5], Out1[29], w839);
  FullAdder U249 (w839, w730, IN30[5], Out1[30], w841);
  FullAdder U250 (w841, w732, IN31[5], Out1[31], w843);
  FullAdder U251 (w843, w734, IN32[5], Out1[32], w845);
  FullAdder U252 (w845, w736, IN33[5], Out1[33], w847);
  FullAdder U253 (w847, w738, IN34[5], Out1[34], w849);
  FullAdder U254 (w849, w740, IN35[5], Out1[35], w851);
  FullAdder U255 (w851, w742, IN36[5], Out1[36], w853);
  FullAdder U256 (w853, w744, IN37[5], Out1[37], w855);
  FullAdder U257 (w855, w746, IN38[5], Out1[38], w857);
  FullAdder U258 (w857, w748, IN39[5], Out1[39], w859);
  FullAdder U259 (w859, w750, IN40[5], Out1[40], w861);
  FullAdder U260 (w861, w752, IN41[5], Out1[41], w863);
  FullAdder U261 (w863, w754, IN42[5], Out1[42], w865);
  FullAdder U262 (w865, w756, IN43[5], Out1[43], w867);
  FullAdder U263 (w867, w758, IN44[5], Out1[44], w869);
  FullAdder U264 (w869, w760, IN45[5], Out1[45], w871);
  FullAdder U265 (w871, w762, IN46[5], Out1[46], w873);
  FullAdder U266 (w873, w764, IN47[5], Out1[47], w875);
  FullAdder U267 (w875, w766, IN48[5], Out1[48], w877);
  FullAdder U268 (w877, w768, IN49[5], Out1[49], w879);
  FullAdder U269 (w879, w770, IN50[5], Out1[50], w881);
  FullAdder U270 (w881, w772, IN51[5], Out1[51], w883);
  FullAdder U271 (w883, w774, IN52[5], Out1[52], w885);
  FullAdder U272 (w885, w776, IN53[5], Out1[53], w887);
  FullAdder U273 (w887, w778, IN54[5], Out1[54], w889);
  FullAdder U274 (w889, w780, IN55[5], Out1[55], w891);
  FullAdder U275 (w891, w782, IN56[5], Out1[56], w893);
  FullAdder U276 (w893, w784, IN57[3], Out1[57], w895);
  FullAdder U277 (w895, w786, IN58[2], Out1[58], w897);
  FullAdder U278 (w897, w788, IN59[1], Out1[59], w899);
  FullAdder U279 (w899, w789, IN60[0], Out1[60], Out1[61]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN57[4];
  assign Out2[1] = IN58[3];
  assign Out2[2] = IN59[2];
  assign Out2[3] = IN60[1];
  assign Out2[4] = IN61[0];

endmodule
module RC_5_5(IN1, IN2, Out);
  input [4:0] IN1;
  input [4:0] IN2;
  output [5:0] Out;
  wire w11;
  wire w13;
  wire w15;
  wire w17;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w11);
  FullAdder U1 (IN1[1], IN2[1], w11, Out[1], w13);
  FullAdder U2 (IN1[2], IN2[2], w13, Out[2], w15);
  FullAdder U3 (IN1[3], IN2[3], w15, Out[3], w17);
  FullAdder U4 (IN1[4], IN2[4], w17, Out[4], Out[5]);

endmodule
module NR_57_6(IN1, IN2, Out);
  input [56:0] IN1;
  input [5:0] IN2;
  output [62:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [5:0] P6;
  wire [5:0] P7;
  wire [5:0] P8;
  wire [5:0] P9;
  wire [5:0] P10;
  wire [5:0] P11;
  wire [5:0] P12;
  wire [5:0] P13;
  wire [5:0] P14;
  wire [5:0] P15;
  wire [5:0] P16;
  wire [5:0] P17;
  wire [5:0] P18;
  wire [5:0] P19;
  wire [5:0] P20;
  wire [5:0] P21;
  wire [5:0] P22;
  wire [5:0] P23;
  wire [5:0] P24;
  wire [5:0] P25;
  wire [5:0] P26;
  wire [5:0] P27;
  wire [5:0] P28;
  wire [5:0] P29;
  wire [5:0] P30;
  wire [5:0] P31;
  wire [5:0] P32;
  wire [5:0] P33;
  wire [5:0] P34;
  wire [5:0] P35;
  wire [5:0] P36;
  wire [5:0] P37;
  wire [5:0] P38;
  wire [5:0] P39;
  wire [5:0] P40;
  wire [5:0] P41;
  wire [5:0] P42;
  wire [5:0] P43;
  wire [5:0] P44;
  wire [5:0] P45;
  wire [5:0] P46;
  wire [5:0] P47;
  wire [5:0] P48;
  wire [5:0] P49;
  wire [5:0] P50;
  wire [5:0] P51;
  wire [5:0] P52;
  wire [5:0] P53;
  wire [5:0] P54;
  wire [5:0] P55;
  wire [5:0] P56;
  wire [4:0] P57;
  wire [3:0] P58;
  wire [2:0] P59;
  wire [1:0] P60;
  wire [0:0] P61;
  wire [61:0] R1;
  wire [4:0] R2;
  wire [62:0] aOut;
  U_SP_57_6 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, R1, R2);
  RC_5_5 S2 (R1[61:57], R2, aOut[62:57]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign Out = aOut[62:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
