
module NR_1_57(
    input [0:0]IN1,
    input [56:0]IN2,
    output [56:0]Out
);
    assign Out = IN2;
endmodule
