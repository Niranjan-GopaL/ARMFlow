
module NR_1_55(
    input [0:0]IN1,
    input [54:0]IN2,
    output [54:0]Out
);
    assign Out = IN2;
endmodule
