
module customAdder41_0(
    input [40 : 0] A,
    input [40 : 0] B,
    output [41 : 0] Sum
);

    assign Sum = A+B;

endmodule
