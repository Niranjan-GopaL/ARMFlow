//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 61
  second input length: 7
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_61_7(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66);
  input [60:0] IN1;
  input [6:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [6:0] P37;
  output [6:0] P38;
  output [6:0] P39;
  output [6:0] P40;
  output [6:0] P41;
  output [6:0] P42;
  output [6:0] P43;
  output [6:0] P44;
  output [6:0] P45;
  output [6:0] P46;
  output [6:0] P47;
  output [6:0] P48;
  output [6:0] P49;
  output [6:0] P50;
  output [6:0] P51;
  output [6:0] P52;
  output [6:0] P53;
  output [6:0] P54;
  output [6:0] P55;
  output [6:0] P56;
  output [6:0] P57;
  output [6:0] P58;
  output [6:0] P59;
  output [6:0] P60;
  output [5:0] P61;
  output [4:0] P62;
  output [3:0] P63;
  output [2:0] P64;
  output [1:0] P65;
  output [0:0] P66;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[0] = IN1[1]&IN2[6];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[1] = IN1[2]&IN2[5];
  assign P8[0] = IN1[2]&IN2[6];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[2] = IN1[3]&IN2[4];
  assign P8[1] = IN1[3]&IN2[5];
  assign P9[0] = IN1[3]&IN2[6];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[3] = IN1[4]&IN2[3];
  assign P8[2] = IN1[4]&IN2[4];
  assign P9[1] = IN1[4]&IN2[5];
  assign P10[0] = IN1[4]&IN2[6];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[4] = IN1[5]&IN2[2];
  assign P8[3] = IN1[5]&IN2[3];
  assign P9[2] = IN1[5]&IN2[4];
  assign P10[1] = IN1[5]&IN2[5];
  assign P11[0] = IN1[5]&IN2[6];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[5] = IN1[6]&IN2[1];
  assign P8[4] = IN1[6]&IN2[2];
  assign P9[3] = IN1[6]&IN2[3];
  assign P10[2] = IN1[6]&IN2[4];
  assign P11[1] = IN1[6]&IN2[5];
  assign P12[0] = IN1[6]&IN2[6];
  assign P7[6] = IN1[7]&IN2[0];
  assign P8[5] = IN1[7]&IN2[1];
  assign P9[4] = IN1[7]&IN2[2];
  assign P10[3] = IN1[7]&IN2[3];
  assign P11[2] = IN1[7]&IN2[4];
  assign P12[1] = IN1[7]&IN2[5];
  assign P13[0] = IN1[7]&IN2[6];
  assign P8[6] = IN1[8]&IN2[0];
  assign P9[5] = IN1[8]&IN2[1];
  assign P10[4] = IN1[8]&IN2[2];
  assign P11[3] = IN1[8]&IN2[3];
  assign P12[2] = IN1[8]&IN2[4];
  assign P13[1] = IN1[8]&IN2[5];
  assign P14[0] = IN1[8]&IN2[6];
  assign P9[6] = IN1[9]&IN2[0];
  assign P10[5] = IN1[9]&IN2[1];
  assign P11[4] = IN1[9]&IN2[2];
  assign P12[3] = IN1[9]&IN2[3];
  assign P13[2] = IN1[9]&IN2[4];
  assign P14[1] = IN1[9]&IN2[5];
  assign P15[0] = IN1[9]&IN2[6];
  assign P10[6] = IN1[10]&IN2[0];
  assign P11[5] = IN1[10]&IN2[1];
  assign P12[4] = IN1[10]&IN2[2];
  assign P13[3] = IN1[10]&IN2[3];
  assign P14[2] = IN1[10]&IN2[4];
  assign P15[1] = IN1[10]&IN2[5];
  assign P16[0] = IN1[10]&IN2[6];
  assign P11[6] = IN1[11]&IN2[0];
  assign P12[5] = IN1[11]&IN2[1];
  assign P13[4] = IN1[11]&IN2[2];
  assign P14[3] = IN1[11]&IN2[3];
  assign P15[2] = IN1[11]&IN2[4];
  assign P16[1] = IN1[11]&IN2[5];
  assign P17[0] = IN1[11]&IN2[6];
  assign P12[6] = IN1[12]&IN2[0];
  assign P13[5] = IN1[12]&IN2[1];
  assign P14[4] = IN1[12]&IN2[2];
  assign P15[3] = IN1[12]&IN2[3];
  assign P16[2] = IN1[12]&IN2[4];
  assign P17[1] = IN1[12]&IN2[5];
  assign P18[0] = IN1[12]&IN2[6];
  assign P13[6] = IN1[13]&IN2[0];
  assign P14[5] = IN1[13]&IN2[1];
  assign P15[4] = IN1[13]&IN2[2];
  assign P16[3] = IN1[13]&IN2[3];
  assign P17[2] = IN1[13]&IN2[4];
  assign P18[1] = IN1[13]&IN2[5];
  assign P19[0] = IN1[13]&IN2[6];
  assign P14[6] = IN1[14]&IN2[0];
  assign P15[5] = IN1[14]&IN2[1];
  assign P16[4] = IN1[14]&IN2[2];
  assign P17[3] = IN1[14]&IN2[3];
  assign P18[2] = IN1[14]&IN2[4];
  assign P19[1] = IN1[14]&IN2[5];
  assign P20[0] = IN1[14]&IN2[6];
  assign P15[6] = IN1[15]&IN2[0];
  assign P16[5] = IN1[15]&IN2[1];
  assign P17[4] = IN1[15]&IN2[2];
  assign P18[3] = IN1[15]&IN2[3];
  assign P19[2] = IN1[15]&IN2[4];
  assign P20[1] = IN1[15]&IN2[5];
  assign P21[0] = IN1[15]&IN2[6];
  assign P16[6] = IN1[16]&IN2[0];
  assign P17[5] = IN1[16]&IN2[1];
  assign P18[4] = IN1[16]&IN2[2];
  assign P19[3] = IN1[16]&IN2[3];
  assign P20[2] = IN1[16]&IN2[4];
  assign P21[1] = IN1[16]&IN2[5];
  assign P22[0] = IN1[16]&IN2[6];
  assign P17[6] = IN1[17]&IN2[0];
  assign P18[5] = IN1[17]&IN2[1];
  assign P19[4] = IN1[17]&IN2[2];
  assign P20[3] = IN1[17]&IN2[3];
  assign P21[2] = IN1[17]&IN2[4];
  assign P22[1] = IN1[17]&IN2[5];
  assign P23[0] = IN1[17]&IN2[6];
  assign P18[6] = IN1[18]&IN2[0];
  assign P19[5] = IN1[18]&IN2[1];
  assign P20[4] = IN1[18]&IN2[2];
  assign P21[3] = IN1[18]&IN2[3];
  assign P22[2] = IN1[18]&IN2[4];
  assign P23[1] = IN1[18]&IN2[5];
  assign P24[0] = IN1[18]&IN2[6];
  assign P19[6] = IN1[19]&IN2[0];
  assign P20[5] = IN1[19]&IN2[1];
  assign P21[4] = IN1[19]&IN2[2];
  assign P22[3] = IN1[19]&IN2[3];
  assign P23[2] = IN1[19]&IN2[4];
  assign P24[1] = IN1[19]&IN2[5];
  assign P25[0] = IN1[19]&IN2[6];
  assign P20[6] = IN1[20]&IN2[0];
  assign P21[5] = IN1[20]&IN2[1];
  assign P22[4] = IN1[20]&IN2[2];
  assign P23[3] = IN1[20]&IN2[3];
  assign P24[2] = IN1[20]&IN2[4];
  assign P25[1] = IN1[20]&IN2[5];
  assign P26[0] = IN1[20]&IN2[6];
  assign P21[6] = IN1[21]&IN2[0];
  assign P22[5] = IN1[21]&IN2[1];
  assign P23[4] = IN1[21]&IN2[2];
  assign P24[3] = IN1[21]&IN2[3];
  assign P25[2] = IN1[21]&IN2[4];
  assign P26[1] = IN1[21]&IN2[5];
  assign P27[0] = IN1[21]&IN2[6];
  assign P22[6] = IN1[22]&IN2[0];
  assign P23[5] = IN1[22]&IN2[1];
  assign P24[4] = IN1[22]&IN2[2];
  assign P25[3] = IN1[22]&IN2[3];
  assign P26[2] = IN1[22]&IN2[4];
  assign P27[1] = IN1[22]&IN2[5];
  assign P28[0] = IN1[22]&IN2[6];
  assign P23[6] = IN1[23]&IN2[0];
  assign P24[5] = IN1[23]&IN2[1];
  assign P25[4] = IN1[23]&IN2[2];
  assign P26[3] = IN1[23]&IN2[3];
  assign P27[2] = IN1[23]&IN2[4];
  assign P28[1] = IN1[23]&IN2[5];
  assign P29[0] = IN1[23]&IN2[6];
  assign P24[6] = IN1[24]&IN2[0];
  assign P25[5] = IN1[24]&IN2[1];
  assign P26[4] = IN1[24]&IN2[2];
  assign P27[3] = IN1[24]&IN2[3];
  assign P28[2] = IN1[24]&IN2[4];
  assign P29[1] = IN1[24]&IN2[5];
  assign P30[0] = IN1[24]&IN2[6];
  assign P25[6] = IN1[25]&IN2[0];
  assign P26[5] = IN1[25]&IN2[1];
  assign P27[4] = IN1[25]&IN2[2];
  assign P28[3] = IN1[25]&IN2[3];
  assign P29[2] = IN1[25]&IN2[4];
  assign P30[1] = IN1[25]&IN2[5];
  assign P31[0] = IN1[25]&IN2[6];
  assign P26[6] = IN1[26]&IN2[0];
  assign P27[5] = IN1[26]&IN2[1];
  assign P28[4] = IN1[26]&IN2[2];
  assign P29[3] = IN1[26]&IN2[3];
  assign P30[2] = IN1[26]&IN2[4];
  assign P31[1] = IN1[26]&IN2[5];
  assign P32[0] = IN1[26]&IN2[6];
  assign P27[6] = IN1[27]&IN2[0];
  assign P28[5] = IN1[27]&IN2[1];
  assign P29[4] = IN1[27]&IN2[2];
  assign P30[3] = IN1[27]&IN2[3];
  assign P31[2] = IN1[27]&IN2[4];
  assign P32[1] = IN1[27]&IN2[5];
  assign P33[0] = IN1[27]&IN2[6];
  assign P28[6] = IN1[28]&IN2[0];
  assign P29[5] = IN1[28]&IN2[1];
  assign P30[4] = IN1[28]&IN2[2];
  assign P31[3] = IN1[28]&IN2[3];
  assign P32[2] = IN1[28]&IN2[4];
  assign P33[1] = IN1[28]&IN2[5];
  assign P34[0] = IN1[28]&IN2[6];
  assign P29[6] = IN1[29]&IN2[0];
  assign P30[5] = IN1[29]&IN2[1];
  assign P31[4] = IN1[29]&IN2[2];
  assign P32[3] = IN1[29]&IN2[3];
  assign P33[2] = IN1[29]&IN2[4];
  assign P34[1] = IN1[29]&IN2[5];
  assign P35[0] = IN1[29]&IN2[6];
  assign P30[6] = IN1[30]&IN2[0];
  assign P31[5] = IN1[30]&IN2[1];
  assign P32[4] = IN1[30]&IN2[2];
  assign P33[3] = IN1[30]&IN2[3];
  assign P34[2] = IN1[30]&IN2[4];
  assign P35[1] = IN1[30]&IN2[5];
  assign P36[0] = IN1[30]&IN2[6];
  assign P31[6] = IN1[31]&IN2[0];
  assign P32[5] = IN1[31]&IN2[1];
  assign P33[4] = IN1[31]&IN2[2];
  assign P34[3] = IN1[31]&IN2[3];
  assign P35[2] = IN1[31]&IN2[4];
  assign P36[1] = IN1[31]&IN2[5];
  assign P37[0] = IN1[31]&IN2[6];
  assign P32[6] = IN1[32]&IN2[0];
  assign P33[5] = IN1[32]&IN2[1];
  assign P34[4] = IN1[32]&IN2[2];
  assign P35[3] = IN1[32]&IN2[3];
  assign P36[2] = IN1[32]&IN2[4];
  assign P37[1] = IN1[32]&IN2[5];
  assign P38[0] = IN1[32]&IN2[6];
  assign P33[6] = IN1[33]&IN2[0];
  assign P34[5] = IN1[33]&IN2[1];
  assign P35[4] = IN1[33]&IN2[2];
  assign P36[3] = IN1[33]&IN2[3];
  assign P37[2] = IN1[33]&IN2[4];
  assign P38[1] = IN1[33]&IN2[5];
  assign P39[0] = IN1[33]&IN2[6];
  assign P34[6] = IN1[34]&IN2[0];
  assign P35[5] = IN1[34]&IN2[1];
  assign P36[4] = IN1[34]&IN2[2];
  assign P37[3] = IN1[34]&IN2[3];
  assign P38[2] = IN1[34]&IN2[4];
  assign P39[1] = IN1[34]&IN2[5];
  assign P40[0] = IN1[34]&IN2[6];
  assign P35[6] = IN1[35]&IN2[0];
  assign P36[5] = IN1[35]&IN2[1];
  assign P37[4] = IN1[35]&IN2[2];
  assign P38[3] = IN1[35]&IN2[3];
  assign P39[2] = IN1[35]&IN2[4];
  assign P40[1] = IN1[35]&IN2[5];
  assign P41[0] = IN1[35]&IN2[6];
  assign P36[6] = IN1[36]&IN2[0];
  assign P37[5] = IN1[36]&IN2[1];
  assign P38[4] = IN1[36]&IN2[2];
  assign P39[3] = IN1[36]&IN2[3];
  assign P40[2] = IN1[36]&IN2[4];
  assign P41[1] = IN1[36]&IN2[5];
  assign P42[0] = IN1[36]&IN2[6];
  assign P37[6] = IN1[37]&IN2[0];
  assign P38[5] = IN1[37]&IN2[1];
  assign P39[4] = IN1[37]&IN2[2];
  assign P40[3] = IN1[37]&IN2[3];
  assign P41[2] = IN1[37]&IN2[4];
  assign P42[1] = IN1[37]&IN2[5];
  assign P43[0] = IN1[37]&IN2[6];
  assign P38[6] = IN1[38]&IN2[0];
  assign P39[5] = IN1[38]&IN2[1];
  assign P40[4] = IN1[38]&IN2[2];
  assign P41[3] = IN1[38]&IN2[3];
  assign P42[2] = IN1[38]&IN2[4];
  assign P43[1] = IN1[38]&IN2[5];
  assign P44[0] = IN1[38]&IN2[6];
  assign P39[6] = IN1[39]&IN2[0];
  assign P40[5] = IN1[39]&IN2[1];
  assign P41[4] = IN1[39]&IN2[2];
  assign P42[3] = IN1[39]&IN2[3];
  assign P43[2] = IN1[39]&IN2[4];
  assign P44[1] = IN1[39]&IN2[5];
  assign P45[0] = IN1[39]&IN2[6];
  assign P40[6] = IN1[40]&IN2[0];
  assign P41[5] = IN1[40]&IN2[1];
  assign P42[4] = IN1[40]&IN2[2];
  assign P43[3] = IN1[40]&IN2[3];
  assign P44[2] = IN1[40]&IN2[4];
  assign P45[1] = IN1[40]&IN2[5];
  assign P46[0] = IN1[40]&IN2[6];
  assign P41[6] = IN1[41]&IN2[0];
  assign P42[5] = IN1[41]&IN2[1];
  assign P43[4] = IN1[41]&IN2[2];
  assign P44[3] = IN1[41]&IN2[3];
  assign P45[2] = IN1[41]&IN2[4];
  assign P46[1] = IN1[41]&IN2[5];
  assign P47[0] = IN1[41]&IN2[6];
  assign P42[6] = IN1[42]&IN2[0];
  assign P43[5] = IN1[42]&IN2[1];
  assign P44[4] = IN1[42]&IN2[2];
  assign P45[3] = IN1[42]&IN2[3];
  assign P46[2] = IN1[42]&IN2[4];
  assign P47[1] = IN1[42]&IN2[5];
  assign P48[0] = IN1[42]&IN2[6];
  assign P43[6] = IN1[43]&IN2[0];
  assign P44[5] = IN1[43]&IN2[1];
  assign P45[4] = IN1[43]&IN2[2];
  assign P46[3] = IN1[43]&IN2[3];
  assign P47[2] = IN1[43]&IN2[4];
  assign P48[1] = IN1[43]&IN2[5];
  assign P49[0] = IN1[43]&IN2[6];
  assign P44[6] = IN1[44]&IN2[0];
  assign P45[5] = IN1[44]&IN2[1];
  assign P46[4] = IN1[44]&IN2[2];
  assign P47[3] = IN1[44]&IN2[3];
  assign P48[2] = IN1[44]&IN2[4];
  assign P49[1] = IN1[44]&IN2[5];
  assign P50[0] = IN1[44]&IN2[6];
  assign P45[6] = IN1[45]&IN2[0];
  assign P46[5] = IN1[45]&IN2[1];
  assign P47[4] = IN1[45]&IN2[2];
  assign P48[3] = IN1[45]&IN2[3];
  assign P49[2] = IN1[45]&IN2[4];
  assign P50[1] = IN1[45]&IN2[5];
  assign P51[0] = IN1[45]&IN2[6];
  assign P46[6] = IN1[46]&IN2[0];
  assign P47[5] = IN1[46]&IN2[1];
  assign P48[4] = IN1[46]&IN2[2];
  assign P49[3] = IN1[46]&IN2[3];
  assign P50[2] = IN1[46]&IN2[4];
  assign P51[1] = IN1[46]&IN2[5];
  assign P52[0] = IN1[46]&IN2[6];
  assign P47[6] = IN1[47]&IN2[0];
  assign P48[5] = IN1[47]&IN2[1];
  assign P49[4] = IN1[47]&IN2[2];
  assign P50[3] = IN1[47]&IN2[3];
  assign P51[2] = IN1[47]&IN2[4];
  assign P52[1] = IN1[47]&IN2[5];
  assign P53[0] = IN1[47]&IN2[6];
  assign P48[6] = IN1[48]&IN2[0];
  assign P49[5] = IN1[48]&IN2[1];
  assign P50[4] = IN1[48]&IN2[2];
  assign P51[3] = IN1[48]&IN2[3];
  assign P52[2] = IN1[48]&IN2[4];
  assign P53[1] = IN1[48]&IN2[5];
  assign P54[0] = IN1[48]&IN2[6];
  assign P49[6] = IN1[49]&IN2[0];
  assign P50[5] = IN1[49]&IN2[1];
  assign P51[4] = IN1[49]&IN2[2];
  assign P52[3] = IN1[49]&IN2[3];
  assign P53[2] = IN1[49]&IN2[4];
  assign P54[1] = IN1[49]&IN2[5];
  assign P55[0] = IN1[49]&IN2[6];
  assign P50[6] = IN1[50]&IN2[0];
  assign P51[5] = IN1[50]&IN2[1];
  assign P52[4] = IN1[50]&IN2[2];
  assign P53[3] = IN1[50]&IN2[3];
  assign P54[2] = IN1[50]&IN2[4];
  assign P55[1] = IN1[50]&IN2[5];
  assign P56[0] = IN1[50]&IN2[6];
  assign P51[6] = IN1[51]&IN2[0];
  assign P52[5] = IN1[51]&IN2[1];
  assign P53[4] = IN1[51]&IN2[2];
  assign P54[3] = IN1[51]&IN2[3];
  assign P55[2] = IN1[51]&IN2[4];
  assign P56[1] = IN1[51]&IN2[5];
  assign P57[0] = IN1[51]&IN2[6];
  assign P52[6] = IN1[52]&IN2[0];
  assign P53[5] = IN1[52]&IN2[1];
  assign P54[4] = IN1[52]&IN2[2];
  assign P55[3] = IN1[52]&IN2[3];
  assign P56[2] = IN1[52]&IN2[4];
  assign P57[1] = IN1[52]&IN2[5];
  assign P58[0] = IN1[52]&IN2[6];
  assign P53[6] = IN1[53]&IN2[0];
  assign P54[5] = IN1[53]&IN2[1];
  assign P55[4] = IN1[53]&IN2[2];
  assign P56[3] = IN1[53]&IN2[3];
  assign P57[2] = IN1[53]&IN2[4];
  assign P58[1] = IN1[53]&IN2[5];
  assign P59[0] = IN1[53]&IN2[6];
  assign P54[6] = IN1[54]&IN2[0];
  assign P55[5] = IN1[54]&IN2[1];
  assign P56[4] = IN1[54]&IN2[2];
  assign P57[3] = IN1[54]&IN2[3];
  assign P58[2] = IN1[54]&IN2[4];
  assign P59[1] = IN1[54]&IN2[5];
  assign P60[0] = IN1[54]&IN2[6];
  assign P55[6] = IN1[55]&IN2[0];
  assign P56[5] = IN1[55]&IN2[1];
  assign P57[4] = IN1[55]&IN2[2];
  assign P58[3] = IN1[55]&IN2[3];
  assign P59[2] = IN1[55]&IN2[4];
  assign P60[1] = IN1[55]&IN2[5];
  assign P61[0] = IN1[55]&IN2[6];
  assign P56[6] = IN1[56]&IN2[0];
  assign P57[5] = IN1[56]&IN2[1];
  assign P58[4] = IN1[56]&IN2[2];
  assign P59[3] = IN1[56]&IN2[3];
  assign P60[2] = IN1[56]&IN2[4];
  assign P61[1] = IN1[56]&IN2[5];
  assign P62[0] = IN1[56]&IN2[6];
  assign P57[6] = IN1[57]&IN2[0];
  assign P58[5] = IN1[57]&IN2[1];
  assign P59[4] = IN1[57]&IN2[2];
  assign P60[3] = IN1[57]&IN2[3];
  assign P61[2] = IN1[57]&IN2[4];
  assign P62[1] = IN1[57]&IN2[5];
  assign P63[0] = IN1[57]&IN2[6];
  assign P58[6] = IN1[58]&IN2[0];
  assign P59[5] = IN1[58]&IN2[1];
  assign P60[4] = IN1[58]&IN2[2];
  assign P61[3] = IN1[58]&IN2[3];
  assign P62[2] = IN1[58]&IN2[4];
  assign P63[1] = IN1[58]&IN2[5];
  assign P64[0] = IN1[58]&IN2[6];
  assign P59[6] = IN1[59]&IN2[0];
  assign P60[5] = IN1[59]&IN2[1];
  assign P61[4] = IN1[59]&IN2[2];
  assign P62[3] = IN1[59]&IN2[3];
  assign P63[2] = IN1[59]&IN2[4];
  assign P64[1] = IN1[59]&IN2[5];
  assign P65[0] = IN1[59]&IN2[6];
  assign P60[6] = IN1[60]&IN2[0];
  assign P61[5] = IN1[60]&IN2[1];
  assign P62[4] = IN1[60]&IN2[2];
  assign P63[3] = IN1[60]&IN2[3];
  assign P64[2] = IN1[60]&IN2[4];
  assign P65[1] = IN1[60]&IN2[5];
  assign P66[0] = IN1[60]&IN2[6];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [6:0] IN37;
  input [6:0] IN38;
  input [6:0] IN39;
  input [6:0] IN40;
  input [6:0] IN41;
  input [6:0] IN42;
  input [6:0] IN43;
  input [6:0] IN44;
  input [6:0] IN45;
  input [6:0] IN46;
  input [6:0] IN47;
  input [6:0] IN48;
  input [6:0] IN49;
  input [6:0] IN50;
  input [6:0] IN51;
  input [6:0] IN52;
  input [6:0] IN53;
  input [6:0] IN54;
  input [6:0] IN55;
  input [6:0] IN56;
  input [6:0] IN57;
  input [6:0] IN58;
  input [6:0] IN59;
  input [6:0] IN60;
  input [5:0] IN61;
  input [4:0] IN62;
  input [3:0] IN63;
  input [2:0] IN64;
  input [1:0] IN65;
  input [0:0] IN66;
  output [66:0] Out1;
  output [5:0] Out2;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1028;
  wire w1030;
  wire w1032;
  wire w1034;
  wire w1036;
  wire w1038;
  wire w1040;
  wire w1042;
  wire w1044;
  wire w1046;
  wire w1048;
  wire w1050;
  wire w1052;
  wire w1054;
  wire w1056;
  wire w1058;
  wire w1060;
  wire w1062;
  wire w1064;
  wire w1066;
  wire w1068;
  wire w1070;
  wire w1072;
  wire w1074;
  wire w1076;
  wire w1078;
  wire w1080;
  wire w1082;
  wire w1084;
  wire w1086;
  wire w1088;
  wire w1090;
  wire w1092;
  wire w1094;
  wire w1096;
  wire w1098;
  wire w1100;
  wire w1102;
  wire w1104;
  wire w1106;
  wire w1108;
  wire w1110;
  wire w1112;
  wire w1114;
  wire w1116;
  wire w1118;
  wire w1120;
  wire w1122;
  wire w1124;
  wire w1126;
  wire w1128;
  wire w1130;
  wire w1132;
  wire w1134;
  wire w1136;
  wire w1138;
  wire w1140;
  wire w1142;
  wire w1144;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w428);
  FullAdder U1 (w428, IN2[0], IN2[1], w429, w430);
  FullAdder U2 (w430, IN3[0], IN3[1], w431, w432);
  FullAdder U3 (w432, IN4[0], IN4[1], w433, w434);
  FullAdder U4 (w434, IN5[0], IN5[1], w435, w436);
  FullAdder U5 (w436, IN6[0], IN6[1], w437, w438);
  FullAdder U6 (w438, IN7[0], IN7[1], w439, w440);
  FullAdder U7 (w440, IN8[0], IN8[1], w441, w442);
  FullAdder U8 (w442, IN9[0], IN9[1], w443, w444);
  FullAdder U9 (w444, IN10[0], IN10[1], w445, w446);
  FullAdder U10 (w446, IN11[0], IN11[1], w447, w448);
  FullAdder U11 (w448, IN12[0], IN12[1], w449, w450);
  FullAdder U12 (w450, IN13[0], IN13[1], w451, w452);
  FullAdder U13 (w452, IN14[0], IN14[1], w453, w454);
  FullAdder U14 (w454, IN15[0], IN15[1], w455, w456);
  FullAdder U15 (w456, IN16[0], IN16[1], w457, w458);
  FullAdder U16 (w458, IN17[0], IN17[1], w459, w460);
  FullAdder U17 (w460, IN18[0], IN18[1], w461, w462);
  FullAdder U18 (w462, IN19[0], IN19[1], w463, w464);
  FullAdder U19 (w464, IN20[0], IN20[1], w465, w466);
  FullAdder U20 (w466, IN21[0], IN21[1], w467, w468);
  FullAdder U21 (w468, IN22[0], IN22[1], w469, w470);
  FullAdder U22 (w470, IN23[0], IN23[1], w471, w472);
  FullAdder U23 (w472, IN24[0], IN24[1], w473, w474);
  FullAdder U24 (w474, IN25[0], IN25[1], w475, w476);
  FullAdder U25 (w476, IN26[0], IN26[1], w477, w478);
  FullAdder U26 (w478, IN27[0], IN27[1], w479, w480);
  FullAdder U27 (w480, IN28[0], IN28[1], w481, w482);
  FullAdder U28 (w482, IN29[0], IN29[1], w483, w484);
  FullAdder U29 (w484, IN30[0], IN30[1], w485, w486);
  FullAdder U30 (w486, IN31[0], IN31[1], w487, w488);
  FullAdder U31 (w488, IN32[0], IN32[1], w489, w490);
  FullAdder U32 (w490, IN33[0], IN33[1], w491, w492);
  FullAdder U33 (w492, IN34[0], IN34[1], w493, w494);
  FullAdder U34 (w494, IN35[0], IN35[1], w495, w496);
  FullAdder U35 (w496, IN36[0], IN36[1], w497, w498);
  FullAdder U36 (w498, IN37[0], IN37[1], w499, w500);
  FullAdder U37 (w500, IN38[0], IN38[1], w501, w502);
  FullAdder U38 (w502, IN39[0], IN39[1], w503, w504);
  FullAdder U39 (w504, IN40[0], IN40[1], w505, w506);
  FullAdder U40 (w506, IN41[0], IN41[1], w507, w508);
  FullAdder U41 (w508, IN42[0], IN42[1], w509, w510);
  FullAdder U42 (w510, IN43[0], IN43[1], w511, w512);
  FullAdder U43 (w512, IN44[0], IN44[1], w513, w514);
  FullAdder U44 (w514, IN45[0], IN45[1], w515, w516);
  FullAdder U45 (w516, IN46[0], IN46[1], w517, w518);
  FullAdder U46 (w518, IN47[0], IN47[1], w519, w520);
  FullAdder U47 (w520, IN48[0], IN48[1], w521, w522);
  FullAdder U48 (w522, IN49[0], IN49[1], w523, w524);
  FullAdder U49 (w524, IN50[0], IN50[1], w525, w526);
  FullAdder U50 (w526, IN51[0], IN51[1], w527, w528);
  FullAdder U51 (w528, IN52[0], IN52[1], w529, w530);
  FullAdder U52 (w530, IN53[0], IN53[1], w531, w532);
  FullAdder U53 (w532, IN54[0], IN54[1], w533, w534);
  FullAdder U54 (w534, IN55[0], IN55[1], w535, w536);
  FullAdder U55 (w536, IN56[0], IN56[1], w537, w538);
  FullAdder U56 (w538, IN57[0], IN57[1], w539, w540);
  FullAdder U57 (w540, IN58[0], IN58[1], w541, w542);
  FullAdder U58 (w542, IN59[0], IN59[1], w543, w544);
  FullAdder U59 (w544, IN60[0], IN60[1], w545, w546);
  HalfAdder U60 (w429, IN2[2], Out1[2], w548);
  FullAdder U61 (w548, w431, IN3[2], w549, w550);
  FullAdder U62 (w550, w433, IN4[2], w551, w552);
  FullAdder U63 (w552, w435, IN5[2], w553, w554);
  FullAdder U64 (w554, w437, IN6[2], w555, w556);
  FullAdder U65 (w556, w439, IN7[2], w557, w558);
  FullAdder U66 (w558, w441, IN8[2], w559, w560);
  FullAdder U67 (w560, w443, IN9[2], w561, w562);
  FullAdder U68 (w562, w445, IN10[2], w563, w564);
  FullAdder U69 (w564, w447, IN11[2], w565, w566);
  FullAdder U70 (w566, w449, IN12[2], w567, w568);
  FullAdder U71 (w568, w451, IN13[2], w569, w570);
  FullAdder U72 (w570, w453, IN14[2], w571, w572);
  FullAdder U73 (w572, w455, IN15[2], w573, w574);
  FullAdder U74 (w574, w457, IN16[2], w575, w576);
  FullAdder U75 (w576, w459, IN17[2], w577, w578);
  FullAdder U76 (w578, w461, IN18[2], w579, w580);
  FullAdder U77 (w580, w463, IN19[2], w581, w582);
  FullAdder U78 (w582, w465, IN20[2], w583, w584);
  FullAdder U79 (w584, w467, IN21[2], w585, w586);
  FullAdder U80 (w586, w469, IN22[2], w587, w588);
  FullAdder U81 (w588, w471, IN23[2], w589, w590);
  FullAdder U82 (w590, w473, IN24[2], w591, w592);
  FullAdder U83 (w592, w475, IN25[2], w593, w594);
  FullAdder U84 (w594, w477, IN26[2], w595, w596);
  FullAdder U85 (w596, w479, IN27[2], w597, w598);
  FullAdder U86 (w598, w481, IN28[2], w599, w600);
  FullAdder U87 (w600, w483, IN29[2], w601, w602);
  FullAdder U88 (w602, w485, IN30[2], w603, w604);
  FullAdder U89 (w604, w487, IN31[2], w605, w606);
  FullAdder U90 (w606, w489, IN32[2], w607, w608);
  FullAdder U91 (w608, w491, IN33[2], w609, w610);
  FullAdder U92 (w610, w493, IN34[2], w611, w612);
  FullAdder U93 (w612, w495, IN35[2], w613, w614);
  FullAdder U94 (w614, w497, IN36[2], w615, w616);
  FullAdder U95 (w616, w499, IN37[2], w617, w618);
  FullAdder U96 (w618, w501, IN38[2], w619, w620);
  FullAdder U97 (w620, w503, IN39[2], w621, w622);
  FullAdder U98 (w622, w505, IN40[2], w623, w624);
  FullAdder U99 (w624, w507, IN41[2], w625, w626);
  FullAdder U100 (w626, w509, IN42[2], w627, w628);
  FullAdder U101 (w628, w511, IN43[2], w629, w630);
  FullAdder U102 (w630, w513, IN44[2], w631, w632);
  FullAdder U103 (w632, w515, IN45[2], w633, w634);
  FullAdder U104 (w634, w517, IN46[2], w635, w636);
  FullAdder U105 (w636, w519, IN47[2], w637, w638);
  FullAdder U106 (w638, w521, IN48[2], w639, w640);
  FullAdder U107 (w640, w523, IN49[2], w641, w642);
  FullAdder U108 (w642, w525, IN50[2], w643, w644);
  FullAdder U109 (w644, w527, IN51[2], w645, w646);
  FullAdder U110 (w646, w529, IN52[2], w647, w648);
  FullAdder U111 (w648, w531, IN53[2], w649, w650);
  FullAdder U112 (w650, w533, IN54[2], w651, w652);
  FullAdder U113 (w652, w535, IN55[2], w653, w654);
  FullAdder U114 (w654, w537, IN56[2], w655, w656);
  FullAdder U115 (w656, w539, IN57[2], w657, w658);
  FullAdder U116 (w658, w541, IN58[2], w659, w660);
  FullAdder U117 (w660, w543, IN59[2], w661, w662);
  FullAdder U118 (w662, w545, IN60[2], w663, w664);
  FullAdder U119 (w664, w546, IN61[0], w665, w666);
  HalfAdder U120 (w549, IN3[3], Out1[3], w668);
  FullAdder U121 (w668, w551, IN4[3], w669, w670);
  FullAdder U122 (w670, w553, IN5[3], w671, w672);
  FullAdder U123 (w672, w555, IN6[3], w673, w674);
  FullAdder U124 (w674, w557, IN7[3], w675, w676);
  FullAdder U125 (w676, w559, IN8[3], w677, w678);
  FullAdder U126 (w678, w561, IN9[3], w679, w680);
  FullAdder U127 (w680, w563, IN10[3], w681, w682);
  FullAdder U128 (w682, w565, IN11[3], w683, w684);
  FullAdder U129 (w684, w567, IN12[3], w685, w686);
  FullAdder U130 (w686, w569, IN13[3], w687, w688);
  FullAdder U131 (w688, w571, IN14[3], w689, w690);
  FullAdder U132 (w690, w573, IN15[3], w691, w692);
  FullAdder U133 (w692, w575, IN16[3], w693, w694);
  FullAdder U134 (w694, w577, IN17[3], w695, w696);
  FullAdder U135 (w696, w579, IN18[3], w697, w698);
  FullAdder U136 (w698, w581, IN19[3], w699, w700);
  FullAdder U137 (w700, w583, IN20[3], w701, w702);
  FullAdder U138 (w702, w585, IN21[3], w703, w704);
  FullAdder U139 (w704, w587, IN22[3], w705, w706);
  FullAdder U140 (w706, w589, IN23[3], w707, w708);
  FullAdder U141 (w708, w591, IN24[3], w709, w710);
  FullAdder U142 (w710, w593, IN25[3], w711, w712);
  FullAdder U143 (w712, w595, IN26[3], w713, w714);
  FullAdder U144 (w714, w597, IN27[3], w715, w716);
  FullAdder U145 (w716, w599, IN28[3], w717, w718);
  FullAdder U146 (w718, w601, IN29[3], w719, w720);
  FullAdder U147 (w720, w603, IN30[3], w721, w722);
  FullAdder U148 (w722, w605, IN31[3], w723, w724);
  FullAdder U149 (w724, w607, IN32[3], w725, w726);
  FullAdder U150 (w726, w609, IN33[3], w727, w728);
  FullAdder U151 (w728, w611, IN34[3], w729, w730);
  FullAdder U152 (w730, w613, IN35[3], w731, w732);
  FullAdder U153 (w732, w615, IN36[3], w733, w734);
  FullAdder U154 (w734, w617, IN37[3], w735, w736);
  FullAdder U155 (w736, w619, IN38[3], w737, w738);
  FullAdder U156 (w738, w621, IN39[3], w739, w740);
  FullAdder U157 (w740, w623, IN40[3], w741, w742);
  FullAdder U158 (w742, w625, IN41[3], w743, w744);
  FullAdder U159 (w744, w627, IN42[3], w745, w746);
  FullAdder U160 (w746, w629, IN43[3], w747, w748);
  FullAdder U161 (w748, w631, IN44[3], w749, w750);
  FullAdder U162 (w750, w633, IN45[3], w751, w752);
  FullAdder U163 (w752, w635, IN46[3], w753, w754);
  FullAdder U164 (w754, w637, IN47[3], w755, w756);
  FullAdder U165 (w756, w639, IN48[3], w757, w758);
  FullAdder U166 (w758, w641, IN49[3], w759, w760);
  FullAdder U167 (w760, w643, IN50[3], w761, w762);
  FullAdder U168 (w762, w645, IN51[3], w763, w764);
  FullAdder U169 (w764, w647, IN52[3], w765, w766);
  FullAdder U170 (w766, w649, IN53[3], w767, w768);
  FullAdder U171 (w768, w651, IN54[3], w769, w770);
  FullAdder U172 (w770, w653, IN55[3], w771, w772);
  FullAdder U173 (w772, w655, IN56[3], w773, w774);
  FullAdder U174 (w774, w657, IN57[3], w775, w776);
  FullAdder U175 (w776, w659, IN58[3], w777, w778);
  FullAdder U176 (w778, w661, IN59[3], w779, w780);
  FullAdder U177 (w780, w663, IN60[3], w781, w782);
  FullAdder U178 (w782, w665, IN61[1], w783, w784);
  FullAdder U179 (w784, w666, IN62[0], w785, w786);
  HalfAdder U180 (w669, IN4[4], Out1[4], w788);
  FullAdder U181 (w788, w671, IN5[4], w789, w790);
  FullAdder U182 (w790, w673, IN6[4], w791, w792);
  FullAdder U183 (w792, w675, IN7[4], w793, w794);
  FullAdder U184 (w794, w677, IN8[4], w795, w796);
  FullAdder U185 (w796, w679, IN9[4], w797, w798);
  FullAdder U186 (w798, w681, IN10[4], w799, w800);
  FullAdder U187 (w800, w683, IN11[4], w801, w802);
  FullAdder U188 (w802, w685, IN12[4], w803, w804);
  FullAdder U189 (w804, w687, IN13[4], w805, w806);
  FullAdder U190 (w806, w689, IN14[4], w807, w808);
  FullAdder U191 (w808, w691, IN15[4], w809, w810);
  FullAdder U192 (w810, w693, IN16[4], w811, w812);
  FullAdder U193 (w812, w695, IN17[4], w813, w814);
  FullAdder U194 (w814, w697, IN18[4], w815, w816);
  FullAdder U195 (w816, w699, IN19[4], w817, w818);
  FullAdder U196 (w818, w701, IN20[4], w819, w820);
  FullAdder U197 (w820, w703, IN21[4], w821, w822);
  FullAdder U198 (w822, w705, IN22[4], w823, w824);
  FullAdder U199 (w824, w707, IN23[4], w825, w826);
  FullAdder U200 (w826, w709, IN24[4], w827, w828);
  FullAdder U201 (w828, w711, IN25[4], w829, w830);
  FullAdder U202 (w830, w713, IN26[4], w831, w832);
  FullAdder U203 (w832, w715, IN27[4], w833, w834);
  FullAdder U204 (w834, w717, IN28[4], w835, w836);
  FullAdder U205 (w836, w719, IN29[4], w837, w838);
  FullAdder U206 (w838, w721, IN30[4], w839, w840);
  FullAdder U207 (w840, w723, IN31[4], w841, w842);
  FullAdder U208 (w842, w725, IN32[4], w843, w844);
  FullAdder U209 (w844, w727, IN33[4], w845, w846);
  FullAdder U210 (w846, w729, IN34[4], w847, w848);
  FullAdder U211 (w848, w731, IN35[4], w849, w850);
  FullAdder U212 (w850, w733, IN36[4], w851, w852);
  FullAdder U213 (w852, w735, IN37[4], w853, w854);
  FullAdder U214 (w854, w737, IN38[4], w855, w856);
  FullAdder U215 (w856, w739, IN39[4], w857, w858);
  FullAdder U216 (w858, w741, IN40[4], w859, w860);
  FullAdder U217 (w860, w743, IN41[4], w861, w862);
  FullAdder U218 (w862, w745, IN42[4], w863, w864);
  FullAdder U219 (w864, w747, IN43[4], w865, w866);
  FullAdder U220 (w866, w749, IN44[4], w867, w868);
  FullAdder U221 (w868, w751, IN45[4], w869, w870);
  FullAdder U222 (w870, w753, IN46[4], w871, w872);
  FullAdder U223 (w872, w755, IN47[4], w873, w874);
  FullAdder U224 (w874, w757, IN48[4], w875, w876);
  FullAdder U225 (w876, w759, IN49[4], w877, w878);
  FullAdder U226 (w878, w761, IN50[4], w879, w880);
  FullAdder U227 (w880, w763, IN51[4], w881, w882);
  FullAdder U228 (w882, w765, IN52[4], w883, w884);
  FullAdder U229 (w884, w767, IN53[4], w885, w886);
  FullAdder U230 (w886, w769, IN54[4], w887, w888);
  FullAdder U231 (w888, w771, IN55[4], w889, w890);
  FullAdder U232 (w890, w773, IN56[4], w891, w892);
  FullAdder U233 (w892, w775, IN57[4], w893, w894);
  FullAdder U234 (w894, w777, IN58[4], w895, w896);
  FullAdder U235 (w896, w779, IN59[4], w897, w898);
  FullAdder U236 (w898, w781, IN60[4], w899, w900);
  FullAdder U237 (w900, w783, IN61[2], w901, w902);
  FullAdder U238 (w902, w785, IN62[1], w903, w904);
  FullAdder U239 (w904, w786, IN63[0], w905, w906);
  HalfAdder U240 (w789, IN5[5], Out1[5], w908);
  FullAdder U241 (w908, w791, IN6[5], w909, w910);
  FullAdder U242 (w910, w793, IN7[5], w911, w912);
  FullAdder U243 (w912, w795, IN8[5], w913, w914);
  FullAdder U244 (w914, w797, IN9[5], w915, w916);
  FullAdder U245 (w916, w799, IN10[5], w917, w918);
  FullAdder U246 (w918, w801, IN11[5], w919, w920);
  FullAdder U247 (w920, w803, IN12[5], w921, w922);
  FullAdder U248 (w922, w805, IN13[5], w923, w924);
  FullAdder U249 (w924, w807, IN14[5], w925, w926);
  FullAdder U250 (w926, w809, IN15[5], w927, w928);
  FullAdder U251 (w928, w811, IN16[5], w929, w930);
  FullAdder U252 (w930, w813, IN17[5], w931, w932);
  FullAdder U253 (w932, w815, IN18[5], w933, w934);
  FullAdder U254 (w934, w817, IN19[5], w935, w936);
  FullAdder U255 (w936, w819, IN20[5], w937, w938);
  FullAdder U256 (w938, w821, IN21[5], w939, w940);
  FullAdder U257 (w940, w823, IN22[5], w941, w942);
  FullAdder U258 (w942, w825, IN23[5], w943, w944);
  FullAdder U259 (w944, w827, IN24[5], w945, w946);
  FullAdder U260 (w946, w829, IN25[5], w947, w948);
  FullAdder U261 (w948, w831, IN26[5], w949, w950);
  FullAdder U262 (w950, w833, IN27[5], w951, w952);
  FullAdder U263 (w952, w835, IN28[5], w953, w954);
  FullAdder U264 (w954, w837, IN29[5], w955, w956);
  FullAdder U265 (w956, w839, IN30[5], w957, w958);
  FullAdder U266 (w958, w841, IN31[5], w959, w960);
  FullAdder U267 (w960, w843, IN32[5], w961, w962);
  FullAdder U268 (w962, w845, IN33[5], w963, w964);
  FullAdder U269 (w964, w847, IN34[5], w965, w966);
  FullAdder U270 (w966, w849, IN35[5], w967, w968);
  FullAdder U271 (w968, w851, IN36[5], w969, w970);
  FullAdder U272 (w970, w853, IN37[5], w971, w972);
  FullAdder U273 (w972, w855, IN38[5], w973, w974);
  FullAdder U274 (w974, w857, IN39[5], w975, w976);
  FullAdder U275 (w976, w859, IN40[5], w977, w978);
  FullAdder U276 (w978, w861, IN41[5], w979, w980);
  FullAdder U277 (w980, w863, IN42[5], w981, w982);
  FullAdder U278 (w982, w865, IN43[5], w983, w984);
  FullAdder U279 (w984, w867, IN44[5], w985, w986);
  FullAdder U280 (w986, w869, IN45[5], w987, w988);
  FullAdder U281 (w988, w871, IN46[5], w989, w990);
  FullAdder U282 (w990, w873, IN47[5], w991, w992);
  FullAdder U283 (w992, w875, IN48[5], w993, w994);
  FullAdder U284 (w994, w877, IN49[5], w995, w996);
  FullAdder U285 (w996, w879, IN50[5], w997, w998);
  FullAdder U286 (w998, w881, IN51[5], w999, w1000);
  FullAdder U287 (w1000, w883, IN52[5], w1001, w1002);
  FullAdder U288 (w1002, w885, IN53[5], w1003, w1004);
  FullAdder U289 (w1004, w887, IN54[5], w1005, w1006);
  FullAdder U290 (w1006, w889, IN55[5], w1007, w1008);
  FullAdder U291 (w1008, w891, IN56[5], w1009, w1010);
  FullAdder U292 (w1010, w893, IN57[5], w1011, w1012);
  FullAdder U293 (w1012, w895, IN58[5], w1013, w1014);
  FullAdder U294 (w1014, w897, IN59[5], w1015, w1016);
  FullAdder U295 (w1016, w899, IN60[5], w1017, w1018);
  FullAdder U296 (w1018, w901, IN61[3], w1019, w1020);
  FullAdder U297 (w1020, w903, IN62[2], w1021, w1022);
  FullAdder U298 (w1022, w905, IN63[1], w1023, w1024);
  FullAdder U299 (w1024, w906, IN64[0], w1025, w1026);
  HalfAdder U300 (w909, IN6[6], Out1[6], w1028);
  FullAdder U301 (w1028, w911, IN7[6], Out1[7], w1030);
  FullAdder U302 (w1030, w913, IN8[6], Out1[8], w1032);
  FullAdder U303 (w1032, w915, IN9[6], Out1[9], w1034);
  FullAdder U304 (w1034, w917, IN10[6], Out1[10], w1036);
  FullAdder U305 (w1036, w919, IN11[6], Out1[11], w1038);
  FullAdder U306 (w1038, w921, IN12[6], Out1[12], w1040);
  FullAdder U307 (w1040, w923, IN13[6], Out1[13], w1042);
  FullAdder U308 (w1042, w925, IN14[6], Out1[14], w1044);
  FullAdder U309 (w1044, w927, IN15[6], Out1[15], w1046);
  FullAdder U310 (w1046, w929, IN16[6], Out1[16], w1048);
  FullAdder U311 (w1048, w931, IN17[6], Out1[17], w1050);
  FullAdder U312 (w1050, w933, IN18[6], Out1[18], w1052);
  FullAdder U313 (w1052, w935, IN19[6], Out1[19], w1054);
  FullAdder U314 (w1054, w937, IN20[6], Out1[20], w1056);
  FullAdder U315 (w1056, w939, IN21[6], Out1[21], w1058);
  FullAdder U316 (w1058, w941, IN22[6], Out1[22], w1060);
  FullAdder U317 (w1060, w943, IN23[6], Out1[23], w1062);
  FullAdder U318 (w1062, w945, IN24[6], Out1[24], w1064);
  FullAdder U319 (w1064, w947, IN25[6], Out1[25], w1066);
  FullAdder U320 (w1066, w949, IN26[6], Out1[26], w1068);
  FullAdder U321 (w1068, w951, IN27[6], Out1[27], w1070);
  FullAdder U322 (w1070, w953, IN28[6], Out1[28], w1072);
  FullAdder U323 (w1072, w955, IN29[6], Out1[29], w1074);
  FullAdder U324 (w1074, w957, IN30[6], Out1[30], w1076);
  FullAdder U325 (w1076, w959, IN31[6], Out1[31], w1078);
  FullAdder U326 (w1078, w961, IN32[6], Out1[32], w1080);
  FullAdder U327 (w1080, w963, IN33[6], Out1[33], w1082);
  FullAdder U328 (w1082, w965, IN34[6], Out1[34], w1084);
  FullAdder U329 (w1084, w967, IN35[6], Out1[35], w1086);
  FullAdder U330 (w1086, w969, IN36[6], Out1[36], w1088);
  FullAdder U331 (w1088, w971, IN37[6], Out1[37], w1090);
  FullAdder U332 (w1090, w973, IN38[6], Out1[38], w1092);
  FullAdder U333 (w1092, w975, IN39[6], Out1[39], w1094);
  FullAdder U334 (w1094, w977, IN40[6], Out1[40], w1096);
  FullAdder U335 (w1096, w979, IN41[6], Out1[41], w1098);
  FullAdder U336 (w1098, w981, IN42[6], Out1[42], w1100);
  FullAdder U337 (w1100, w983, IN43[6], Out1[43], w1102);
  FullAdder U338 (w1102, w985, IN44[6], Out1[44], w1104);
  FullAdder U339 (w1104, w987, IN45[6], Out1[45], w1106);
  FullAdder U340 (w1106, w989, IN46[6], Out1[46], w1108);
  FullAdder U341 (w1108, w991, IN47[6], Out1[47], w1110);
  FullAdder U342 (w1110, w993, IN48[6], Out1[48], w1112);
  FullAdder U343 (w1112, w995, IN49[6], Out1[49], w1114);
  FullAdder U344 (w1114, w997, IN50[6], Out1[50], w1116);
  FullAdder U345 (w1116, w999, IN51[6], Out1[51], w1118);
  FullAdder U346 (w1118, w1001, IN52[6], Out1[52], w1120);
  FullAdder U347 (w1120, w1003, IN53[6], Out1[53], w1122);
  FullAdder U348 (w1122, w1005, IN54[6], Out1[54], w1124);
  FullAdder U349 (w1124, w1007, IN55[6], Out1[55], w1126);
  FullAdder U350 (w1126, w1009, IN56[6], Out1[56], w1128);
  FullAdder U351 (w1128, w1011, IN57[6], Out1[57], w1130);
  FullAdder U352 (w1130, w1013, IN58[6], Out1[58], w1132);
  FullAdder U353 (w1132, w1015, IN59[6], Out1[59], w1134);
  FullAdder U354 (w1134, w1017, IN60[6], Out1[60], w1136);
  FullAdder U355 (w1136, w1019, IN61[4], Out1[61], w1138);
  FullAdder U356 (w1138, w1021, IN62[3], Out1[62], w1140);
  FullAdder U357 (w1140, w1023, IN63[2], Out1[63], w1142);
  FullAdder U358 (w1142, w1025, IN64[1], Out1[64], w1144);
  FullAdder U359 (w1144, w1026, IN65[0], Out1[65], Out1[66]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN61[5];
  assign Out2[1] = IN62[4];
  assign Out2[2] = IN63[3];
  assign Out2[3] = IN64[2];
  assign Out2[4] = IN65[1];
  assign Out2[5] = IN66[0];

endmodule
module RC_6_6(IN1, IN2, Out);
  input [5:0] IN1;
  input [5:0] IN2;
  output [6:0] Out;
  wire w13;
  wire w15;
  wire w17;
  wire w19;
  wire w21;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w13);
  FullAdder U1 (IN1[1], IN2[1], w13, Out[1], w15);
  FullAdder U2 (IN1[2], IN2[2], w15, Out[2], w17);
  FullAdder U3 (IN1[3], IN2[3], w17, Out[3], w19);
  FullAdder U4 (IN1[4], IN2[4], w19, Out[4], w21);
  FullAdder U5 (IN1[5], IN2[5], w21, Out[5], Out[6]);

endmodule
module NR_61_7(IN1, IN2, Out);
  input [60:0] IN1;
  input [6:0] IN2;
  output [67:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [6:0] P37;
  wire [6:0] P38;
  wire [6:0] P39;
  wire [6:0] P40;
  wire [6:0] P41;
  wire [6:0] P42;
  wire [6:0] P43;
  wire [6:0] P44;
  wire [6:0] P45;
  wire [6:0] P46;
  wire [6:0] P47;
  wire [6:0] P48;
  wire [6:0] P49;
  wire [6:0] P50;
  wire [6:0] P51;
  wire [6:0] P52;
  wire [6:0] P53;
  wire [6:0] P54;
  wire [6:0] P55;
  wire [6:0] P56;
  wire [6:0] P57;
  wire [6:0] P58;
  wire [6:0] P59;
  wire [6:0] P60;
  wire [5:0] P61;
  wire [4:0] P62;
  wire [3:0] P63;
  wire [2:0] P64;
  wire [1:0] P65;
  wire [0:0] P66;
  wire [66:0] R1;
  wire [5:0] R2;
  wire [67:0] aOut;
  U_SP_61_7 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, R1, R2);
  RC_6_6 S2 (R1[66:61], R2, aOut[67:61]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign aOut[57] = R1[57];
  assign aOut[58] = R1[58];
  assign aOut[59] = R1[59];
  assign aOut[60] = R1[60];
  assign Out = aOut[67:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
