
module customAdder44_0(
    input [43 : 0] A,
    input [43 : 0] B,
    output [44 : 0] Sum
);

    assign Sum = A+B;

endmodule
