//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 8
  second input length: 56
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_8_56(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  input [7:0] IN1;
  input [55:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [7:0] P8;
  output [7:0] P9;
  output [7:0] P10;
  output [7:0] P11;
  output [7:0] P12;
  output [7:0] P13;
  output [7:0] P14;
  output [7:0] P15;
  output [7:0] P16;
  output [7:0] P17;
  output [7:0] P18;
  output [7:0] P19;
  output [7:0] P20;
  output [7:0] P21;
  output [7:0] P22;
  output [7:0] P23;
  output [7:0] P24;
  output [7:0] P25;
  output [7:0] P26;
  output [7:0] P27;
  output [7:0] P28;
  output [7:0] P29;
  output [7:0] P30;
  output [7:0] P31;
  output [7:0] P32;
  output [7:0] P33;
  output [7:0] P34;
  output [7:0] P35;
  output [7:0] P36;
  output [7:0] P37;
  output [7:0] P38;
  output [7:0] P39;
  output [7:0] P40;
  output [7:0] P41;
  output [7:0] P42;
  output [7:0] P43;
  output [7:0] P44;
  output [7:0] P45;
  output [7:0] P46;
  output [7:0] P47;
  output [7:0] P48;
  output [7:0] P49;
  output [7:0] P50;
  output [7:0] P51;
  output [7:0] P52;
  output [7:0] P53;
  output [7:0] P54;
  output [7:0] P55;
  output [6:0] P56;
  output [5:0] P57;
  output [4:0] P58;
  output [3:0] P59;
  output [2:0] P60;
  output [1:0] P61;
  output [0:0] P62;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[0] = IN1[1]&IN2[55];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[1] = IN1[2]&IN2[54];
  assign P57[0] = IN1[2]&IN2[55];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[2] = IN1[3]&IN2[53];
  assign P57[1] = IN1[3]&IN2[54];
  assign P58[0] = IN1[3]&IN2[55];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[3] = IN1[4]&IN2[52];
  assign P57[2] = IN1[4]&IN2[53];
  assign P58[1] = IN1[4]&IN2[54];
  assign P59[0] = IN1[4]&IN2[55];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[4] = IN1[5]&IN2[51];
  assign P57[3] = IN1[5]&IN2[52];
  assign P58[2] = IN1[5]&IN2[53];
  assign P59[1] = IN1[5]&IN2[54];
  assign P60[0] = IN1[5]&IN2[55];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[5] = IN1[6]&IN2[50];
  assign P57[4] = IN1[6]&IN2[51];
  assign P58[3] = IN1[6]&IN2[52];
  assign P59[2] = IN1[6]&IN2[53];
  assign P60[1] = IN1[6]&IN2[54];
  assign P61[0] = IN1[6]&IN2[55];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[7] = IN1[7]&IN2[47];
  assign P55[7] = IN1[7]&IN2[48];
  assign P56[6] = IN1[7]&IN2[49];
  assign P57[5] = IN1[7]&IN2[50];
  assign P58[4] = IN1[7]&IN2[51];
  assign P59[3] = IN1[7]&IN2[52];
  assign P60[2] = IN1[7]&IN2[53];
  assign P61[1] = IN1[7]&IN2[54];
  assign P62[0] = IN1[7]&IN2[55];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [7:0] IN8;
  input [7:0] IN9;
  input [7:0] IN10;
  input [7:0] IN11;
  input [7:0] IN12;
  input [7:0] IN13;
  input [7:0] IN14;
  input [7:0] IN15;
  input [7:0] IN16;
  input [7:0] IN17;
  input [7:0] IN18;
  input [7:0] IN19;
  input [7:0] IN20;
  input [7:0] IN21;
  input [7:0] IN22;
  input [7:0] IN23;
  input [7:0] IN24;
  input [7:0] IN25;
  input [7:0] IN26;
  input [7:0] IN27;
  input [7:0] IN28;
  input [7:0] IN29;
  input [7:0] IN30;
  input [7:0] IN31;
  input [7:0] IN32;
  input [7:0] IN33;
  input [7:0] IN34;
  input [7:0] IN35;
  input [7:0] IN36;
  input [7:0] IN37;
  input [7:0] IN38;
  input [7:0] IN39;
  input [7:0] IN40;
  input [7:0] IN41;
  input [7:0] IN42;
  input [7:0] IN43;
  input [7:0] IN44;
  input [7:0] IN45;
  input [7:0] IN46;
  input [7:0] IN47;
  input [7:0] IN48;
  input [7:0] IN49;
  input [7:0] IN50;
  input [7:0] IN51;
  input [7:0] IN52;
  input [7:0] IN53;
  input [7:0] IN54;
  input [7:0] IN55;
  input [6:0] IN56;
  input [5:0] IN57;
  input [4:0] IN58;
  input [3:0] IN59;
  input [2:0] IN60;
  input [1:0] IN61;
  input [0:0] IN62;
  output [62:0] Out1;
  output [54:0] Out2;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1205;
  wire w1207;
  wire w1209;
  wire w1211;
  wire w1213;
  wire w1215;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w449);
  FullAdder U1 (w449, IN2[0], IN2[1], w450, w451);
  FullAdder U2 (w451, IN3[0], IN3[1], w452, w453);
  FullAdder U3 (w453, IN4[0], IN4[1], w454, w455);
  FullAdder U4 (w455, IN5[0], IN5[1], w456, w457);
  FullAdder U5 (w457, IN6[0], IN6[1], w458, w459);
  FullAdder U6 (w459, IN7[0], IN7[1], w460, w461);
  HalfAdder U7 (w450, IN2[2], Out1[2], w463);
  FullAdder U8 (w463, w452, IN3[2], w464, w465);
  FullAdder U9 (w465, w454, IN4[2], w466, w467);
  FullAdder U10 (w467, w456, IN5[2], w468, w469);
  FullAdder U11 (w469, w458, IN6[2], w470, w471);
  FullAdder U12 (w471, w460, IN7[2], w472, w473);
  FullAdder U13 (w473, w461, IN8[0], w474, w475);
  HalfAdder U14 (w464, IN3[3], Out1[3], w477);
  FullAdder U15 (w477, w466, IN4[3], w478, w479);
  FullAdder U16 (w479, w468, IN5[3], w480, w481);
  FullAdder U17 (w481, w470, IN6[3], w482, w483);
  FullAdder U18 (w483, w472, IN7[3], w484, w485);
  FullAdder U19 (w485, w474, IN8[1], w486, w487);
  FullAdder U20 (w487, w475, IN9[0], w488, w489);
  HalfAdder U21 (w478, IN4[4], Out1[4], w491);
  FullAdder U22 (w491, w480, IN5[4], w492, w493);
  FullAdder U23 (w493, w482, IN6[4], w494, w495);
  FullAdder U24 (w495, w484, IN7[4], w496, w497);
  FullAdder U25 (w497, w486, IN8[2], w498, w499);
  FullAdder U26 (w499, w488, IN9[1], w500, w501);
  FullAdder U27 (w501, w489, IN10[0], w502, w503);
  HalfAdder U28 (w492, IN5[5], Out1[5], w505);
  FullAdder U29 (w505, w494, IN6[5], w506, w507);
  FullAdder U30 (w507, w496, IN7[5], w508, w509);
  FullAdder U31 (w509, w498, IN8[3], w510, w511);
  FullAdder U32 (w511, w500, IN9[2], w512, w513);
  FullAdder U33 (w513, w502, IN10[1], w514, w515);
  FullAdder U34 (w515, w503, IN11[0], w516, w517);
  HalfAdder U35 (w506, IN6[6], Out1[6], w519);
  FullAdder U36 (w519, w508, IN7[6], w520, w521);
  FullAdder U37 (w521, w510, IN8[4], w522, w523);
  FullAdder U38 (w523, w512, IN9[3], w524, w525);
  FullAdder U39 (w525, w514, IN10[2], w526, w527);
  FullAdder U40 (w527, w516, IN11[1], w528, w529);
  FullAdder U41 (w529, w517, IN12[0], w530, w531);
  HalfAdder U42 (w520, IN7[7], Out1[7], w533);
  FullAdder U43 (w533, w522, IN8[5], w534, w535);
  FullAdder U44 (w535, w524, IN9[4], w536, w537);
  FullAdder U45 (w537, w526, IN10[3], w538, w539);
  FullAdder U46 (w539, w528, IN11[2], w540, w541);
  FullAdder U47 (w541, w530, IN12[1], w542, w543);
  FullAdder U48 (w543, w531, IN13[0], w544, w545);
  HalfAdder U49 (w534, IN8[6], Out1[8], w547);
  FullAdder U50 (w547, w536, IN9[5], w548, w549);
  FullAdder U51 (w549, w538, IN10[4], w550, w551);
  FullAdder U52 (w551, w540, IN11[3], w552, w553);
  FullAdder U53 (w553, w542, IN12[2], w554, w555);
  FullAdder U54 (w555, w544, IN13[1], w556, w557);
  FullAdder U55 (w557, w545, IN14[0], w558, w559);
  HalfAdder U56 (w548, IN9[6], Out1[9], w561);
  FullAdder U57 (w561, w550, IN10[5], w562, w563);
  FullAdder U58 (w563, w552, IN11[4], w564, w565);
  FullAdder U59 (w565, w554, IN12[3], w566, w567);
  FullAdder U60 (w567, w556, IN13[2], w568, w569);
  FullAdder U61 (w569, w558, IN14[1], w570, w571);
  FullAdder U62 (w571, w559, IN15[0], w572, w573);
  HalfAdder U63 (w562, IN10[6], Out1[10], w575);
  FullAdder U64 (w575, w564, IN11[5], w576, w577);
  FullAdder U65 (w577, w566, IN12[4], w578, w579);
  FullAdder U66 (w579, w568, IN13[3], w580, w581);
  FullAdder U67 (w581, w570, IN14[2], w582, w583);
  FullAdder U68 (w583, w572, IN15[1], w584, w585);
  FullAdder U69 (w585, w573, IN16[0], w586, w587);
  HalfAdder U70 (w576, IN11[6], Out1[11], w589);
  FullAdder U71 (w589, w578, IN12[5], w590, w591);
  FullAdder U72 (w591, w580, IN13[4], w592, w593);
  FullAdder U73 (w593, w582, IN14[3], w594, w595);
  FullAdder U74 (w595, w584, IN15[2], w596, w597);
  FullAdder U75 (w597, w586, IN16[1], w598, w599);
  FullAdder U76 (w599, w587, IN17[0], w600, w601);
  HalfAdder U77 (w590, IN12[6], Out1[12], w603);
  FullAdder U78 (w603, w592, IN13[5], w604, w605);
  FullAdder U79 (w605, w594, IN14[4], w606, w607);
  FullAdder U80 (w607, w596, IN15[3], w608, w609);
  FullAdder U81 (w609, w598, IN16[2], w610, w611);
  FullAdder U82 (w611, w600, IN17[1], w612, w613);
  FullAdder U83 (w613, w601, IN18[0], w614, w615);
  HalfAdder U84 (w604, IN13[6], Out1[13], w617);
  FullAdder U85 (w617, w606, IN14[5], w618, w619);
  FullAdder U86 (w619, w608, IN15[4], w620, w621);
  FullAdder U87 (w621, w610, IN16[3], w622, w623);
  FullAdder U88 (w623, w612, IN17[2], w624, w625);
  FullAdder U89 (w625, w614, IN18[1], w626, w627);
  FullAdder U90 (w627, w615, IN19[0], w628, w629);
  HalfAdder U91 (w618, IN14[6], Out1[14], w631);
  FullAdder U92 (w631, w620, IN15[5], w632, w633);
  FullAdder U93 (w633, w622, IN16[4], w634, w635);
  FullAdder U94 (w635, w624, IN17[3], w636, w637);
  FullAdder U95 (w637, w626, IN18[2], w638, w639);
  FullAdder U96 (w639, w628, IN19[1], w640, w641);
  FullAdder U97 (w641, w629, IN20[0], w642, w643);
  HalfAdder U98 (w632, IN15[6], Out1[15], w645);
  FullAdder U99 (w645, w634, IN16[5], w646, w647);
  FullAdder U100 (w647, w636, IN17[4], w648, w649);
  FullAdder U101 (w649, w638, IN18[3], w650, w651);
  FullAdder U102 (w651, w640, IN19[2], w652, w653);
  FullAdder U103 (w653, w642, IN20[1], w654, w655);
  FullAdder U104 (w655, w643, IN21[0], w656, w657);
  HalfAdder U105 (w646, IN16[6], Out1[16], w659);
  FullAdder U106 (w659, w648, IN17[5], w660, w661);
  FullAdder U107 (w661, w650, IN18[4], w662, w663);
  FullAdder U108 (w663, w652, IN19[3], w664, w665);
  FullAdder U109 (w665, w654, IN20[2], w666, w667);
  FullAdder U110 (w667, w656, IN21[1], w668, w669);
  FullAdder U111 (w669, w657, IN22[0], w670, w671);
  HalfAdder U112 (w660, IN17[6], Out1[17], w673);
  FullAdder U113 (w673, w662, IN18[5], w674, w675);
  FullAdder U114 (w675, w664, IN19[4], w676, w677);
  FullAdder U115 (w677, w666, IN20[3], w678, w679);
  FullAdder U116 (w679, w668, IN21[2], w680, w681);
  FullAdder U117 (w681, w670, IN22[1], w682, w683);
  FullAdder U118 (w683, w671, IN23[0], w684, w685);
  HalfAdder U119 (w674, IN18[6], Out1[18], w687);
  FullAdder U120 (w687, w676, IN19[5], w688, w689);
  FullAdder U121 (w689, w678, IN20[4], w690, w691);
  FullAdder U122 (w691, w680, IN21[3], w692, w693);
  FullAdder U123 (w693, w682, IN22[2], w694, w695);
  FullAdder U124 (w695, w684, IN23[1], w696, w697);
  FullAdder U125 (w697, w685, IN24[0], w698, w699);
  HalfAdder U126 (w688, IN19[6], Out1[19], w701);
  FullAdder U127 (w701, w690, IN20[5], w702, w703);
  FullAdder U128 (w703, w692, IN21[4], w704, w705);
  FullAdder U129 (w705, w694, IN22[3], w706, w707);
  FullAdder U130 (w707, w696, IN23[2], w708, w709);
  FullAdder U131 (w709, w698, IN24[1], w710, w711);
  FullAdder U132 (w711, w699, IN25[0], w712, w713);
  HalfAdder U133 (w702, IN20[6], Out1[20], w715);
  FullAdder U134 (w715, w704, IN21[5], w716, w717);
  FullAdder U135 (w717, w706, IN22[4], w718, w719);
  FullAdder U136 (w719, w708, IN23[3], w720, w721);
  FullAdder U137 (w721, w710, IN24[2], w722, w723);
  FullAdder U138 (w723, w712, IN25[1], w724, w725);
  FullAdder U139 (w725, w713, IN26[0], w726, w727);
  HalfAdder U140 (w716, IN21[6], Out1[21], w729);
  FullAdder U141 (w729, w718, IN22[5], w730, w731);
  FullAdder U142 (w731, w720, IN23[4], w732, w733);
  FullAdder U143 (w733, w722, IN24[3], w734, w735);
  FullAdder U144 (w735, w724, IN25[2], w736, w737);
  FullAdder U145 (w737, w726, IN26[1], w738, w739);
  FullAdder U146 (w739, w727, IN27[0], w740, w741);
  HalfAdder U147 (w730, IN22[6], Out1[22], w743);
  FullAdder U148 (w743, w732, IN23[5], w744, w745);
  FullAdder U149 (w745, w734, IN24[4], w746, w747);
  FullAdder U150 (w747, w736, IN25[3], w748, w749);
  FullAdder U151 (w749, w738, IN26[2], w750, w751);
  FullAdder U152 (w751, w740, IN27[1], w752, w753);
  FullAdder U153 (w753, w741, IN28[0], w754, w755);
  HalfAdder U154 (w744, IN23[6], Out1[23], w757);
  FullAdder U155 (w757, w746, IN24[5], w758, w759);
  FullAdder U156 (w759, w748, IN25[4], w760, w761);
  FullAdder U157 (w761, w750, IN26[3], w762, w763);
  FullAdder U158 (w763, w752, IN27[2], w764, w765);
  FullAdder U159 (w765, w754, IN28[1], w766, w767);
  FullAdder U160 (w767, w755, IN29[0], w768, w769);
  HalfAdder U161 (w758, IN24[6], Out1[24], w771);
  FullAdder U162 (w771, w760, IN25[5], w772, w773);
  FullAdder U163 (w773, w762, IN26[4], w774, w775);
  FullAdder U164 (w775, w764, IN27[3], w776, w777);
  FullAdder U165 (w777, w766, IN28[2], w778, w779);
  FullAdder U166 (w779, w768, IN29[1], w780, w781);
  FullAdder U167 (w781, w769, IN30[0], w782, w783);
  HalfAdder U168 (w772, IN25[6], Out1[25], w785);
  FullAdder U169 (w785, w774, IN26[5], w786, w787);
  FullAdder U170 (w787, w776, IN27[4], w788, w789);
  FullAdder U171 (w789, w778, IN28[3], w790, w791);
  FullAdder U172 (w791, w780, IN29[2], w792, w793);
  FullAdder U173 (w793, w782, IN30[1], w794, w795);
  FullAdder U174 (w795, w783, IN31[0], w796, w797);
  HalfAdder U175 (w786, IN26[6], Out1[26], w799);
  FullAdder U176 (w799, w788, IN27[5], w800, w801);
  FullAdder U177 (w801, w790, IN28[4], w802, w803);
  FullAdder U178 (w803, w792, IN29[3], w804, w805);
  FullAdder U179 (w805, w794, IN30[2], w806, w807);
  FullAdder U180 (w807, w796, IN31[1], w808, w809);
  FullAdder U181 (w809, w797, IN32[0], w810, w811);
  HalfAdder U182 (w800, IN27[6], Out1[27], w813);
  FullAdder U183 (w813, w802, IN28[5], w814, w815);
  FullAdder U184 (w815, w804, IN29[4], w816, w817);
  FullAdder U185 (w817, w806, IN30[3], w818, w819);
  FullAdder U186 (w819, w808, IN31[2], w820, w821);
  FullAdder U187 (w821, w810, IN32[1], w822, w823);
  FullAdder U188 (w823, w811, IN33[0], w824, w825);
  HalfAdder U189 (w814, IN28[6], Out1[28], w827);
  FullAdder U190 (w827, w816, IN29[5], w828, w829);
  FullAdder U191 (w829, w818, IN30[4], w830, w831);
  FullAdder U192 (w831, w820, IN31[3], w832, w833);
  FullAdder U193 (w833, w822, IN32[2], w834, w835);
  FullAdder U194 (w835, w824, IN33[1], w836, w837);
  FullAdder U195 (w837, w825, IN34[0], w838, w839);
  HalfAdder U196 (w828, IN29[6], Out1[29], w841);
  FullAdder U197 (w841, w830, IN30[5], w842, w843);
  FullAdder U198 (w843, w832, IN31[4], w844, w845);
  FullAdder U199 (w845, w834, IN32[3], w846, w847);
  FullAdder U200 (w847, w836, IN33[2], w848, w849);
  FullAdder U201 (w849, w838, IN34[1], w850, w851);
  FullAdder U202 (w851, w839, IN35[0], w852, w853);
  HalfAdder U203 (w842, IN30[6], Out1[30], w855);
  FullAdder U204 (w855, w844, IN31[5], w856, w857);
  FullAdder U205 (w857, w846, IN32[4], w858, w859);
  FullAdder U206 (w859, w848, IN33[3], w860, w861);
  FullAdder U207 (w861, w850, IN34[2], w862, w863);
  FullAdder U208 (w863, w852, IN35[1], w864, w865);
  FullAdder U209 (w865, w853, IN36[0], w866, w867);
  HalfAdder U210 (w856, IN31[6], Out1[31], w869);
  FullAdder U211 (w869, w858, IN32[5], w870, w871);
  FullAdder U212 (w871, w860, IN33[4], w872, w873);
  FullAdder U213 (w873, w862, IN34[3], w874, w875);
  FullAdder U214 (w875, w864, IN35[2], w876, w877);
  FullAdder U215 (w877, w866, IN36[1], w878, w879);
  FullAdder U216 (w879, w867, IN37[0], w880, w881);
  HalfAdder U217 (w870, IN32[6], Out1[32], w883);
  FullAdder U218 (w883, w872, IN33[5], w884, w885);
  FullAdder U219 (w885, w874, IN34[4], w886, w887);
  FullAdder U220 (w887, w876, IN35[3], w888, w889);
  FullAdder U221 (w889, w878, IN36[2], w890, w891);
  FullAdder U222 (w891, w880, IN37[1], w892, w893);
  FullAdder U223 (w893, w881, IN38[0], w894, w895);
  HalfAdder U224 (w884, IN33[6], Out1[33], w897);
  FullAdder U225 (w897, w886, IN34[5], w898, w899);
  FullAdder U226 (w899, w888, IN35[4], w900, w901);
  FullAdder U227 (w901, w890, IN36[3], w902, w903);
  FullAdder U228 (w903, w892, IN37[2], w904, w905);
  FullAdder U229 (w905, w894, IN38[1], w906, w907);
  FullAdder U230 (w907, w895, IN39[0], w908, w909);
  HalfAdder U231 (w898, IN34[6], Out1[34], w911);
  FullAdder U232 (w911, w900, IN35[5], w912, w913);
  FullAdder U233 (w913, w902, IN36[4], w914, w915);
  FullAdder U234 (w915, w904, IN37[3], w916, w917);
  FullAdder U235 (w917, w906, IN38[2], w918, w919);
  FullAdder U236 (w919, w908, IN39[1], w920, w921);
  FullAdder U237 (w921, w909, IN40[0], w922, w923);
  HalfAdder U238 (w912, IN35[6], Out1[35], w925);
  FullAdder U239 (w925, w914, IN36[5], w926, w927);
  FullAdder U240 (w927, w916, IN37[4], w928, w929);
  FullAdder U241 (w929, w918, IN38[3], w930, w931);
  FullAdder U242 (w931, w920, IN39[2], w932, w933);
  FullAdder U243 (w933, w922, IN40[1], w934, w935);
  FullAdder U244 (w935, w923, IN41[0], w936, w937);
  HalfAdder U245 (w926, IN36[6], Out1[36], w939);
  FullAdder U246 (w939, w928, IN37[5], w940, w941);
  FullAdder U247 (w941, w930, IN38[4], w942, w943);
  FullAdder U248 (w943, w932, IN39[3], w944, w945);
  FullAdder U249 (w945, w934, IN40[2], w946, w947);
  FullAdder U250 (w947, w936, IN41[1], w948, w949);
  FullAdder U251 (w949, w937, IN42[0], w950, w951);
  HalfAdder U252 (w940, IN37[6], Out1[37], w953);
  FullAdder U253 (w953, w942, IN38[5], w954, w955);
  FullAdder U254 (w955, w944, IN39[4], w956, w957);
  FullAdder U255 (w957, w946, IN40[3], w958, w959);
  FullAdder U256 (w959, w948, IN41[2], w960, w961);
  FullAdder U257 (w961, w950, IN42[1], w962, w963);
  FullAdder U258 (w963, w951, IN43[0], w964, w965);
  HalfAdder U259 (w954, IN38[6], Out1[38], w967);
  FullAdder U260 (w967, w956, IN39[5], w968, w969);
  FullAdder U261 (w969, w958, IN40[4], w970, w971);
  FullAdder U262 (w971, w960, IN41[3], w972, w973);
  FullAdder U263 (w973, w962, IN42[2], w974, w975);
  FullAdder U264 (w975, w964, IN43[1], w976, w977);
  FullAdder U265 (w977, w965, IN44[0], w978, w979);
  HalfAdder U266 (w968, IN39[6], Out1[39], w981);
  FullAdder U267 (w981, w970, IN40[5], w982, w983);
  FullAdder U268 (w983, w972, IN41[4], w984, w985);
  FullAdder U269 (w985, w974, IN42[3], w986, w987);
  FullAdder U270 (w987, w976, IN43[2], w988, w989);
  FullAdder U271 (w989, w978, IN44[1], w990, w991);
  FullAdder U272 (w991, w979, IN45[0], w992, w993);
  HalfAdder U273 (w982, IN40[6], Out1[40], w995);
  FullAdder U274 (w995, w984, IN41[5], w996, w997);
  FullAdder U275 (w997, w986, IN42[4], w998, w999);
  FullAdder U276 (w999, w988, IN43[3], w1000, w1001);
  FullAdder U277 (w1001, w990, IN44[2], w1002, w1003);
  FullAdder U278 (w1003, w992, IN45[1], w1004, w1005);
  FullAdder U279 (w1005, w993, IN46[0], w1006, w1007);
  HalfAdder U280 (w996, IN41[6], Out1[41], w1009);
  FullAdder U281 (w1009, w998, IN42[5], w1010, w1011);
  FullAdder U282 (w1011, w1000, IN43[4], w1012, w1013);
  FullAdder U283 (w1013, w1002, IN44[3], w1014, w1015);
  FullAdder U284 (w1015, w1004, IN45[2], w1016, w1017);
  FullAdder U285 (w1017, w1006, IN46[1], w1018, w1019);
  FullAdder U286 (w1019, w1007, IN47[0], w1020, w1021);
  HalfAdder U287 (w1010, IN42[6], Out1[42], w1023);
  FullAdder U288 (w1023, w1012, IN43[5], w1024, w1025);
  FullAdder U289 (w1025, w1014, IN44[4], w1026, w1027);
  FullAdder U290 (w1027, w1016, IN45[3], w1028, w1029);
  FullAdder U291 (w1029, w1018, IN46[2], w1030, w1031);
  FullAdder U292 (w1031, w1020, IN47[1], w1032, w1033);
  FullAdder U293 (w1033, w1021, IN48[0], w1034, w1035);
  HalfAdder U294 (w1024, IN43[6], Out1[43], w1037);
  FullAdder U295 (w1037, w1026, IN44[5], w1038, w1039);
  FullAdder U296 (w1039, w1028, IN45[4], w1040, w1041);
  FullAdder U297 (w1041, w1030, IN46[3], w1042, w1043);
  FullAdder U298 (w1043, w1032, IN47[2], w1044, w1045);
  FullAdder U299 (w1045, w1034, IN48[1], w1046, w1047);
  FullAdder U300 (w1047, w1035, IN49[0], w1048, w1049);
  HalfAdder U301 (w1038, IN44[6], Out1[44], w1051);
  FullAdder U302 (w1051, w1040, IN45[5], w1052, w1053);
  FullAdder U303 (w1053, w1042, IN46[4], w1054, w1055);
  FullAdder U304 (w1055, w1044, IN47[3], w1056, w1057);
  FullAdder U305 (w1057, w1046, IN48[2], w1058, w1059);
  FullAdder U306 (w1059, w1048, IN49[1], w1060, w1061);
  FullAdder U307 (w1061, w1049, IN50[0], w1062, w1063);
  HalfAdder U308 (w1052, IN45[6], Out1[45], w1065);
  FullAdder U309 (w1065, w1054, IN46[5], w1066, w1067);
  FullAdder U310 (w1067, w1056, IN47[4], w1068, w1069);
  FullAdder U311 (w1069, w1058, IN48[3], w1070, w1071);
  FullAdder U312 (w1071, w1060, IN49[2], w1072, w1073);
  FullAdder U313 (w1073, w1062, IN50[1], w1074, w1075);
  FullAdder U314 (w1075, w1063, IN51[0], w1076, w1077);
  HalfAdder U315 (w1066, IN46[6], Out1[46], w1079);
  FullAdder U316 (w1079, w1068, IN47[5], w1080, w1081);
  FullAdder U317 (w1081, w1070, IN48[4], w1082, w1083);
  FullAdder U318 (w1083, w1072, IN49[3], w1084, w1085);
  FullAdder U319 (w1085, w1074, IN50[2], w1086, w1087);
  FullAdder U320 (w1087, w1076, IN51[1], w1088, w1089);
  FullAdder U321 (w1089, w1077, IN52[0], w1090, w1091);
  HalfAdder U322 (w1080, IN47[6], Out1[47], w1093);
  FullAdder U323 (w1093, w1082, IN48[5], w1094, w1095);
  FullAdder U324 (w1095, w1084, IN49[4], w1096, w1097);
  FullAdder U325 (w1097, w1086, IN50[3], w1098, w1099);
  FullAdder U326 (w1099, w1088, IN51[2], w1100, w1101);
  FullAdder U327 (w1101, w1090, IN52[1], w1102, w1103);
  FullAdder U328 (w1103, w1091, IN53[0], w1104, w1105);
  HalfAdder U329 (w1094, IN48[6], Out1[48], w1107);
  FullAdder U330 (w1107, w1096, IN49[5], w1108, w1109);
  FullAdder U331 (w1109, w1098, IN50[4], w1110, w1111);
  FullAdder U332 (w1111, w1100, IN51[3], w1112, w1113);
  FullAdder U333 (w1113, w1102, IN52[2], w1114, w1115);
  FullAdder U334 (w1115, w1104, IN53[1], w1116, w1117);
  FullAdder U335 (w1117, w1105, IN54[0], w1118, w1119);
  HalfAdder U336 (w1108, IN49[6], Out1[49], w1121);
  FullAdder U337 (w1121, w1110, IN50[5], w1122, w1123);
  FullAdder U338 (w1123, w1112, IN51[4], w1124, w1125);
  FullAdder U339 (w1125, w1114, IN52[3], w1126, w1127);
  FullAdder U340 (w1127, w1116, IN53[2], w1128, w1129);
  FullAdder U341 (w1129, w1118, IN54[1], w1130, w1131);
  FullAdder U342 (w1131, w1119, IN55[0], w1132, w1133);
  HalfAdder U343 (w1122, IN50[6], Out1[50], w1135);
  FullAdder U344 (w1135, w1124, IN51[5], w1136, w1137);
  FullAdder U345 (w1137, w1126, IN52[4], w1138, w1139);
  FullAdder U346 (w1139, w1128, IN53[3], w1140, w1141);
  FullAdder U347 (w1141, w1130, IN54[2], w1142, w1143);
  FullAdder U348 (w1143, w1132, IN55[1], w1144, w1145);
  FullAdder U349 (w1145, w1133, IN56[0], w1146, w1147);
  HalfAdder U350 (w1136, IN51[6], Out1[51], w1149);
  FullAdder U351 (w1149, w1138, IN52[5], w1150, w1151);
  FullAdder U352 (w1151, w1140, IN53[4], w1152, w1153);
  FullAdder U353 (w1153, w1142, IN54[3], w1154, w1155);
  FullAdder U354 (w1155, w1144, IN55[2], w1156, w1157);
  FullAdder U355 (w1157, w1146, IN56[1], w1158, w1159);
  FullAdder U356 (w1159, w1147, IN57[0], w1160, w1161);
  HalfAdder U357 (w1150, IN52[6], Out1[52], w1163);
  FullAdder U358 (w1163, w1152, IN53[5], w1164, w1165);
  FullAdder U359 (w1165, w1154, IN54[4], w1166, w1167);
  FullAdder U360 (w1167, w1156, IN55[3], w1168, w1169);
  FullAdder U361 (w1169, w1158, IN56[2], w1170, w1171);
  FullAdder U362 (w1171, w1160, IN57[1], w1172, w1173);
  FullAdder U363 (w1173, w1161, IN58[0], w1174, w1175);
  HalfAdder U364 (w1164, IN53[6], Out1[53], w1177);
  FullAdder U365 (w1177, w1166, IN54[5], w1178, w1179);
  FullAdder U366 (w1179, w1168, IN55[4], w1180, w1181);
  FullAdder U367 (w1181, w1170, IN56[3], w1182, w1183);
  FullAdder U368 (w1183, w1172, IN57[2], w1184, w1185);
  FullAdder U369 (w1185, w1174, IN58[1], w1186, w1187);
  FullAdder U370 (w1187, w1175, IN59[0], w1188, w1189);
  HalfAdder U371 (w1178, IN54[6], Out1[54], w1191);
  FullAdder U372 (w1191, w1180, IN55[5], w1192, w1193);
  FullAdder U373 (w1193, w1182, IN56[4], w1194, w1195);
  FullAdder U374 (w1195, w1184, IN57[3], w1196, w1197);
  FullAdder U375 (w1197, w1186, IN58[2], w1198, w1199);
  FullAdder U376 (w1199, w1188, IN59[1], w1200, w1201);
  FullAdder U377 (w1201, w1189, IN60[0], w1202, w1203);
  HalfAdder U378 (w1192, IN55[6], Out1[55], w1205);
  FullAdder U379 (w1205, w1194, IN56[5], Out1[56], w1207);
  FullAdder U380 (w1207, w1196, IN57[4], Out1[57], w1209);
  FullAdder U381 (w1209, w1198, IN58[3], Out1[58], w1211);
  FullAdder U382 (w1211, w1200, IN59[2], Out1[59], w1213);
  FullAdder U383 (w1213, w1202, IN60[1], Out1[60], w1215);
  FullAdder U384 (w1215, w1203, IN61[0], Out1[61], Out1[62]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN8[7];
  assign Out2[1] = IN9[7];
  assign Out2[2] = IN10[7];
  assign Out2[3] = IN11[7];
  assign Out2[4] = IN12[7];
  assign Out2[5] = IN13[7];
  assign Out2[6] = IN14[7];
  assign Out2[7] = IN15[7];
  assign Out2[8] = IN16[7];
  assign Out2[9] = IN17[7];
  assign Out2[10] = IN18[7];
  assign Out2[11] = IN19[7];
  assign Out2[12] = IN20[7];
  assign Out2[13] = IN21[7];
  assign Out2[14] = IN22[7];
  assign Out2[15] = IN23[7];
  assign Out2[16] = IN24[7];
  assign Out2[17] = IN25[7];
  assign Out2[18] = IN26[7];
  assign Out2[19] = IN27[7];
  assign Out2[20] = IN28[7];
  assign Out2[21] = IN29[7];
  assign Out2[22] = IN30[7];
  assign Out2[23] = IN31[7];
  assign Out2[24] = IN32[7];
  assign Out2[25] = IN33[7];
  assign Out2[26] = IN34[7];
  assign Out2[27] = IN35[7];
  assign Out2[28] = IN36[7];
  assign Out2[29] = IN37[7];
  assign Out2[30] = IN38[7];
  assign Out2[31] = IN39[7];
  assign Out2[32] = IN40[7];
  assign Out2[33] = IN41[7];
  assign Out2[34] = IN42[7];
  assign Out2[35] = IN43[7];
  assign Out2[36] = IN44[7];
  assign Out2[37] = IN45[7];
  assign Out2[38] = IN46[7];
  assign Out2[39] = IN47[7];
  assign Out2[40] = IN48[7];
  assign Out2[41] = IN49[7];
  assign Out2[42] = IN50[7];
  assign Out2[43] = IN51[7];
  assign Out2[44] = IN52[7];
  assign Out2[45] = IN53[7];
  assign Out2[46] = IN54[7];
  assign Out2[47] = IN55[7];
  assign Out2[48] = IN56[6];
  assign Out2[49] = IN57[5];
  assign Out2[50] = IN58[4];
  assign Out2[51] = IN59[3];
  assign Out2[52] = IN60[2];
  assign Out2[53] = IN61[1];
  assign Out2[54] = IN62[0];

endmodule
module RC_55_55(IN1, IN2, Out);
  input [54:0] IN1;
  input [54:0] IN2;
  output [55:0] Out;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w111);
  FullAdder U1 (IN1[1], IN2[1], w111, Out[1], w113);
  FullAdder U2 (IN1[2], IN2[2], w113, Out[2], w115);
  FullAdder U3 (IN1[3], IN2[3], w115, Out[3], w117);
  FullAdder U4 (IN1[4], IN2[4], w117, Out[4], w119);
  FullAdder U5 (IN1[5], IN2[5], w119, Out[5], w121);
  FullAdder U6 (IN1[6], IN2[6], w121, Out[6], w123);
  FullAdder U7 (IN1[7], IN2[7], w123, Out[7], w125);
  FullAdder U8 (IN1[8], IN2[8], w125, Out[8], w127);
  FullAdder U9 (IN1[9], IN2[9], w127, Out[9], w129);
  FullAdder U10 (IN1[10], IN2[10], w129, Out[10], w131);
  FullAdder U11 (IN1[11], IN2[11], w131, Out[11], w133);
  FullAdder U12 (IN1[12], IN2[12], w133, Out[12], w135);
  FullAdder U13 (IN1[13], IN2[13], w135, Out[13], w137);
  FullAdder U14 (IN1[14], IN2[14], w137, Out[14], w139);
  FullAdder U15 (IN1[15], IN2[15], w139, Out[15], w141);
  FullAdder U16 (IN1[16], IN2[16], w141, Out[16], w143);
  FullAdder U17 (IN1[17], IN2[17], w143, Out[17], w145);
  FullAdder U18 (IN1[18], IN2[18], w145, Out[18], w147);
  FullAdder U19 (IN1[19], IN2[19], w147, Out[19], w149);
  FullAdder U20 (IN1[20], IN2[20], w149, Out[20], w151);
  FullAdder U21 (IN1[21], IN2[21], w151, Out[21], w153);
  FullAdder U22 (IN1[22], IN2[22], w153, Out[22], w155);
  FullAdder U23 (IN1[23], IN2[23], w155, Out[23], w157);
  FullAdder U24 (IN1[24], IN2[24], w157, Out[24], w159);
  FullAdder U25 (IN1[25], IN2[25], w159, Out[25], w161);
  FullAdder U26 (IN1[26], IN2[26], w161, Out[26], w163);
  FullAdder U27 (IN1[27], IN2[27], w163, Out[27], w165);
  FullAdder U28 (IN1[28], IN2[28], w165, Out[28], w167);
  FullAdder U29 (IN1[29], IN2[29], w167, Out[29], w169);
  FullAdder U30 (IN1[30], IN2[30], w169, Out[30], w171);
  FullAdder U31 (IN1[31], IN2[31], w171, Out[31], w173);
  FullAdder U32 (IN1[32], IN2[32], w173, Out[32], w175);
  FullAdder U33 (IN1[33], IN2[33], w175, Out[33], w177);
  FullAdder U34 (IN1[34], IN2[34], w177, Out[34], w179);
  FullAdder U35 (IN1[35], IN2[35], w179, Out[35], w181);
  FullAdder U36 (IN1[36], IN2[36], w181, Out[36], w183);
  FullAdder U37 (IN1[37], IN2[37], w183, Out[37], w185);
  FullAdder U38 (IN1[38], IN2[38], w185, Out[38], w187);
  FullAdder U39 (IN1[39], IN2[39], w187, Out[39], w189);
  FullAdder U40 (IN1[40], IN2[40], w189, Out[40], w191);
  FullAdder U41 (IN1[41], IN2[41], w191, Out[41], w193);
  FullAdder U42 (IN1[42], IN2[42], w193, Out[42], w195);
  FullAdder U43 (IN1[43], IN2[43], w195, Out[43], w197);
  FullAdder U44 (IN1[44], IN2[44], w197, Out[44], w199);
  FullAdder U45 (IN1[45], IN2[45], w199, Out[45], w201);
  FullAdder U46 (IN1[46], IN2[46], w201, Out[46], w203);
  FullAdder U47 (IN1[47], IN2[47], w203, Out[47], w205);
  FullAdder U48 (IN1[48], IN2[48], w205, Out[48], w207);
  FullAdder U49 (IN1[49], IN2[49], w207, Out[49], w209);
  FullAdder U50 (IN1[50], IN2[50], w209, Out[50], w211);
  FullAdder U51 (IN1[51], IN2[51], w211, Out[51], w213);
  FullAdder U52 (IN1[52], IN2[52], w213, Out[52], w215);
  FullAdder U53 (IN1[53], IN2[53], w215, Out[53], w217);
  FullAdder U54 (IN1[54], IN2[54], w217, Out[54], Out[55]);

endmodule
module NR_8_56(IN1, IN2, Out);
  input [7:0] IN1;
  input [55:0] IN2;
  output [63:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [7:0] P8;
  wire [7:0] P9;
  wire [7:0] P10;
  wire [7:0] P11;
  wire [7:0] P12;
  wire [7:0] P13;
  wire [7:0] P14;
  wire [7:0] P15;
  wire [7:0] P16;
  wire [7:0] P17;
  wire [7:0] P18;
  wire [7:0] P19;
  wire [7:0] P20;
  wire [7:0] P21;
  wire [7:0] P22;
  wire [7:0] P23;
  wire [7:0] P24;
  wire [7:0] P25;
  wire [7:0] P26;
  wire [7:0] P27;
  wire [7:0] P28;
  wire [7:0] P29;
  wire [7:0] P30;
  wire [7:0] P31;
  wire [7:0] P32;
  wire [7:0] P33;
  wire [7:0] P34;
  wire [7:0] P35;
  wire [7:0] P36;
  wire [7:0] P37;
  wire [7:0] P38;
  wire [7:0] P39;
  wire [7:0] P40;
  wire [7:0] P41;
  wire [7:0] P42;
  wire [7:0] P43;
  wire [7:0] P44;
  wire [7:0] P45;
  wire [7:0] P46;
  wire [7:0] P47;
  wire [7:0] P48;
  wire [7:0] P49;
  wire [7:0] P50;
  wire [7:0] P51;
  wire [7:0] P52;
  wire [7:0] P53;
  wire [7:0] P54;
  wire [7:0] P55;
  wire [6:0] P56;
  wire [5:0] P57;
  wire [4:0] P58;
  wire [3:0] P59;
  wire [2:0] P60;
  wire [1:0] P61;
  wire [0:0] P62;
  wire [62:0] R1;
  wire [54:0] R2;
  wire [63:0] aOut;
  U_SP_8_56 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, R1, R2);
  RC_55_55 S2 (R1[62:8], R2, aOut[63:8]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign Out = aOut[63:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
