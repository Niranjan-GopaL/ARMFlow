
module NR_43_1(
    input [42:0]IN1,
    input [0:0]IN2,
    output [42:0]Out
);
    assign Out = IN2;
endmodule
