
module NR_51_1(
    input [50:0]IN1,
    input [0:0]IN2,
    output [50:0]Out
);
    assign Out = IN2;
endmodule
