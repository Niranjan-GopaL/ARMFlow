
module customAdder60_0(
    input [59 : 0] A,
    input [59 : 0] B,
    output [60 : 0] Sum
);

    assign Sum = A+B;

endmodule
