
module NR_59_1(
    input [58:0]IN1,
    input [0:0]IN2,
    output [58:0]Out
);
    assign Out = IN2;
endmodule
