//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 14
  second input length: 60
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_14_60(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72);
  input [13:0] IN1;
  input [59:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [13:0] P14;
  output [13:0] P15;
  output [13:0] P16;
  output [13:0] P17;
  output [13:0] P18;
  output [13:0] P19;
  output [13:0] P20;
  output [13:0] P21;
  output [13:0] P22;
  output [13:0] P23;
  output [13:0] P24;
  output [13:0] P25;
  output [13:0] P26;
  output [13:0] P27;
  output [13:0] P28;
  output [13:0] P29;
  output [13:0] P30;
  output [13:0] P31;
  output [13:0] P32;
  output [13:0] P33;
  output [13:0] P34;
  output [13:0] P35;
  output [13:0] P36;
  output [13:0] P37;
  output [13:0] P38;
  output [13:0] P39;
  output [13:0] P40;
  output [13:0] P41;
  output [13:0] P42;
  output [13:0] P43;
  output [13:0] P44;
  output [13:0] P45;
  output [13:0] P46;
  output [13:0] P47;
  output [13:0] P48;
  output [13:0] P49;
  output [13:0] P50;
  output [13:0] P51;
  output [13:0] P52;
  output [13:0] P53;
  output [13:0] P54;
  output [13:0] P55;
  output [13:0] P56;
  output [13:0] P57;
  output [13:0] P58;
  output [13:0] P59;
  output [12:0] P60;
  output [11:0] P61;
  output [10:0] P62;
  output [9:0] P63;
  output [8:0] P64;
  output [7:0] P65;
  output [6:0] P66;
  output [5:0] P67;
  output [4:0] P68;
  output [3:0] P69;
  output [2:0] P70;
  output [1:0] P71;
  output [0:0] P72;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P59[0] = IN1[0]&IN2[59];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[1] = IN1[1]&IN2[58];
  assign P60[0] = IN1[1]&IN2[59];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[2] = IN1[2]&IN2[57];
  assign P60[1] = IN1[2]&IN2[58];
  assign P61[0] = IN1[2]&IN2[59];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[3] = IN1[3]&IN2[56];
  assign P60[2] = IN1[3]&IN2[57];
  assign P61[1] = IN1[3]&IN2[58];
  assign P62[0] = IN1[3]&IN2[59];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[4] = IN1[4]&IN2[55];
  assign P60[3] = IN1[4]&IN2[56];
  assign P61[2] = IN1[4]&IN2[57];
  assign P62[1] = IN1[4]&IN2[58];
  assign P63[0] = IN1[4]&IN2[59];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[5] = IN1[5]&IN2[54];
  assign P60[4] = IN1[5]&IN2[55];
  assign P61[3] = IN1[5]&IN2[56];
  assign P62[2] = IN1[5]&IN2[57];
  assign P63[1] = IN1[5]&IN2[58];
  assign P64[0] = IN1[5]&IN2[59];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[6] = IN1[6]&IN2[53];
  assign P60[5] = IN1[6]&IN2[54];
  assign P61[4] = IN1[6]&IN2[55];
  assign P62[3] = IN1[6]&IN2[56];
  assign P63[2] = IN1[6]&IN2[57];
  assign P64[1] = IN1[6]&IN2[58];
  assign P65[0] = IN1[6]&IN2[59];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[7] = IN1[7]&IN2[47];
  assign P55[7] = IN1[7]&IN2[48];
  assign P56[7] = IN1[7]&IN2[49];
  assign P57[7] = IN1[7]&IN2[50];
  assign P58[7] = IN1[7]&IN2[51];
  assign P59[7] = IN1[7]&IN2[52];
  assign P60[6] = IN1[7]&IN2[53];
  assign P61[5] = IN1[7]&IN2[54];
  assign P62[4] = IN1[7]&IN2[55];
  assign P63[3] = IN1[7]&IN2[56];
  assign P64[2] = IN1[7]&IN2[57];
  assign P65[1] = IN1[7]&IN2[58];
  assign P66[0] = IN1[7]&IN2[59];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[8] = IN1[8]&IN2[45];
  assign P54[8] = IN1[8]&IN2[46];
  assign P55[8] = IN1[8]&IN2[47];
  assign P56[8] = IN1[8]&IN2[48];
  assign P57[8] = IN1[8]&IN2[49];
  assign P58[8] = IN1[8]&IN2[50];
  assign P59[8] = IN1[8]&IN2[51];
  assign P60[7] = IN1[8]&IN2[52];
  assign P61[6] = IN1[8]&IN2[53];
  assign P62[5] = IN1[8]&IN2[54];
  assign P63[4] = IN1[8]&IN2[55];
  assign P64[3] = IN1[8]&IN2[56];
  assign P65[2] = IN1[8]&IN2[57];
  assign P66[1] = IN1[8]&IN2[58];
  assign P67[0] = IN1[8]&IN2[59];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[9] = IN1[9]&IN2[44];
  assign P54[9] = IN1[9]&IN2[45];
  assign P55[9] = IN1[9]&IN2[46];
  assign P56[9] = IN1[9]&IN2[47];
  assign P57[9] = IN1[9]&IN2[48];
  assign P58[9] = IN1[9]&IN2[49];
  assign P59[9] = IN1[9]&IN2[50];
  assign P60[8] = IN1[9]&IN2[51];
  assign P61[7] = IN1[9]&IN2[52];
  assign P62[6] = IN1[9]&IN2[53];
  assign P63[5] = IN1[9]&IN2[54];
  assign P64[4] = IN1[9]&IN2[55];
  assign P65[3] = IN1[9]&IN2[56];
  assign P66[2] = IN1[9]&IN2[57];
  assign P67[1] = IN1[9]&IN2[58];
  assign P68[0] = IN1[9]&IN2[59];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[10] = IN1[10]&IN2[39];
  assign P50[10] = IN1[10]&IN2[40];
  assign P51[10] = IN1[10]&IN2[41];
  assign P52[10] = IN1[10]&IN2[42];
  assign P53[10] = IN1[10]&IN2[43];
  assign P54[10] = IN1[10]&IN2[44];
  assign P55[10] = IN1[10]&IN2[45];
  assign P56[10] = IN1[10]&IN2[46];
  assign P57[10] = IN1[10]&IN2[47];
  assign P58[10] = IN1[10]&IN2[48];
  assign P59[10] = IN1[10]&IN2[49];
  assign P60[9] = IN1[10]&IN2[50];
  assign P61[8] = IN1[10]&IN2[51];
  assign P62[7] = IN1[10]&IN2[52];
  assign P63[6] = IN1[10]&IN2[53];
  assign P64[5] = IN1[10]&IN2[54];
  assign P65[4] = IN1[10]&IN2[55];
  assign P66[3] = IN1[10]&IN2[56];
  assign P67[2] = IN1[10]&IN2[57];
  assign P68[1] = IN1[10]&IN2[58];
  assign P69[0] = IN1[10]&IN2[59];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[11] = IN1[11]&IN2[38];
  assign P50[11] = IN1[11]&IN2[39];
  assign P51[11] = IN1[11]&IN2[40];
  assign P52[11] = IN1[11]&IN2[41];
  assign P53[11] = IN1[11]&IN2[42];
  assign P54[11] = IN1[11]&IN2[43];
  assign P55[11] = IN1[11]&IN2[44];
  assign P56[11] = IN1[11]&IN2[45];
  assign P57[11] = IN1[11]&IN2[46];
  assign P58[11] = IN1[11]&IN2[47];
  assign P59[11] = IN1[11]&IN2[48];
  assign P60[10] = IN1[11]&IN2[49];
  assign P61[9] = IN1[11]&IN2[50];
  assign P62[8] = IN1[11]&IN2[51];
  assign P63[7] = IN1[11]&IN2[52];
  assign P64[6] = IN1[11]&IN2[53];
  assign P65[5] = IN1[11]&IN2[54];
  assign P66[4] = IN1[11]&IN2[55];
  assign P67[3] = IN1[11]&IN2[56];
  assign P68[2] = IN1[11]&IN2[57];
  assign P69[1] = IN1[11]&IN2[58];
  assign P70[0] = IN1[11]&IN2[59];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[12] = IN1[12]&IN2[37];
  assign P50[12] = IN1[12]&IN2[38];
  assign P51[12] = IN1[12]&IN2[39];
  assign P52[12] = IN1[12]&IN2[40];
  assign P53[12] = IN1[12]&IN2[41];
  assign P54[12] = IN1[12]&IN2[42];
  assign P55[12] = IN1[12]&IN2[43];
  assign P56[12] = IN1[12]&IN2[44];
  assign P57[12] = IN1[12]&IN2[45];
  assign P58[12] = IN1[12]&IN2[46];
  assign P59[12] = IN1[12]&IN2[47];
  assign P60[11] = IN1[12]&IN2[48];
  assign P61[10] = IN1[12]&IN2[49];
  assign P62[9] = IN1[12]&IN2[50];
  assign P63[8] = IN1[12]&IN2[51];
  assign P64[7] = IN1[12]&IN2[52];
  assign P65[6] = IN1[12]&IN2[53];
  assign P66[5] = IN1[12]&IN2[54];
  assign P67[4] = IN1[12]&IN2[55];
  assign P68[3] = IN1[12]&IN2[56];
  assign P69[2] = IN1[12]&IN2[57];
  assign P70[1] = IN1[12]&IN2[58];
  assign P71[0] = IN1[12]&IN2[59];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[13] = IN1[13]&IN2[36];
  assign P50[13] = IN1[13]&IN2[37];
  assign P51[13] = IN1[13]&IN2[38];
  assign P52[13] = IN1[13]&IN2[39];
  assign P53[13] = IN1[13]&IN2[40];
  assign P54[13] = IN1[13]&IN2[41];
  assign P55[13] = IN1[13]&IN2[42];
  assign P56[13] = IN1[13]&IN2[43];
  assign P57[13] = IN1[13]&IN2[44];
  assign P58[13] = IN1[13]&IN2[45];
  assign P59[13] = IN1[13]&IN2[46];
  assign P60[12] = IN1[13]&IN2[47];
  assign P61[11] = IN1[13]&IN2[48];
  assign P62[10] = IN1[13]&IN2[49];
  assign P63[9] = IN1[13]&IN2[50];
  assign P64[8] = IN1[13]&IN2[51];
  assign P65[7] = IN1[13]&IN2[52];
  assign P66[6] = IN1[13]&IN2[53];
  assign P67[5] = IN1[13]&IN2[54];
  assign P68[4] = IN1[13]&IN2[55];
  assign P69[3] = IN1[13]&IN2[56];
  assign P70[2] = IN1[13]&IN2[57];
  assign P71[1] = IN1[13]&IN2[58];
  assign P72[0] = IN1[13]&IN2[59];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [13:0] IN14;
  input [13:0] IN15;
  input [13:0] IN16;
  input [13:0] IN17;
  input [13:0] IN18;
  input [13:0] IN19;
  input [13:0] IN20;
  input [13:0] IN21;
  input [13:0] IN22;
  input [13:0] IN23;
  input [13:0] IN24;
  input [13:0] IN25;
  input [13:0] IN26;
  input [13:0] IN27;
  input [13:0] IN28;
  input [13:0] IN29;
  input [13:0] IN30;
  input [13:0] IN31;
  input [13:0] IN32;
  input [13:0] IN33;
  input [13:0] IN34;
  input [13:0] IN35;
  input [13:0] IN36;
  input [13:0] IN37;
  input [13:0] IN38;
  input [13:0] IN39;
  input [13:0] IN40;
  input [13:0] IN41;
  input [13:0] IN42;
  input [13:0] IN43;
  input [13:0] IN44;
  input [13:0] IN45;
  input [13:0] IN46;
  input [13:0] IN47;
  input [13:0] IN48;
  input [13:0] IN49;
  input [13:0] IN50;
  input [13:0] IN51;
  input [13:0] IN52;
  input [13:0] IN53;
  input [13:0] IN54;
  input [13:0] IN55;
  input [13:0] IN56;
  input [13:0] IN57;
  input [13:0] IN58;
  input [13:0] IN59;
  input [12:0] IN60;
  input [11:0] IN61;
  input [10:0] IN62;
  input [9:0] IN63;
  input [8:0] IN64;
  input [7:0] IN65;
  input [6:0] IN66;
  input [5:0] IN67;
  input [4:0] IN68;
  input [3:0] IN69;
  input [2:0] IN70;
  input [1:0] IN71;
  input [0:0] IN72;
  output [72:0] Out1;
  output [58:0] Out2;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1231;
  wire w1232;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1257;
  wire w1258;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1283;
  wire w1284;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1309;
  wire w1310;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1335;
  wire w1336;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1361;
  wire w1362;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1387;
  wire w1388;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1413;
  wire w1414;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1439;
  wire w1440;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1465;
  wire w1466;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1491;
  wire w1492;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1517;
  wire w1518;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1543;
  wire w1544;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1569;
  wire w1570;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1595;
  wire w1596;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1621;
  wire w1622;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1647;
  wire w1648;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1673;
  wire w1674;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1699;
  wire w1700;
  wire w1701;
  wire w1702;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1725;
  wire w1726;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1751;
  wire w1752;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1777;
  wire w1778;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1803;
  wire w1804;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1829;
  wire w1830;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1855;
  wire w1856;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1881;
  wire w1882;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1907;
  wire w1908;
  wire w1909;
  wire w1910;
  wire w1911;
  wire w1912;
  wire w1913;
  wire w1914;
  wire w1915;
  wire w1916;
  wire w1917;
  wire w1918;
  wire w1919;
  wire w1920;
  wire w1921;
  wire w1922;
  wire w1923;
  wire w1924;
  wire w1925;
  wire w1926;
  wire w1927;
  wire w1928;
  wire w1929;
  wire w1930;
  wire w1931;
  wire w1933;
  wire w1934;
  wire w1935;
  wire w1936;
  wire w1937;
  wire w1938;
  wire w1939;
  wire w1940;
  wire w1941;
  wire w1942;
  wire w1943;
  wire w1944;
  wire w1945;
  wire w1946;
  wire w1947;
  wire w1948;
  wire w1949;
  wire w1950;
  wire w1951;
  wire w1952;
  wire w1953;
  wire w1954;
  wire w1955;
  wire w1956;
  wire w1957;
  wire w1959;
  wire w1960;
  wire w1961;
  wire w1962;
  wire w1963;
  wire w1964;
  wire w1965;
  wire w1966;
  wire w1967;
  wire w1968;
  wire w1969;
  wire w1970;
  wire w1971;
  wire w1972;
  wire w1973;
  wire w1974;
  wire w1975;
  wire w1976;
  wire w1977;
  wire w1978;
  wire w1979;
  wire w1980;
  wire w1981;
  wire w1982;
  wire w1983;
  wire w1985;
  wire w1986;
  wire w1987;
  wire w1988;
  wire w1989;
  wire w1990;
  wire w1991;
  wire w1992;
  wire w1993;
  wire w1994;
  wire w1995;
  wire w1996;
  wire w1997;
  wire w1998;
  wire w1999;
  wire w2000;
  wire w2001;
  wire w2002;
  wire w2003;
  wire w2004;
  wire w2005;
  wire w2006;
  wire w2007;
  wire w2008;
  wire w2009;
  wire w2011;
  wire w2012;
  wire w2013;
  wire w2014;
  wire w2015;
  wire w2016;
  wire w2017;
  wire w2018;
  wire w2019;
  wire w2020;
  wire w2021;
  wire w2022;
  wire w2023;
  wire w2024;
  wire w2025;
  wire w2026;
  wire w2027;
  wire w2028;
  wire w2029;
  wire w2030;
  wire w2031;
  wire w2032;
  wire w2033;
  wire w2034;
  wire w2035;
  wire w2037;
  wire w2038;
  wire w2039;
  wire w2040;
  wire w2041;
  wire w2042;
  wire w2043;
  wire w2044;
  wire w2045;
  wire w2046;
  wire w2047;
  wire w2048;
  wire w2049;
  wire w2050;
  wire w2051;
  wire w2052;
  wire w2053;
  wire w2054;
  wire w2055;
  wire w2056;
  wire w2057;
  wire w2058;
  wire w2059;
  wire w2060;
  wire w2061;
  wire w2063;
  wire w2064;
  wire w2065;
  wire w2066;
  wire w2067;
  wire w2068;
  wire w2069;
  wire w2070;
  wire w2071;
  wire w2072;
  wire w2073;
  wire w2074;
  wire w2075;
  wire w2076;
  wire w2077;
  wire w2078;
  wire w2079;
  wire w2080;
  wire w2081;
  wire w2082;
  wire w2083;
  wire w2084;
  wire w2085;
  wire w2086;
  wire w2087;
  wire w2089;
  wire w2090;
  wire w2091;
  wire w2092;
  wire w2093;
  wire w2094;
  wire w2095;
  wire w2096;
  wire w2097;
  wire w2098;
  wire w2099;
  wire w2100;
  wire w2101;
  wire w2102;
  wire w2103;
  wire w2104;
  wire w2105;
  wire w2106;
  wire w2107;
  wire w2108;
  wire w2109;
  wire w2110;
  wire w2111;
  wire w2112;
  wire w2113;
  wire w2115;
  wire w2116;
  wire w2117;
  wire w2118;
  wire w2119;
  wire w2120;
  wire w2121;
  wire w2122;
  wire w2123;
  wire w2124;
  wire w2125;
  wire w2126;
  wire w2127;
  wire w2128;
  wire w2129;
  wire w2130;
  wire w2131;
  wire w2132;
  wire w2133;
  wire w2134;
  wire w2135;
  wire w2136;
  wire w2137;
  wire w2138;
  wire w2139;
  wire w2141;
  wire w2142;
  wire w2143;
  wire w2144;
  wire w2145;
  wire w2146;
  wire w2147;
  wire w2148;
  wire w2149;
  wire w2150;
  wire w2151;
  wire w2152;
  wire w2153;
  wire w2154;
  wire w2155;
  wire w2156;
  wire w2157;
  wire w2158;
  wire w2159;
  wire w2160;
  wire w2161;
  wire w2162;
  wire w2163;
  wire w2164;
  wire w2165;
  wire w2167;
  wire w2168;
  wire w2169;
  wire w2170;
  wire w2171;
  wire w2172;
  wire w2173;
  wire w2174;
  wire w2175;
  wire w2176;
  wire w2177;
  wire w2178;
  wire w2179;
  wire w2180;
  wire w2181;
  wire w2182;
  wire w2183;
  wire w2184;
  wire w2185;
  wire w2186;
  wire w2187;
  wire w2188;
  wire w2189;
  wire w2190;
  wire w2191;
  wire w2193;
  wire w2194;
  wire w2195;
  wire w2196;
  wire w2197;
  wire w2198;
  wire w2199;
  wire w2200;
  wire w2201;
  wire w2202;
  wire w2203;
  wire w2204;
  wire w2205;
  wire w2206;
  wire w2207;
  wire w2208;
  wire w2209;
  wire w2210;
  wire w2211;
  wire w2212;
  wire w2213;
  wire w2214;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2294;
  wire w2295;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2349;
  wire w2351;
  wire w2353;
  wire w2355;
  wire w2357;
  wire w2359;
  wire w2361;
  wire w2363;
  wire w2365;
  wire w2367;
  wire w2369;
  wire w2371;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w841);
  FullAdder U1 (w841, IN2[0], IN2[1], w842, w843);
  FullAdder U2 (w843, IN3[0], IN3[1], w844, w845);
  FullAdder U3 (w845, IN4[0], IN4[1], w846, w847);
  FullAdder U4 (w847, IN5[0], IN5[1], w848, w849);
  FullAdder U5 (w849, IN6[0], IN6[1], w850, w851);
  FullAdder U6 (w851, IN7[0], IN7[1], w852, w853);
  FullAdder U7 (w853, IN8[0], IN8[1], w854, w855);
  FullAdder U8 (w855, IN9[0], IN9[1], w856, w857);
  FullAdder U9 (w857, IN10[0], IN10[1], w858, w859);
  FullAdder U10 (w859, IN11[0], IN11[1], w860, w861);
  FullAdder U11 (w861, IN12[0], IN12[1], w862, w863);
  FullAdder U12 (w863, IN13[0], IN13[1], w864, w865);
  HalfAdder U13 (w842, IN2[2], Out1[2], w867);
  FullAdder U14 (w867, w844, IN3[2], w868, w869);
  FullAdder U15 (w869, w846, IN4[2], w870, w871);
  FullAdder U16 (w871, w848, IN5[2], w872, w873);
  FullAdder U17 (w873, w850, IN6[2], w874, w875);
  FullAdder U18 (w875, w852, IN7[2], w876, w877);
  FullAdder U19 (w877, w854, IN8[2], w878, w879);
  FullAdder U20 (w879, w856, IN9[2], w880, w881);
  FullAdder U21 (w881, w858, IN10[2], w882, w883);
  FullAdder U22 (w883, w860, IN11[2], w884, w885);
  FullAdder U23 (w885, w862, IN12[2], w886, w887);
  FullAdder U24 (w887, w864, IN13[2], w888, w889);
  FullAdder U25 (w889, w865, IN14[0], w890, w891);
  HalfAdder U26 (w868, IN3[3], Out1[3], w893);
  FullAdder U27 (w893, w870, IN4[3], w894, w895);
  FullAdder U28 (w895, w872, IN5[3], w896, w897);
  FullAdder U29 (w897, w874, IN6[3], w898, w899);
  FullAdder U30 (w899, w876, IN7[3], w900, w901);
  FullAdder U31 (w901, w878, IN8[3], w902, w903);
  FullAdder U32 (w903, w880, IN9[3], w904, w905);
  FullAdder U33 (w905, w882, IN10[3], w906, w907);
  FullAdder U34 (w907, w884, IN11[3], w908, w909);
  FullAdder U35 (w909, w886, IN12[3], w910, w911);
  FullAdder U36 (w911, w888, IN13[3], w912, w913);
  FullAdder U37 (w913, w890, IN14[1], w914, w915);
  FullAdder U38 (w915, w891, IN15[0], w916, w917);
  HalfAdder U39 (w894, IN4[4], Out1[4], w919);
  FullAdder U40 (w919, w896, IN5[4], w920, w921);
  FullAdder U41 (w921, w898, IN6[4], w922, w923);
  FullAdder U42 (w923, w900, IN7[4], w924, w925);
  FullAdder U43 (w925, w902, IN8[4], w926, w927);
  FullAdder U44 (w927, w904, IN9[4], w928, w929);
  FullAdder U45 (w929, w906, IN10[4], w930, w931);
  FullAdder U46 (w931, w908, IN11[4], w932, w933);
  FullAdder U47 (w933, w910, IN12[4], w934, w935);
  FullAdder U48 (w935, w912, IN13[4], w936, w937);
  FullAdder U49 (w937, w914, IN14[2], w938, w939);
  FullAdder U50 (w939, w916, IN15[1], w940, w941);
  FullAdder U51 (w941, w917, IN16[0], w942, w943);
  HalfAdder U52 (w920, IN5[5], Out1[5], w945);
  FullAdder U53 (w945, w922, IN6[5], w946, w947);
  FullAdder U54 (w947, w924, IN7[5], w948, w949);
  FullAdder U55 (w949, w926, IN8[5], w950, w951);
  FullAdder U56 (w951, w928, IN9[5], w952, w953);
  FullAdder U57 (w953, w930, IN10[5], w954, w955);
  FullAdder U58 (w955, w932, IN11[5], w956, w957);
  FullAdder U59 (w957, w934, IN12[5], w958, w959);
  FullAdder U60 (w959, w936, IN13[5], w960, w961);
  FullAdder U61 (w961, w938, IN14[3], w962, w963);
  FullAdder U62 (w963, w940, IN15[2], w964, w965);
  FullAdder U63 (w965, w942, IN16[1], w966, w967);
  FullAdder U64 (w967, w943, IN17[0], w968, w969);
  HalfAdder U65 (w946, IN6[6], Out1[6], w971);
  FullAdder U66 (w971, w948, IN7[6], w972, w973);
  FullAdder U67 (w973, w950, IN8[6], w974, w975);
  FullAdder U68 (w975, w952, IN9[6], w976, w977);
  FullAdder U69 (w977, w954, IN10[6], w978, w979);
  FullAdder U70 (w979, w956, IN11[6], w980, w981);
  FullAdder U71 (w981, w958, IN12[6], w982, w983);
  FullAdder U72 (w983, w960, IN13[6], w984, w985);
  FullAdder U73 (w985, w962, IN14[4], w986, w987);
  FullAdder U74 (w987, w964, IN15[3], w988, w989);
  FullAdder U75 (w989, w966, IN16[2], w990, w991);
  FullAdder U76 (w991, w968, IN17[1], w992, w993);
  FullAdder U77 (w993, w969, IN18[0], w994, w995);
  HalfAdder U78 (w972, IN7[7], Out1[7], w997);
  FullAdder U79 (w997, w974, IN8[7], w998, w999);
  FullAdder U80 (w999, w976, IN9[7], w1000, w1001);
  FullAdder U81 (w1001, w978, IN10[7], w1002, w1003);
  FullAdder U82 (w1003, w980, IN11[7], w1004, w1005);
  FullAdder U83 (w1005, w982, IN12[7], w1006, w1007);
  FullAdder U84 (w1007, w984, IN13[7], w1008, w1009);
  FullAdder U85 (w1009, w986, IN14[5], w1010, w1011);
  FullAdder U86 (w1011, w988, IN15[4], w1012, w1013);
  FullAdder U87 (w1013, w990, IN16[3], w1014, w1015);
  FullAdder U88 (w1015, w992, IN17[2], w1016, w1017);
  FullAdder U89 (w1017, w994, IN18[1], w1018, w1019);
  FullAdder U90 (w1019, w995, IN19[0], w1020, w1021);
  HalfAdder U91 (w998, IN8[8], Out1[8], w1023);
  FullAdder U92 (w1023, w1000, IN9[8], w1024, w1025);
  FullAdder U93 (w1025, w1002, IN10[8], w1026, w1027);
  FullAdder U94 (w1027, w1004, IN11[8], w1028, w1029);
  FullAdder U95 (w1029, w1006, IN12[8], w1030, w1031);
  FullAdder U96 (w1031, w1008, IN13[8], w1032, w1033);
  FullAdder U97 (w1033, w1010, IN14[6], w1034, w1035);
  FullAdder U98 (w1035, w1012, IN15[5], w1036, w1037);
  FullAdder U99 (w1037, w1014, IN16[4], w1038, w1039);
  FullAdder U100 (w1039, w1016, IN17[3], w1040, w1041);
  FullAdder U101 (w1041, w1018, IN18[2], w1042, w1043);
  FullAdder U102 (w1043, w1020, IN19[1], w1044, w1045);
  FullAdder U103 (w1045, w1021, IN20[0], w1046, w1047);
  HalfAdder U104 (w1024, IN9[9], Out1[9], w1049);
  FullAdder U105 (w1049, w1026, IN10[9], w1050, w1051);
  FullAdder U106 (w1051, w1028, IN11[9], w1052, w1053);
  FullAdder U107 (w1053, w1030, IN12[9], w1054, w1055);
  FullAdder U108 (w1055, w1032, IN13[9], w1056, w1057);
  FullAdder U109 (w1057, w1034, IN14[7], w1058, w1059);
  FullAdder U110 (w1059, w1036, IN15[6], w1060, w1061);
  FullAdder U111 (w1061, w1038, IN16[5], w1062, w1063);
  FullAdder U112 (w1063, w1040, IN17[4], w1064, w1065);
  FullAdder U113 (w1065, w1042, IN18[3], w1066, w1067);
  FullAdder U114 (w1067, w1044, IN19[2], w1068, w1069);
  FullAdder U115 (w1069, w1046, IN20[1], w1070, w1071);
  FullAdder U116 (w1071, w1047, IN21[0], w1072, w1073);
  HalfAdder U117 (w1050, IN10[10], Out1[10], w1075);
  FullAdder U118 (w1075, w1052, IN11[10], w1076, w1077);
  FullAdder U119 (w1077, w1054, IN12[10], w1078, w1079);
  FullAdder U120 (w1079, w1056, IN13[10], w1080, w1081);
  FullAdder U121 (w1081, w1058, IN14[8], w1082, w1083);
  FullAdder U122 (w1083, w1060, IN15[7], w1084, w1085);
  FullAdder U123 (w1085, w1062, IN16[6], w1086, w1087);
  FullAdder U124 (w1087, w1064, IN17[5], w1088, w1089);
  FullAdder U125 (w1089, w1066, IN18[4], w1090, w1091);
  FullAdder U126 (w1091, w1068, IN19[3], w1092, w1093);
  FullAdder U127 (w1093, w1070, IN20[2], w1094, w1095);
  FullAdder U128 (w1095, w1072, IN21[1], w1096, w1097);
  FullAdder U129 (w1097, w1073, IN22[0], w1098, w1099);
  HalfAdder U130 (w1076, IN11[11], Out1[11], w1101);
  FullAdder U131 (w1101, w1078, IN12[11], w1102, w1103);
  FullAdder U132 (w1103, w1080, IN13[11], w1104, w1105);
  FullAdder U133 (w1105, w1082, IN14[9], w1106, w1107);
  FullAdder U134 (w1107, w1084, IN15[8], w1108, w1109);
  FullAdder U135 (w1109, w1086, IN16[7], w1110, w1111);
  FullAdder U136 (w1111, w1088, IN17[6], w1112, w1113);
  FullAdder U137 (w1113, w1090, IN18[5], w1114, w1115);
  FullAdder U138 (w1115, w1092, IN19[4], w1116, w1117);
  FullAdder U139 (w1117, w1094, IN20[3], w1118, w1119);
  FullAdder U140 (w1119, w1096, IN21[2], w1120, w1121);
  FullAdder U141 (w1121, w1098, IN22[1], w1122, w1123);
  FullAdder U142 (w1123, w1099, IN23[0], w1124, w1125);
  HalfAdder U143 (w1102, IN12[12], Out1[12], w1127);
  FullAdder U144 (w1127, w1104, IN13[12], w1128, w1129);
  FullAdder U145 (w1129, w1106, IN14[10], w1130, w1131);
  FullAdder U146 (w1131, w1108, IN15[9], w1132, w1133);
  FullAdder U147 (w1133, w1110, IN16[8], w1134, w1135);
  FullAdder U148 (w1135, w1112, IN17[7], w1136, w1137);
  FullAdder U149 (w1137, w1114, IN18[6], w1138, w1139);
  FullAdder U150 (w1139, w1116, IN19[5], w1140, w1141);
  FullAdder U151 (w1141, w1118, IN20[4], w1142, w1143);
  FullAdder U152 (w1143, w1120, IN21[3], w1144, w1145);
  FullAdder U153 (w1145, w1122, IN22[2], w1146, w1147);
  FullAdder U154 (w1147, w1124, IN23[1], w1148, w1149);
  FullAdder U155 (w1149, w1125, IN24[0], w1150, w1151);
  HalfAdder U156 (w1128, IN13[13], Out1[13], w1153);
  FullAdder U157 (w1153, w1130, IN14[11], w1154, w1155);
  FullAdder U158 (w1155, w1132, IN15[10], w1156, w1157);
  FullAdder U159 (w1157, w1134, IN16[9], w1158, w1159);
  FullAdder U160 (w1159, w1136, IN17[8], w1160, w1161);
  FullAdder U161 (w1161, w1138, IN18[7], w1162, w1163);
  FullAdder U162 (w1163, w1140, IN19[6], w1164, w1165);
  FullAdder U163 (w1165, w1142, IN20[5], w1166, w1167);
  FullAdder U164 (w1167, w1144, IN21[4], w1168, w1169);
  FullAdder U165 (w1169, w1146, IN22[3], w1170, w1171);
  FullAdder U166 (w1171, w1148, IN23[2], w1172, w1173);
  FullAdder U167 (w1173, w1150, IN24[1], w1174, w1175);
  FullAdder U168 (w1175, w1151, IN25[0], w1176, w1177);
  HalfAdder U169 (w1154, IN14[12], Out1[14], w1179);
  FullAdder U170 (w1179, w1156, IN15[11], w1180, w1181);
  FullAdder U171 (w1181, w1158, IN16[10], w1182, w1183);
  FullAdder U172 (w1183, w1160, IN17[9], w1184, w1185);
  FullAdder U173 (w1185, w1162, IN18[8], w1186, w1187);
  FullAdder U174 (w1187, w1164, IN19[7], w1188, w1189);
  FullAdder U175 (w1189, w1166, IN20[6], w1190, w1191);
  FullAdder U176 (w1191, w1168, IN21[5], w1192, w1193);
  FullAdder U177 (w1193, w1170, IN22[4], w1194, w1195);
  FullAdder U178 (w1195, w1172, IN23[3], w1196, w1197);
  FullAdder U179 (w1197, w1174, IN24[2], w1198, w1199);
  FullAdder U180 (w1199, w1176, IN25[1], w1200, w1201);
  FullAdder U181 (w1201, w1177, IN26[0], w1202, w1203);
  HalfAdder U182 (w1180, IN15[12], Out1[15], w1205);
  FullAdder U183 (w1205, w1182, IN16[11], w1206, w1207);
  FullAdder U184 (w1207, w1184, IN17[10], w1208, w1209);
  FullAdder U185 (w1209, w1186, IN18[9], w1210, w1211);
  FullAdder U186 (w1211, w1188, IN19[8], w1212, w1213);
  FullAdder U187 (w1213, w1190, IN20[7], w1214, w1215);
  FullAdder U188 (w1215, w1192, IN21[6], w1216, w1217);
  FullAdder U189 (w1217, w1194, IN22[5], w1218, w1219);
  FullAdder U190 (w1219, w1196, IN23[4], w1220, w1221);
  FullAdder U191 (w1221, w1198, IN24[3], w1222, w1223);
  FullAdder U192 (w1223, w1200, IN25[2], w1224, w1225);
  FullAdder U193 (w1225, w1202, IN26[1], w1226, w1227);
  FullAdder U194 (w1227, w1203, IN27[0], w1228, w1229);
  HalfAdder U195 (w1206, IN16[12], Out1[16], w1231);
  FullAdder U196 (w1231, w1208, IN17[11], w1232, w1233);
  FullAdder U197 (w1233, w1210, IN18[10], w1234, w1235);
  FullAdder U198 (w1235, w1212, IN19[9], w1236, w1237);
  FullAdder U199 (w1237, w1214, IN20[8], w1238, w1239);
  FullAdder U200 (w1239, w1216, IN21[7], w1240, w1241);
  FullAdder U201 (w1241, w1218, IN22[6], w1242, w1243);
  FullAdder U202 (w1243, w1220, IN23[5], w1244, w1245);
  FullAdder U203 (w1245, w1222, IN24[4], w1246, w1247);
  FullAdder U204 (w1247, w1224, IN25[3], w1248, w1249);
  FullAdder U205 (w1249, w1226, IN26[2], w1250, w1251);
  FullAdder U206 (w1251, w1228, IN27[1], w1252, w1253);
  FullAdder U207 (w1253, w1229, IN28[0], w1254, w1255);
  HalfAdder U208 (w1232, IN17[12], Out1[17], w1257);
  FullAdder U209 (w1257, w1234, IN18[11], w1258, w1259);
  FullAdder U210 (w1259, w1236, IN19[10], w1260, w1261);
  FullAdder U211 (w1261, w1238, IN20[9], w1262, w1263);
  FullAdder U212 (w1263, w1240, IN21[8], w1264, w1265);
  FullAdder U213 (w1265, w1242, IN22[7], w1266, w1267);
  FullAdder U214 (w1267, w1244, IN23[6], w1268, w1269);
  FullAdder U215 (w1269, w1246, IN24[5], w1270, w1271);
  FullAdder U216 (w1271, w1248, IN25[4], w1272, w1273);
  FullAdder U217 (w1273, w1250, IN26[3], w1274, w1275);
  FullAdder U218 (w1275, w1252, IN27[2], w1276, w1277);
  FullAdder U219 (w1277, w1254, IN28[1], w1278, w1279);
  FullAdder U220 (w1279, w1255, IN29[0], w1280, w1281);
  HalfAdder U221 (w1258, IN18[12], Out1[18], w1283);
  FullAdder U222 (w1283, w1260, IN19[11], w1284, w1285);
  FullAdder U223 (w1285, w1262, IN20[10], w1286, w1287);
  FullAdder U224 (w1287, w1264, IN21[9], w1288, w1289);
  FullAdder U225 (w1289, w1266, IN22[8], w1290, w1291);
  FullAdder U226 (w1291, w1268, IN23[7], w1292, w1293);
  FullAdder U227 (w1293, w1270, IN24[6], w1294, w1295);
  FullAdder U228 (w1295, w1272, IN25[5], w1296, w1297);
  FullAdder U229 (w1297, w1274, IN26[4], w1298, w1299);
  FullAdder U230 (w1299, w1276, IN27[3], w1300, w1301);
  FullAdder U231 (w1301, w1278, IN28[2], w1302, w1303);
  FullAdder U232 (w1303, w1280, IN29[1], w1304, w1305);
  FullAdder U233 (w1305, w1281, IN30[0], w1306, w1307);
  HalfAdder U234 (w1284, IN19[12], Out1[19], w1309);
  FullAdder U235 (w1309, w1286, IN20[11], w1310, w1311);
  FullAdder U236 (w1311, w1288, IN21[10], w1312, w1313);
  FullAdder U237 (w1313, w1290, IN22[9], w1314, w1315);
  FullAdder U238 (w1315, w1292, IN23[8], w1316, w1317);
  FullAdder U239 (w1317, w1294, IN24[7], w1318, w1319);
  FullAdder U240 (w1319, w1296, IN25[6], w1320, w1321);
  FullAdder U241 (w1321, w1298, IN26[5], w1322, w1323);
  FullAdder U242 (w1323, w1300, IN27[4], w1324, w1325);
  FullAdder U243 (w1325, w1302, IN28[3], w1326, w1327);
  FullAdder U244 (w1327, w1304, IN29[2], w1328, w1329);
  FullAdder U245 (w1329, w1306, IN30[1], w1330, w1331);
  FullAdder U246 (w1331, w1307, IN31[0], w1332, w1333);
  HalfAdder U247 (w1310, IN20[12], Out1[20], w1335);
  FullAdder U248 (w1335, w1312, IN21[11], w1336, w1337);
  FullAdder U249 (w1337, w1314, IN22[10], w1338, w1339);
  FullAdder U250 (w1339, w1316, IN23[9], w1340, w1341);
  FullAdder U251 (w1341, w1318, IN24[8], w1342, w1343);
  FullAdder U252 (w1343, w1320, IN25[7], w1344, w1345);
  FullAdder U253 (w1345, w1322, IN26[6], w1346, w1347);
  FullAdder U254 (w1347, w1324, IN27[5], w1348, w1349);
  FullAdder U255 (w1349, w1326, IN28[4], w1350, w1351);
  FullAdder U256 (w1351, w1328, IN29[3], w1352, w1353);
  FullAdder U257 (w1353, w1330, IN30[2], w1354, w1355);
  FullAdder U258 (w1355, w1332, IN31[1], w1356, w1357);
  FullAdder U259 (w1357, w1333, IN32[0], w1358, w1359);
  HalfAdder U260 (w1336, IN21[12], Out1[21], w1361);
  FullAdder U261 (w1361, w1338, IN22[11], w1362, w1363);
  FullAdder U262 (w1363, w1340, IN23[10], w1364, w1365);
  FullAdder U263 (w1365, w1342, IN24[9], w1366, w1367);
  FullAdder U264 (w1367, w1344, IN25[8], w1368, w1369);
  FullAdder U265 (w1369, w1346, IN26[7], w1370, w1371);
  FullAdder U266 (w1371, w1348, IN27[6], w1372, w1373);
  FullAdder U267 (w1373, w1350, IN28[5], w1374, w1375);
  FullAdder U268 (w1375, w1352, IN29[4], w1376, w1377);
  FullAdder U269 (w1377, w1354, IN30[3], w1378, w1379);
  FullAdder U270 (w1379, w1356, IN31[2], w1380, w1381);
  FullAdder U271 (w1381, w1358, IN32[1], w1382, w1383);
  FullAdder U272 (w1383, w1359, IN33[0], w1384, w1385);
  HalfAdder U273 (w1362, IN22[12], Out1[22], w1387);
  FullAdder U274 (w1387, w1364, IN23[11], w1388, w1389);
  FullAdder U275 (w1389, w1366, IN24[10], w1390, w1391);
  FullAdder U276 (w1391, w1368, IN25[9], w1392, w1393);
  FullAdder U277 (w1393, w1370, IN26[8], w1394, w1395);
  FullAdder U278 (w1395, w1372, IN27[7], w1396, w1397);
  FullAdder U279 (w1397, w1374, IN28[6], w1398, w1399);
  FullAdder U280 (w1399, w1376, IN29[5], w1400, w1401);
  FullAdder U281 (w1401, w1378, IN30[4], w1402, w1403);
  FullAdder U282 (w1403, w1380, IN31[3], w1404, w1405);
  FullAdder U283 (w1405, w1382, IN32[2], w1406, w1407);
  FullAdder U284 (w1407, w1384, IN33[1], w1408, w1409);
  FullAdder U285 (w1409, w1385, IN34[0], w1410, w1411);
  HalfAdder U286 (w1388, IN23[12], Out1[23], w1413);
  FullAdder U287 (w1413, w1390, IN24[11], w1414, w1415);
  FullAdder U288 (w1415, w1392, IN25[10], w1416, w1417);
  FullAdder U289 (w1417, w1394, IN26[9], w1418, w1419);
  FullAdder U290 (w1419, w1396, IN27[8], w1420, w1421);
  FullAdder U291 (w1421, w1398, IN28[7], w1422, w1423);
  FullAdder U292 (w1423, w1400, IN29[6], w1424, w1425);
  FullAdder U293 (w1425, w1402, IN30[5], w1426, w1427);
  FullAdder U294 (w1427, w1404, IN31[4], w1428, w1429);
  FullAdder U295 (w1429, w1406, IN32[3], w1430, w1431);
  FullAdder U296 (w1431, w1408, IN33[2], w1432, w1433);
  FullAdder U297 (w1433, w1410, IN34[1], w1434, w1435);
  FullAdder U298 (w1435, w1411, IN35[0], w1436, w1437);
  HalfAdder U299 (w1414, IN24[12], Out1[24], w1439);
  FullAdder U300 (w1439, w1416, IN25[11], w1440, w1441);
  FullAdder U301 (w1441, w1418, IN26[10], w1442, w1443);
  FullAdder U302 (w1443, w1420, IN27[9], w1444, w1445);
  FullAdder U303 (w1445, w1422, IN28[8], w1446, w1447);
  FullAdder U304 (w1447, w1424, IN29[7], w1448, w1449);
  FullAdder U305 (w1449, w1426, IN30[6], w1450, w1451);
  FullAdder U306 (w1451, w1428, IN31[5], w1452, w1453);
  FullAdder U307 (w1453, w1430, IN32[4], w1454, w1455);
  FullAdder U308 (w1455, w1432, IN33[3], w1456, w1457);
  FullAdder U309 (w1457, w1434, IN34[2], w1458, w1459);
  FullAdder U310 (w1459, w1436, IN35[1], w1460, w1461);
  FullAdder U311 (w1461, w1437, IN36[0], w1462, w1463);
  HalfAdder U312 (w1440, IN25[12], Out1[25], w1465);
  FullAdder U313 (w1465, w1442, IN26[11], w1466, w1467);
  FullAdder U314 (w1467, w1444, IN27[10], w1468, w1469);
  FullAdder U315 (w1469, w1446, IN28[9], w1470, w1471);
  FullAdder U316 (w1471, w1448, IN29[8], w1472, w1473);
  FullAdder U317 (w1473, w1450, IN30[7], w1474, w1475);
  FullAdder U318 (w1475, w1452, IN31[6], w1476, w1477);
  FullAdder U319 (w1477, w1454, IN32[5], w1478, w1479);
  FullAdder U320 (w1479, w1456, IN33[4], w1480, w1481);
  FullAdder U321 (w1481, w1458, IN34[3], w1482, w1483);
  FullAdder U322 (w1483, w1460, IN35[2], w1484, w1485);
  FullAdder U323 (w1485, w1462, IN36[1], w1486, w1487);
  FullAdder U324 (w1487, w1463, IN37[0], w1488, w1489);
  HalfAdder U325 (w1466, IN26[12], Out1[26], w1491);
  FullAdder U326 (w1491, w1468, IN27[11], w1492, w1493);
  FullAdder U327 (w1493, w1470, IN28[10], w1494, w1495);
  FullAdder U328 (w1495, w1472, IN29[9], w1496, w1497);
  FullAdder U329 (w1497, w1474, IN30[8], w1498, w1499);
  FullAdder U330 (w1499, w1476, IN31[7], w1500, w1501);
  FullAdder U331 (w1501, w1478, IN32[6], w1502, w1503);
  FullAdder U332 (w1503, w1480, IN33[5], w1504, w1505);
  FullAdder U333 (w1505, w1482, IN34[4], w1506, w1507);
  FullAdder U334 (w1507, w1484, IN35[3], w1508, w1509);
  FullAdder U335 (w1509, w1486, IN36[2], w1510, w1511);
  FullAdder U336 (w1511, w1488, IN37[1], w1512, w1513);
  FullAdder U337 (w1513, w1489, IN38[0], w1514, w1515);
  HalfAdder U338 (w1492, IN27[12], Out1[27], w1517);
  FullAdder U339 (w1517, w1494, IN28[11], w1518, w1519);
  FullAdder U340 (w1519, w1496, IN29[10], w1520, w1521);
  FullAdder U341 (w1521, w1498, IN30[9], w1522, w1523);
  FullAdder U342 (w1523, w1500, IN31[8], w1524, w1525);
  FullAdder U343 (w1525, w1502, IN32[7], w1526, w1527);
  FullAdder U344 (w1527, w1504, IN33[6], w1528, w1529);
  FullAdder U345 (w1529, w1506, IN34[5], w1530, w1531);
  FullAdder U346 (w1531, w1508, IN35[4], w1532, w1533);
  FullAdder U347 (w1533, w1510, IN36[3], w1534, w1535);
  FullAdder U348 (w1535, w1512, IN37[2], w1536, w1537);
  FullAdder U349 (w1537, w1514, IN38[1], w1538, w1539);
  FullAdder U350 (w1539, w1515, IN39[0], w1540, w1541);
  HalfAdder U351 (w1518, IN28[12], Out1[28], w1543);
  FullAdder U352 (w1543, w1520, IN29[11], w1544, w1545);
  FullAdder U353 (w1545, w1522, IN30[10], w1546, w1547);
  FullAdder U354 (w1547, w1524, IN31[9], w1548, w1549);
  FullAdder U355 (w1549, w1526, IN32[8], w1550, w1551);
  FullAdder U356 (w1551, w1528, IN33[7], w1552, w1553);
  FullAdder U357 (w1553, w1530, IN34[6], w1554, w1555);
  FullAdder U358 (w1555, w1532, IN35[5], w1556, w1557);
  FullAdder U359 (w1557, w1534, IN36[4], w1558, w1559);
  FullAdder U360 (w1559, w1536, IN37[3], w1560, w1561);
  FullAdder U361 (w1561, w1538, IN38[2], w1562, w1563);
  FullAdder U362 (w1563, w1540, IN39[1], w1564, w1565);
  FullAdder U363 (w1565, w1541, IN40[0], w1566, w1567);
  HalfAdder U364 (w1544, IN29[12], Out1[29], w1569);
  FullAdder U365 (w1569, w1546, IN30[11], w1570, w1571);
  FullAdder U366 (w1571, w1548, IN31[10], w1572, w1573);
  FullAdder U367 (w1573, w1550, IN32[9], w1574, w1575);
  FullAdder U368 (w1575, w1552, IN33[8], w1576, w1577);
  FullAdder U369 (w1577, w1554, IN34[7], w1578, w1579);
  FullAdder U370 (w1579, w1556, IN35[6], w1580, w1581);
  FullAdder U371 (w1581, w1558, IN36[5], w1582, w1583);
  FullAdder U372 (w1583, w1560, IN37[4], w1584, w1585);
  FullAdder U373 (w1585, w1562, IN38[3], w1586, w1587);
  FullAdder U374 (w1587, w1564, IN39[2], w1588, w1589);
  FullAdder U375 (w1589, w1566, IN40[1], w1590, w1591);
  FullAdder U376 (w1591, w1567, IN41[0], w1592, w1593);
  HalfAdder U377 (w1570, IN30[12], Out1[30], w1595);
  FullAdder U378 (w1595, w1572, IN31[11], w1596, w1597);
  FullAdder U379 (w1597, w1574, IN32[10], w1598, w1599);
  FullAdder U380 (w1599, w1576, IN33[9], w1600, w1601);
  FullAdder U381 (w1601, w1578, IN34[8], w1602, w1603);
  FullAdder U382 (w1603, w1580, IN35[7], w1604, w1605);
  FullAdder U383 (w1605, w1582, IN36[6], w1606, w1607);
  FullAdder U384 (w1607, w1584, IN37[5], w1608, w1609);
  FullAdder U385 (w1609, w1586, IN38[4], w1610, w1611);
  FullAdder U386 (w1611, w1588, IN39[3], w1612, w1613);
  FullAdder U387 (w1613, w1590, IN40[2], w1614, w1615);
  FullAdder U388 (w1615, w1592, IN41[1], w1616, w1617);
  FullAdder U389 (w1617, w1593, IN42[0], w1618, w1619);
  HalfAdder U390 (w1596, IN31[12], Out1[31], w1621);
  FullAdder U391 (w1621, w1598, IN32[11], w1622, w1623);
  FullAdder U392 (w1623, w1600, IN33[10], w1624, w1625);
  FullAdder U393 (w1625, w1602, IN34[9], w1626, w1627);
  FullAdder U394 (w1627, w1604, IN35[8], w1628, w1629);
  FullAdder U395 (w1629, w1606, IN36[7], w1630, w1631);
  FullAdder U396 (w1631, w1608, IN37[6], w1632, w1633);
  FullAdder U397 (w1633, w1610, IN38[5], w1634, w1635);
  FullAdder U398 (w1635, w1612, IN39[4], w1636, w1637);
  FullAdder U399 (w1637, w1614, IN40[3], w1638, w1639);
  FullAdder U400 (w1639, w1616, IN41[2], w1640, w1641);
  FullAdder U401 (w1641, w1618, IN42[1], w1642, w1643);
  FullAdder U402 (w1643, w1619, IN43[0], w1644, w1645);
  HalfAdder U403 (w1622, IN32[12], Out1[32], w1647);
  FullAdder U404 (w1647, w1624, IN33[11], w1648, w1649);
  FullAdder U405 (w1649, w1626, IN34[10], w1650, w1651);
  FullAdder U406 (w1651, w1628, IN35[9], w1652, w1653);
  FullAdder U407 (w1653, w1630, IN36[8], w1654, w1655);
  FullAdder U408 (w1655, w1632, IN37[7], w1656, w1657);
  FullAdder U409 (w1657, w1634, IN38[6], w1658, w1659);
  FullAdder U410 (w1659, w1636, IN39[5], w1660, w1661);
  FullAdder U411 (w1661, w1638, IN40[4], w1662, w1663);
  FullAdder U412 (w1663, w1640, IN41[3], w1664, w1665);
  FullAdder U413 (w1665, w1642, IN42[2], w1666, w1667);
  FullAdder U414 (w1667, w1644, IN43[1], w1668, w1669);
  FullAdder U415 (w1669, w1645, IN44[0], w1670, w1671);
  HalfAdder U416 (w1648, IN33[12], Out1[33], w1673);
  FullAdder U417 (w1673, w1650, IN34[11], w1674, w1675);
  FullAdder U418 (w1675, w1652, IN35[10], w1676, w1677);
  FullAdder U419 (w1677, w1654, IN36[9], w1678, w1679);
  FullAdder U420 (w1679, w1656, IN37[8], w1680, w1681);
  FullAdder U421 (w1681, w1658, IN38[7], w1682, w1683);
  FullAdder U422 (w1683, w1660, IN39[6], w1684, w1685);
  FullAdder U423 (w1685, w1662, IN40[5], w1686, w1687);
  FullAdder U424 (w1687, w1664, IN41[4], w1688, w1689);
  FullAdder U425 (w1689, w1666, IN42[3], w1690, w1691);
  FullAdder U426 (w1691, w1668, IN43[2], w1692, w1693);
  FullAdder U427 (w1693, w1670, IN44[1], w1694, w1695);
  FullAdder U428 (w1695, w1671, IN45[0], w1696, w1697);
  HalfAdder U429 (w1674, IN34[12], Out1[34], w1699);
  FullAdder U430 (w1699, w1676, IN35[11], w1700, w1701);
  FullAdder U431 (w1701, w1678, IN36[10], w1702, w1703);
  FullAdder U432 (w1703, w1680, IN37[9], w1704, w1705);
  FullAdder U433 (w1705, w1682, IN38[8], w1706, w1707);
  FullAdder U434 (w1707, w1684, IN39[7], w1708, w1709);
  FullAdder U435 (w1709, w1686, IN40[6], w1710, w1711);
  FullAdder U436 (w1711, w1688, IN41[5], w1712, w1713);
  FullAdder U437 (w1713, w1690, IN42[4], w1714, w1715);
  FullAdder U438 (w1715, w1692, IN43[3], w1716, w1717);
  FullAdder U439 (w1717, w1694, IN44[2], w1718, w1719);
  FullAdder U440 (w1719, w1696, IN45[1], w1720, w1721);
  FullAdder U441 (w1721, w1697, IN46[0], w1722, w1723);
  HalfAdder U442 (w1700, IN35[12], Out1[35], w1725);
  FullAdder U443 (w1725, w1702, IN36[11], w1726, w1727);
  FullAdder U444 (w1727, w1704, IN37[10], w1728, w1729);
  FullAdder U445 (w1729, w1706, IN38[9], w1730, w1731);
  FullAdder U446 (w1731, w1708, IN39[8], w1732, w1733);
  FullAdder U447 (w1733, w1710, IN40[7], w1734, w1735);
  FullAdder U448 (w1735, w1712, IN41[6], w1736, w1737);
  FullAdder U449 (w1737, w1714, IN42[5], w1738, w1739);
  FullAdder U450 (w1739, w1716, IN43[4], w1740, w1741);
  FullAdder U451 (w1741, w1718, IN44[3], w1742, w1743);
  FullAdder U452 (w1743, w1720, IN45[2], w1744, w1745);
  FullAdder U453 (w1745, w1722, IN46[1], w1746, w1747);
  FullAdder U454 (w1747, w1723, IN47[0], w1748, w1749);
  HalfAdder U455 (w1726, IN36[12], Out1[36], w1751);
  FullAdder U456 (w1751, w1728, IN37[11], w1752, w1753);
  FullAdder U457 (w1753, w1730, IN38[10], w1754, w1755);
  FullAdder U458 (w1755, w1732, IN39[9], w1756, w1757);
  FullAdder U459 (w1757, w1734, IN40[8], w1758, w1759);
  FullAdder U460 (w1759, w1736, IN41[7], w1760, w1761);
  FullAdder U461 (w1761, w1738, IN42[6], w1762, w1763);
  FullAdder U462 (w1763, w1740, IN43[5], w1764, w1765);
  FullAdder U463 (w1765, w1742, IN44[4], w1766, w1767);
  FullAdder U464 (w1767, w1744, IN45[3], w1768, w1769);
  FullAdder U465 (w1769, w1746, IN46[2], w1770, w1771);
  FullAdder U466 (w1771, w1748, IN47[1], w1772, w1773);
  FullAdder U467 (w1773, w1749, IN48[0], w1774, w1775);
  HalfAdder U468 (w1752, IN37[12], Out1[37], w1777);
  FullAdder U469 (w1777, w1754, IN38[11], w1778, w1779);
  FullAdder U470 (w1779, w1756, IN39[10], w1780, w1781);
  FullAdder U471 (w1781, w1758, IN40[9], w1782, w1783);
  FullAdder U472 (w1783, w1760, IN41[8], w1784, w1785);
  FullAdder U473 (w1785, w1762, IN42[7], w1786, w1787);
  FullAdder U474 (w1787, w1764, IN43[6], w1788, w1789);
  FullAdder U475 (w1789, w1766, IN44[5], w1790, w1791);
  FullAdder U476 (w1791, w1768, IN45[4], w1792, w1793);
  FullAdder U477 (w1793, w1770, IN46[3], w1794, w1795);
  FullAdder U478 (w1795, w1772, IN47[2], w1796, w1797);
  FullAdder U479 (w1797, w1774, IN48[1], w1798, w1799);
  FullAdder U480 (w1799, w1775, IN49[0], w1800, w1801);
  HalfAdder U481 (w1778, IN38[12], Out1[38], w1803);
  FullAdder U482 (w1803, w1780, IN39[11], w1804, w1805);
  FullAdder U483 (w1805, w1782, IN40[10], w1806, w1807);
  FullAdder U484 (w1807, w1784, IN41[9], w1808, w1809);
  FullAdder U485 (w1809, w1786, IN42[8], w1810, w1811);
  FullAdder U486 (w1811, w1788, IN43[7], w1812, w1813);
  FullAdder U487 (w1813, w1790, IN44[6], w1814, w1815);
  FullAdder U488 (w1815, w1792, IN45[5], w1816, w1817);
  FullAdder U489 (w1817, w1794, IN46[4], w1818, w1819);
  FullAdder U490 (w1819, w1796, IN47[3], w1820, w1821);
  FullAdder U491 (w1821, w1798, IN48[2], w1822, w1823);
  FullAdder U492 (w1823, w1800, IN49[1], w1824, w1825);
  FullAdder U493 (w1825, w1801, IN50[0], w1826, w1827);
  HalfAdder U494 (w1804, IN39[12], Out1[39], w1829);
  FullAdder U495 (w1829, w1806, IN40[11], w1830, w1831);
  FullAdder U496 (w1831, w1808, IN41[10], w1832, w1833);
  FullAdder U497 (w1833, w1810, IN42[9], w1834, w1835);
  FullAdder U498 (w1835, w1812, IN43[8], w1836, w1837);
  FullAdder U499 (w1837, w1814, IN44[7], w1838, w1839);
  FullAdder U500 (w1839, w1816, IN45[6], w1840, w1841);
  FullAdder U501 (w1841, w1818, IN46[5], w1842, w1843);
  FullAdder U502 (w1843, w1820, IN47[4], w1844, w1845);
  FullAdder U503 (w1845, w1822, IN48[3], w1846, w1847);
  FullAdder U504 (w1847, w1824, IN49[2], w1848, w1849);
  FullAdder U505 (w1849, w1826, IN50[1], w1850, w1851);
  FullAdder U506 (w1851, w1827, IN51[0], w1852, w1853);
  HalfAdder U507 (w1830, IN40[12], Out1[40], w1855);
  FullAdder U508 (w1855, w1832, IN41[11], w1856, w1857);
  FullAdder U509 (w1857, w1834, IN42[10], w1858, w1859);
  FullAdder U510 (w1859, w1836, IN43[9], w1860, w1861);
  FullAdder U511 (w1861, w1838, IN44[8], w1862, w1863);
  FullAdder U512 (w1863, w1840, IN45[7], w1864, w1865);
  FullAdder U513 (w1865, w1842, IN46[6], w1866, w1867);
  FullAdder U514 (w1867, w1844, IN47[5], w1868, w1869);
  FullAdder U515 (w1869, w1846, IN48[4], w1870, w1871);
  FullAdder U516 (w1871, w1848, IN49[3], w1872, w1873);
  FullAdder U517 (w1873, w1850, IN50[2], w1874, w1875);
  FullAdder U518 (w1875, w1852, IN51[1], w1876, w1877);
  FullAdder U519 (w1877, w1853, IN52[0], w1878, w1879);
  HalfAdder U520 (w1856, IN41[12], Out1[41], w1881);
  FullAdder U521 (w1881, w1858, IN42[11], w1882, w1883);
  FullAdder U522 (w1883, w1860, IN43[10], w1884, w1885);
  FullAdder U523 (w1885, w1862, IN44[9], w1886, w1887);
  FullAdder U524 (w1887, w1864, IN45[8], w1888, w1889);
  FullAdder U525 (w1889, w1866, IN46[7], w1890, w1891);
  FullAdder U526 (w1891, w1868, IN47[6], w1892, w1893);
  FullAdder U527 (w1893, w1870, IN48[5], w1894, w1895);
  FullAdder U528 (w1895, w1872, IN49[4], w1896, w1897);
  FullAdder U529 (w1897, w1874, IN50[3], w1898, w1899);
  FullAdder U530 (w1899, w1876, IN51[2], w1900, w1901);
  FullAdder U531 (w1901, w1878, IN52[1], w1902, w1903);
  FullAdder U532 (w1903, w1879, IN53[0], w1904, w1905);
  HalfAdder U533 (w1882, IN42[12], Out1[42], w1907);
  FullAdder U534 (w1907, w1884, IN43[11], w1908, w1909);
  FullAdder U535 (w1909, w1886, IN44[10], w1910, w1911);
  FullAdder U536 (w1911, w1888, IN45[9], w1912, w1913);
  FullAdder U537 (w1913, w1890, IN46[8], w1914, w1915);
  FullAdder U538 (w1915, w1892, IN47[7], w1916, w1917);
  FullAdder U539 (w1917, w1894, IN48[6], w1918, w1919);
  FullAdder U540 (w1919, w1896, IN49[5], w1920, w1921);
  FullAdder U541 (w1921, w1898, IN50[4], w1922, w1923);
  FullAdder U542 (w1923, w1900, IN51[3], w1924, w1925);
  FullAdder U543 (w1925, w1902, IN52[2], w1926, w1927);
  FullAdder U544 (w1927, w1904, IN53[1], w1928, w1929);
  FullAdder U545 (w1929, w1905, IN54[0], w1930, w1931);
  HalfAdder U546 (w1908, IN43[12], Out1[43], w1933);
  FullAdder U547 (w1933, w1910, IN44[11], w1934, w1935);
  FullAdder U548 (w1935, w1912, IN45[10], w1936, w1937);
  FullAdder U549 (w1937, w1914, IN46[9], w1938, w1939);
  FullAdder U550 (w1939, w1916, IN47[8], w1940, w1941);
  FullAdder U551 (w1941, w1918, IN48[7], w1942, w1943);
  FullAdder U552 (w1943, w1920, IN49[6], w1944, w1945);
  FullAdder U553 (w1945, w1922, IN50[5], w1946, w1947);
  FullAdder U554 (w1947, w1924, IN51[4], w1948, w1949);
  FullAdder U555 (w1949, w1926, IN52[3], w1950, w1951);
  FullAdder U556 (w1951, w1928, IN53[2], w1952, w1953);
  FullAdder U557 (w1953, w1930, IN54[1], w1954, w1955);
  FullAdder U558 (w1955, w1931, IN55[0], w1956, w1957);
  HalfAdder U559 (w1934, IN44[12], Out1[44], w1959);
  FullAdder U560 (w1959, w1936, IN45[11], w1960, w1961);
  FullAdder U561 (w1961, w1938, IN46[10], w1962, w1963);
  FullAdder U562 (w1963, w1940, IN47[9], w1964, w1965);
  FullAdder U563 (w1965, w1942, IN48[8], w1966, w1967);
  FullAdder U564 (w1967, w1944, IN49[7], w1968, w1969);
  FullAdder U565 (w1969, w1946, IN50[6], w1970, w1971);
  FullAdder U566 (w1971, w1948, IN51[5], w1972, w1973);
  FullAdder U567 (w1973, w1950, IN52[4], w1974, w1975);
  FullAdder U568 (w1975, w1952, IN53[3], w1976, w1977);
  FullAdder U569 (w1977, w1954, IN54[2], w1978, w1979);
  FullAdder U570 (w1979, w1956, IN55[1], w1980, w1981);
  FullAdder U571 (w1981, w1957, IN56[0], w1982, w1983);
  HalfAdder U572 (w1960, IN45[12], Out1[45], w1985);
  FullAdder U573 (w1985, w1962, IN46[11], w1986, w1987);
  FullAdder U574 (w1987, w1964, IN47[10], w1988, w1989);
  FullAdder U575 (w1989, w1966, IN48[9], w1990, w1991);
  FullAdder U576 (w1991, w1968, IN49[8], w1992, w1993);
  FullAdder U577 (w1993, w1970, IN50[7], w1994, w1995);
  FullAdder U578 (w1995, w1972, IN51[6], w1996, w1997);
  FullAdder U579 (w1997, w1974, IN52[5], w1998, w1999);
  FullAdder U580 (w1999, w1976, IN53[4], w2000, w2001);
  FullAdder U581 (w2001, w1978, IN54[3], w2002, w2003);
  FullAdder U582 (w2003, w1980, IN55[2], w2004, w2005);
  FullAdder U583 (w2005, w1982, IN56[1], w2006, w2007);
  FullAdder U584 (w2007, w1983, IN57[0], w2008, w2009);
  HalfAdder U585 (w1986, IN46[12], Out1[46], w2011);
  FullAdder U586 (w2011, w1988, IN47[11], w2012, w2013);
  FullAdder U587 (w2013, w1990, IN48[10], w2014, w2015);
  FullAdder U588 (w2015, w1992, IN49[9], w2016, w2017);
  FullAdder U589 (w2017, w1994, IN50[8], w2018, w2019);
  FullAdder U590 (w2019, w1996, IN51[7], w2020, w2021);
  FullAdder U591 (w2021, w1998, IN52[6], w2022, w2023);
  FullAdder U592 (w2023, w2000, IN53[5], w2024, w2025);
  FullAdder U593 (w2025, w2002, IN54[4], w2026, w2027);
  FullAdder U594 (w2027, w2004, IN55[3], w2028, w2029);
  FullAdder U595 (w2029, w2006, IN56[2], w2030, w2031);
  FullAdder U596 (w2031, w2008, IN57[1], w2032, w2033);
  FullAdder U597 (w2033, w2009, IN58[0], w2034, w2035);
  HalfAdder U598 (w2012, IN47[12], Out1[47], w2037);
  FullAdder U599 (w2037, w2014, IN48[11], w2038, w2039);
  FullAdder U600 (w2039, w2016, IN49[10], w2040, w2041);
  FullAdder U601 (w2041, w2018, IN50[9], w2042, w2043);
  FullAdder U602 (w2043, w2020, IN51[8], w2044, w2045);
  FullAdder U603 (w2045, w2022, IN52[7], w2046, w2047);
  FullAdder U604 (w2047, w2024, IN53[6], w2048, w2049);
  FullAdder U605 (w2049, w2026, IN54[5], w2050, w2051);
  FullAdder U606 (w2051, w2028, IN55[4], w2052, w2053);
  FullAdder U607 (w2053, w2030, IN56[3], w2054, w2055);
  FullAdder U608 (w2055, w2032, IN57[2], w2056, w2057);
  FullAdder U609 (w2057, w2034, IN58[1], w2058, w2059);
  FullAdder U610 (w2059, w2035, IN59[0], w2060, w2061);
  HalfAdder U611 (w2038, IN48[12], Out1[48], w2063);
  FullAdder U612 (w2063, w2040, IN49[11], w2064, w2065);
  FullAdder U613 (w2065, w2042, IN50[10], w2066, w2067);
  FullAdder U614 (w2067, w2044, IN51[9], w2068, w2069);
  FullAdder U615 (w2069, w2046, IN52[8], w2070, w2071);
  FullAdder U616 (w2071, w2048, IN53[7], w2072, w2073);
  FullAdder U617 (w2073, w2050, IN54[6], w2074, w2075);
  FullAdder U618 (w2075, w2052, IN55[5], w2076, w2077);
  FullAdder U619 (w2077, w2054, IN56[4], w2078, w2079);
  FullAdder U620 (w2079, w2056, IN57[3], w2080, w2081);
  FullAdder U621 (w2081, w2058, IN58[2], w2082, w2083);
  FullAdder U622 (w2083, w2060, IN59[1], w2084, w2085);
  FullAdder U623 (w2085, w2061, IN60[0], w2086, w2087);
  HalfAdder U624 (w2064, IN49[12], Out1[49], w2089);
  FullAdder U625 (w2089, w2066, IN50[11], w2090, w2091);
  FullAdder U626 (w2091, w2068, IN51[10], w2092, w2093);
  FullAdder U627 (w2093, w2070, IN52[9], w2094, w2095);
  FullAdder U628 (w2095, w2072, IN53[8], w2096, w2097);
  FullAdder U629 (w2097, w2074, IN54[7], w2098, w2099);
  FullAdder U630 (w2099, w2076, IN55[6], w2100, w2101);
  FullAdder U631 (w2101, w2078, IN56[5], w2102, w2103);
  FullAdder U632 (w2103, w2080, IN57[4], w2104, w2105);
  FullAdder U633 (w2105, w2082, IN58[3], w2106, w2107);
  FullAdder U634 (w2107, w2084, IN59[2], w2108, w2109);
  FullAdder U635 (w2109, w2086, IN60[1], w2110, w2111);
  FullAdder U636 (w2111, w2087, IN61[0], w2112, w2113);
  HalfAdder U637 (w2090, IN50[12], Out1[50], w2115);
  FullAdder U638 (w2115, w2092, IN51[11], w2116, w2117);
  FullAdder U639 (w2117, w2094, IN52[10], w2118, w2119);
  FullAdder U640 (w2119, w2096, IN53[9], w2120, w2121);
  FullAdder U641 (w2121, w2098, IN54[8], w2122, w2123);
  FullAdder U642 (w2123, w2100, IN55[7], w2124, w2125);
  FullAdder U643 (w2125, w2102, IN56[6], w2126, w2127);
  FullAdder U644 (w2127, w2104, IN57[5], w2128, w2129);
  FullAdder U645 (w2129, w2106, IN58[4], w2130, w2131);
  FullAdder U646 (w2131, w2108, IN59[3], w2132, w2133);
  FullAdder U647 (w2133, w2110, IN60[2], w2134, w2135);
  FullAdder U648 (w2135, w2112, IN61[1], w2136, w2137);
  FullAdder U649 (w2137, w2113, IN62[0], w2138, w2139);
  HalfAdder U650 (w2116, IN51[12], Out1[51], w2141);
  FullAdder U651 (w2141, w2118, IN52[11], w2142, w2143);
  FullAdder U652 (w2143, w2120, IN53[10], w2144, w2145);
  FullAdder U653 (w2145, w2122, IN54[9], w2146, w2147);
  FullAdder U654 (w2147, w2124, IN55[8], w2148, w2149);
  FullAdder U655 (w2149, w2126, IN56[7], w2150, w2151);
  FullAdder U656 (w2151, w2128, IN57[6], w2152, w2153);
  FullAdder U657 (w2153, w2130, IN58[5], w2154, w2155);
  FullAdder U658 (w2155, w2132, IN59[4], w2156, w2157);
  FullAdder U659 (w2157, w2134, IN60[3], w2158, w2159);
  FullAdder U660 (w2159, w2136, IN61[2], w2160, w2161);
  FullAdder U661 (w2161, w2138, IN62[1], w2162, w2163);
  FullAdder U662 (w2163, w2139, IN63[0], w2164, w2165);
  HalfAdder U663 (w2142, IN52[12], Out1[52], w2167);
  FullAdder U664 (w2167, w2144, IN53[11], w2168, w2169);
  FullAdder U665 (w2169, w2146, IN54[10], w2170, w2171);
  FullAdder U666 (w2171, w2148, IN55[9], w2172, w2173);
  FullAdder U667 (w2173, w2150, IN56[8], w2174, w2175);
  FullAdder U668 (w2175, w2152, IN57[7], w2176, w2177);
  FullAdder U669 (w2177, w2154, IN58[6], w2178, w2179);
  FullAdder U670 (w2179, w2156, IN59[5], w2180, w2181);
  FullAdder U671 (w2181, w2158, IN60[4], w2182, w2183);
  FullAdder U672 (w2183, w2160, IN61[3], w2184, w2185);
  FullAdder U673 (w2185, w2162, IN62[2], w2186, w2187);
  FullAdder U674 (w2187, w2164, IN63[1], w2188, w2189);
  FullAdder U675 (w2189, w2165, IN64[0], w2190, w2191);
  HalfAdder U676 (w2168, IN53[12], Out1[53], w2193);
  FullAdder U677 (w2193, w2170, IN54[11], w2194, w2195);
  FullAdder U678 (w2195, w2172, IN55[10], w2196, w2197);
  FullAdder U679 (w2197, w2174, IN56[9], w2198, w2199);
  FullAdder U680 (w2199, w2176, IN57[8], w2200, w2201);
  FullAdder U681 (w2201, w2178, IN58[7], w2202, w2203);
  FullAdder U682 (w2203, w2180, IN59[6], w2204, w2205);
  FullAdder U683 (w2205, w2182, IN60[5], w2206, w2207);
  FullAdder U684 (w2207, w2184, IN61[4], w2208, w2209);
  FullAdder U685 (w2209, w2186, IN62[3], w2210, w2211);
  FullAdder U686 (w2211, w2188, IN63[2], w2212, w2213);
  FullAdder U687 (w2213, w2190, IN64[1], w2214, w2215);
  FullAdder U688 (w2215, w2191, IN65[0], w2216, w2217);
  HalfAdder U689 (w2194, IN54[12], Out1[54], w2219);
  FullAdder U690 (w2219, w2196, IN55[11], w2220, w2221);
  FullAdder U691 (w2221, w2198, IN56[10], w2222, w2223);
  FullAdder U692 (w2223, w2200, IN57[9], w2224, w2225);
  FullAdder U693 (w2225, w2202, IN58[8], w2226, w2227);
  FullAdder U694 (w2227, w2204, IN59[7], w2228, w2229);
  FullAdder U695 (w2229, w2206, IN60[6], w2230, w2231);
  FullAdder U696 (w2231, w2208, IN61[5], w2232, w2233);
  FullAdder U697 (w2233, w2210, IN62[4], w2234, w2235);
  FullAdder U698 (w2235, w2212, IN63[3], w2236, w2237);
  FullAdder U699 (w2237, w2214, IN64[2], w2238, w2239);
  FullAdder U700 (w2239, w2216, IN65[1], w2240, w2241);
  FullAdder U701 (w2241, w2217, IN66[0], w2242, w2243);
  HalfAdder U702 (w2220, IN55[12], Out1[55], w2245);
  FullAdder U703 (w2245, w2222, IN56[11], w2246, w2247);
  FullAdder U704 (w2247, w2224, IN57[10], w2248, w2249);
  FullAdder U705 (w2249, w2226, IN58[9], w2250, w2251);
  FullAdder U706 (w2251, w2228, IN59[8], w2252, w2253);
  FullAdder U707 (w2253, w2230, IN60[7], w2254, w2255);
  FullAdder U708 (w2255, w2232, IN61[6], w2256, w2257);
  FullAdder U709 (w2257, w2234, IN62[5], w2258, w2259);
  FullAdder U710 (w2259, w2236, IN63[4], w2260, w2261);
  FullAdder U711 (w2261, w2238, IN64[3], w2262, w2263);
  FullAdder U712 (w2263, w2240, IN65[2], w2264, w2265);
  FullAdder U713 (w2265, w2242, IN66[1], w2266, w2267);
  FullAdder U714 (w2267, w2243, IN67[0], w2268, w2269);
  HalfAdder U715 (w2246, IN56[12], Out1[56], w2271);
  FullAdder U716 (w2271, w2248, IN57[11], w2272, w2273);
  FullAdder U717 (w2273, w2250, IN58[10], w2274, w2275);
  FullAdder U718 (w2275, w2252, IN59[9], w2276, w2277);
  FullAdder U719 (w2277, w2254, IN60[8], w2278, w2279);
  FullAdder U720 (w2279, w2256, IN61[7], w2280, w2281);
  FullAdder U721 (w2281, w2258, IN62[6], w2282, w2283);
  FullAdder U722 (w2283, w2260, IN63[5], w2284, w2285);
  FullAdder U723 (w2285, w2262, IN64[4], w2286, w2287);
  FullAdder U724 (w2287, w2264, IN65[3], w2288, w2289);
  FullAdder U725 (w2289, w2266, IN66[2], w2290, w2291);
  FullAdder U726 (w2291, w2268, IN67[1], w2292, w2293);
  FullAdder U727 (w2293, w2269, IN68[0], w2294, w2295);
  HalfAdder U728 (w2272, IN57[12], Out1[57], w2297);
  FullAdder U729 (w2297, w2274, IN58[11], w2298, w2299);
  FullAdder U730 (w2299, w2276, IN59[10], w2300, w2301);
  FullAdder U731 (w2301, w2278, IN60[9], w2302, w2303);
  FullAdder U732 (w2303, w2280, IN61[8], w2304, w2305);
  FullAdder U733 (w2305, w2282, IN62[7], w2306, w2307);
  FullAdder U734 (w2307, w2284, IN63[6], w2308, w2309);
  FullAdder U735 (w2309, w2286, IN64[5], w2310, w2311);
  FullAdder U736 (w2311, w2288, IN65[4], w2312, w2313);
  FullAdder U737 (w2313, w2290, IN66[3], w2314, w2315);
  FullAdder U738 (w2315, w2292, IN67[2], w2316, w2317);
  FullAdder U739 (w2317, w2294, IN68[1], w2318, w2319);
  FullAdder U740 (w2319, w2295, IN69[0], w2320, w2321);
  HalfAdder U741 (w2298, IN58[12], Out1[58], w2323);
  FullAdder U742 (w2323, w2300, IN59[11], w2324, w2325);
  FullAdder U743 (w2325, w2302, IN60[10], w2326, w2327);
  FullAdder U744 (w2327, w2304, IN61[9], w2328, w2329);
  FullAdder U745 (w2329, w2306, IN62[8], w2330, w2331);
  FullAdder U746 (w2331, w2308, IN63[7], w2332, w2333);
  FullAdder U747 (w2333, w2310, IN64[6], w2334, w2335);
  FullAdder U748 (w2335, w2312, IN65[5], w2336, w2337);
  FullAdder U749 (w2337, w2314, IN66[4], w2338, w2339);
  FullAdder U750 (w2339, w2316, IN67[3], w2340, w2341);
  FullAdder U751 (w2341, w2318, IN68[2], w2342, w2343);
  FullAdder U752 (w2343, w2320, IN69[1], w2344, w2345);
  FullAdder U753 (w2345, w2321, IN70[0], w2346, w2347);
  HalfAdder U754 (w2324, IN59[12], Out1[59], w2349);
  FullAdder U755 (w2349, w2326, IN60[11], Out1[60], w2351);
  FullAdder U756 (w2351, w2328, IN61[10], Out1[61], w2353);
  FullAdder U757 (w2353, w2330, IN62[9], Out1[62], w2355);
  FullAdder U758 (w2355, w2332, IN63[8], Out1[63], w2357);
  FullAdder U759 (w2357, w2334, IN64[7], Out1[64], w2359);
  FullAdder U760 (w2359, w2336, IN65[6], Out1[65], w2361);
  FullAdder U761 (w2361, w2338, IN66[5], Out1[66], w2363);
  FullAdder U762 (w2363, w2340, IN67[4], Out1[67], w2365);
  FullAdder U763 (w2365, w2342, IN68[3], Out1[68], w2367);
  FullAdder U764 (w2367, w2344, IN69[2], Out1[69], w2369);
  FullAdder U765 (w2369, w2346, IN70[1], Out1[70], w2371);
  FullAdder U766 (w2371, w2347, IN71[0], Out1[71], Out1[72]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN14[13];
  assign Out2[1] = IN15[13];
  assign Out2[2] = IN16[13];
  assign Out2[3] = IN17[13];
  assign Out2[4] = IN18[13];
  assign Out2[5] = IN19[13];
  assign Out2[6] = IN20[13];
  assign Out2[7] = IN21[13];
  assign Out2[8] = IN22[13];
  assign Out2[9] = IN23[13];
  assign Out2[10] = IN24[13];
  assign Out2[11] = IN25[13];
  assign Out2[12] = IN26[13];
  assign Out2[13] = IN27[13];
  assign Out2[14] = IN28[13];
  assign Out2[15] = IN29[13];
  assign Out2[16] = IN30[13];
  assign Out2[17] = IN31[13];
  assign Out2[18] = IN32[13];
  assign Out2[19] = IN33[13];
  assign Out2[20] = IN34[13];
  assign Out2[21] = IN35[13];
  assign Out2[22] = IN36[13];
  assign Out2[23] = IN37[13];
  assign Out2[24] = IN38[13];
  assign Out2[25] = IN39[13];
  assign Out2[26] = IN40[13];
  assign Out2[27] = IN41[13];
  assign Out2[28] = IN42[13];
  assign Out2[29] = IN43[13];
  assign Out2[30] = IN44[13];
  assign Out2[31] = IN45[13];
  assign Out2[32] = IN46[13];
  assign Out2[33] = IN47[13];
  assign Out2[34] = IN48[13];
  assign Out2[35] = IN49[13];
  assign Out2[36] = IN50[13];
  assign Out2[37] = IN51[13];
  assign Out2[38] = IN52[13];
  assign Out2[39] = IN53[13];
  assign Out2[40] = IN54[13];
  assign Out2[41] = IN55[13];
  assign Out2[42] = IN56[13];
  assign Out2[43] = IN57[13];
  assign Out2[44] = IN58[13];
  assign Out2[45] = IN59[13];
  assign Out2[46] = IN60[12];
  assign Out2[47] = IN61[11];
  assign Out2[48] = IN62[10];
  assign Out2[49] = IN63[9];
  assign Out2[50] = IN64[8];
  assign Out2[51] = IN65[7];
  assign Out2[52] = IN66[6];
  assign Out2[53] = IN67[5];
  assign Out2[54] = IN68[4];
  assign Out2[55] = IN69[3];
  assign Out2[56] = IN70[2];
  assign Out2[57] = IN71[1];
  assign Out2[58] = IN72[0];

endmodule
module RC_59_59(IN1, IN2, Out);
  input [58:0] IN1;
  input [58:0] IN2;
  output [59:0] Out;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  wire w231;
  wire w233;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w119);
  FullAdder U1 (IN1[1], IN2[1], w119, Out[1], w121);
  FullAdder U2 (IN1[2], IN2[2], w121, Out[2], w123);
  FullAdder U3 (IN1[3], IN2[3], w123, Out[3], w125);
  FullAdder U4 (IN1[4], IN2[4], w125, Out[4], w127);
  FullAdder U5 (IN1[5], IN2[5], w127, Out[5], w129);
  FullAdder U6 (IN1[6], IN2[6], w129, Out[6], w131);
  FullAdder U7 (IN1[7], IN2[7], w131, Out[7], w133);
  FullAdder U8 (IN1[8], IN2[8], w133, Out[8], w135);
  FullAdder U9 (IN1[9], IN2[9], w135, Out[9], w137);
  FullAdder U10 (IN1[10], IN2[10], w137, Out[10], w139);
  FullAdder U11 (IN1[11], IN2[11], w139, Out[11], w141);
  FullAdder U12 (IN1[12], IN2[12], w141, Out[12], w143);
  FullAdder U13 (IN1[13], IN2[13], w143, Out[13], w145);
  FullAdder U14 (IN1[14], IN2[14], w145, Out[14], w147);
  FullAdder U15 (IN1[15], IN2[15], w147, Out[15], w149);
  FullAdder U16 (IN1[16], IN2[16], w149, Out[16], w151);
  FullAdder U17 (IN1[17], IN2[17], w151, Out[17], w153);
  FullAdder U18 (IN1[18], IN2[18], w153, Out[18], w155);
  FullAdder U19 (IN1[19], IN2[19], w155, Out[19], w157);
  FullAdder U20 (IN1[20], IN2[20], w157, Out[20], w159);
  FullAdder U21 (IN1[21], IN2[21], w159, Out[21], w161);
  FullAdder U22 (IN1[22], IN2[22], w161, Out[22], w163);
  FullAdder U23 (IN1[23], IN2[23], w163, Out[23], w165);
  FullAdder U24 (IN1[24], IN2[24], w165, Out[24], w167);
  FullAdder U25 (IN1[25], IN2[25], w167, Out[25], w169);
  FullAdder U26 (IN1[26], IN2[26], w169, Out[26], w171);
  FullAdder U27 (IN1[27], IN2[27], w171, Out[27], w173);
  FullAdder U28 (IN1[28], IN2[28], w173, Out[28], w175);
  FullAdder U29 (IN1[29], IN2[29], w175, Out[29], w177);
  FullAdder U30 (IN1[30], IN2[30], w177, Out[30], w179);
  FullAdder U31 (IN1[31], IN2[31], w179, Out[31], w181);
  FullAdder U32 (IN1[32], IN2[32], w181, Out[32], w183);
  FullAdder U33 (IN1[33], IN2[33], w183, Out[33], w185);
  FullAdder U34 (IN1[34], IN2[34], w185, Out[34], w187);
  FullAdder U35 (IN1[35], IN2[35], w187, Out[35], w189);
  FullAdder U36 (IN1[36], IN2[36], w189, Out[36], w191);
  FullAdder U37 (IN1[37], IN2[37], w191, Out[37], w193);
  FullAdder U38 (IN1[38], IN2[38], w193, Out[38], w195);
  FullAdder U39 (IN1[39], IN2[39], w195, Out[39], w197);
  FullAdder U40 (IN1[40], IN2[40], w197, Out[40], w199);
  FullAdder U41 (IN1[41], IN2[41], w199, Out[41], w201);
  FullAdder U42 (IN1[42], IN2[42], w201, Out[42], w203);
  FullAdder U43 (IN1[43], IN2[43], w203, Out[43], w205);
  FullAdder U44 (IN1[44], IN2[44], w205, Out[44], w207);
  FullAdder U45 (IN1[45], IN2[45], w207, Out[45], w209);
  FullAdder U46 (IN1[46], IN2[46], w209, Out[46], w211);
  FullAdder U47 (IN1[47], IN2[47], w211, Out[47], w213);
  FullAdder U48 (IN1[48], IN2[48], w213, Out[48], w215);
  FullAdder U49 (IN1[49], IN2[49], w215, Out[49], w217);
  FullAdder U50 (IN1[50], IN2[50], w217, Out[50], w219);
  FullAdder U51 (IN1[51], IN2[51], w219, Out[51], w221);
  FullAdder U52 (IN1[52], IN2[52], w221, Out[52], w223);
  FullAdder U53 (IN1[53], IN2[53], w223, Out[53], w225);
  FullAdder U54 (IN1[54], IN2[54], w225, Out[54], w227);
  FullAdder U55 (IN1[55], IN2[55], w227, Out[55], w229);
  FullAdder U56 (IN1[56], IN2[56], w229, Out[56], w231);
  FullAdder U57 (IN1[57], IN2[57], w231, Out[57], w233);
  FullAdder U58 (IN1[58], IN2[58], w233, Out[58], Out[59]);

endmodule
module NR_14_60(IN1, IN2, Out);
  input [13:0] IN1;
  input [59:0] IN2;
  output [73:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [13:0] P14;
  wire [13:0] P15;
  wire [13:0] P16;
  wire [13:0] P17;
  wire [13:0] P18;
  wire [13:0] P19;
  wire [13:0] P20;
  wire [13:0] P21;
  wire [13:0] P22;
  wire [13:0] P23;
  wire [13:0] P24;
  wire [13:0] P25;
  wire [13:0] P26;
  wire [13:0] P27;
  wire [13:0] P28;
  wire [13:0] P29;
  wire [13:0] P30;
  wire [13:0] P31;
  wire [13:0] P32;
  wire [13:0] P33;
  wire [13:0] P34;
  wire [13:0] P35;
  wire [13:0] P36;
  wire [13:0] P37;
  wire [13:0] P38;
  wire [13:0] P39;
  wire [13:0] P40;
  wire [13:0] P41;
  wire [13:0] P42;
  wire [13:0] P43;
  wire [13:0] P44;
  wire [13:0] P45;
  wire [13:0] P46;
  wire [13:0] P47;
  wire [13:0] P48;
  wire [13:0] P49;
  wire [13:0] P50;
  wire [13:0] P51;
  wire [13:0] P52;
  wire [13:0] P53;
  wire [13:0] P54;
  wire [13:0] P55;
  wire [13:0] P56;
  wire [13:0] P57;
  wire [13:0] P58;
  wire [13:0] P59;
  wire [12:0] P60;
  wire [11:0] P61;
  wire [10:0] P62;
  wire [9:0] P63;
  wire [8:0] P64;
  wire [7:0] P65;
  wire [6:0] P66;
  wire [5:0] P67;
  wire [4:0] P68;
  wire [3:0] P69;
  wire [2:0] P70;
  wire [1:0] P71;
  wire [0:0] P72;
  wire [72:0] R1;
  wire [58:0] R2;
  wire [73:0] aOut;
  U_SP_14_60 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, R1, R2);
  RC_59_59 S2 (R1[72:14], R2, aOut[73:14]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign Out = aOut[73:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
