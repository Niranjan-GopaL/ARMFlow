
module customAdder46_0(
    input [45 : 0] A,
    input [45 : 0] B,
    output [46 : 0] Sum
);

    assign Sum = A+B;

endmodule
