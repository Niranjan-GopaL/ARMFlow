
module customAdder37_0(
    input [36 : 0] A,
    input [36 : 0] B,
    output [37 : 0] Sum
);

    assign Sum = A+B;

endmodule
