
module customAdder55_0(
    input [54 : 0] A,
    input [54 : 0] B,
    output [55 : 0] Sum
);

    assign Sum = A+B;

endmodule
