
module NR_1_40(
    input [0:0]IN1,
    input [39:0]IN2,
    output [39:0]Out
);
    assign Out = IN2;
endmodule
