//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 8
  second input length: 45
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_8_45(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51);
  input [7:0] IN1;
  input [44:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [7:0] P8;
  output [7:0] P9;
  output [7:0] P10;
  output [7:0] P11;
  output [7:0] P12;
  output [7:0] P13;
  output [7:0] P14;
  output [7:0] P15;
  output [7:0] P16;
  output [7:0] P17;
  output [7:0] P18;
  output [7:0] P19;
  output [7:0] P20;
  output [7:0] P21;
  output [7:0] P22;
  output [7:0] P23;
  output [7:0] P24;
  output [7:0] P25;
  output [7:0] P26;
  output [7:0] P27;
  output [7:0] P28;
  output [7:0] P29;
  output [7:0] P30;
  output [7:0] P31;
  output [7:0] P32;
  output [7:0] P33;
  output [7:0] P34;
  output [7:0] P35;
  output [7:0] P36;
  output [7:0] P37;
  output [7:0] P38;
  output [7:0] P39;
  output [7:0] P40;
  output [7:0] P41;
  output [7:0] P42;
  output [7:0] P43;
  output [7:0] P44;
  output [6:0] P45;
  output [5:0] P46;
  output [4:0] P47;
  output [3:0] P48;
  output [2:0] P49;
  output [1:0] P50;
  output [0:0] P51;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[0] = IN1[1]&IN2[44];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[1] = IN1[2]&IN2[43];
  assign P46[0] = IN1[2]&IN2[44];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[2] = IN1[3]&IN2[42];
  assign P46[1] = IN1[3]&IN2[43];
  assign P47[0] = IN1[3]&IN2[44];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[3] = IN1[4]&IN2[41];
  assign P46[2] = IN1[4]&IN2[42];
  assign P47[1] = IN1[4]&IN2[43];
  assign P48[0] = IN1[4]&IN2[44];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[4] = IN1[5]&IN2[40];
  assign P46[3] = IN1[5]&IN2[41];
  assign P47[2] = IN1[5]&IN2[42];
  assign P48[1] = IN1[5]&IN2[43];
  assign P49[0] = IN1[5]&IN2[44];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[5] = IN1[6]&IN2[39];
  assign P46[4] = IN1[6]&IN2[40];
  assign P47[3] = IN1[6]&IN2[41];
  assign P48[2] = IN1[6]&IN2[42];
  assign P49[1] = IN1[6]&IN2[43];
  assign P50[0] = IN1[6]&IN2[44];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[6] = IN1[7]&IN2[38];
  assign P46[5] = IN1[7]&IN2[39];
  assign P47[4] = IN1[7]&IN2[40];
  assign P48[3] = IN1[7]&IN2[41];
  assign P49[2] = IN1[7]&IN2[42];
  assign P50[1] = IN1[7]&IN2[43];
  assign P51[0] = IN1[7]&IN2[44];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [7:0] IN8;
  input [7:0] IN9;
  input [7:0] IN10;
  input [7:0] IN11;
  input [7:0] IN12;
  input [7:0] IN13;
  input [7:0] IN14;
  input [7:0] IN15;
  input [7:0] IN16;
  input [7:0] IN17;
  input [7:0] IN18;
  input [7:0] IN19;
  input [7:0] IN20;
  input [7:0] IN21;
  input [7:0] IN22;
  input [7:0] IN23;
  input [7:0] IN24;
  input [7:0] IN25;
  input [7:0] IN26;
  input [7:0] IN27;
  input [7:0] IN28;
  input [7:0] IN29;
  input [7:0] IN30;
  input [7:0] IN31;
  input [7:0] IN32;
  input [7:0] IN33;
  input [7:0] IN34;
  input [7:0] IN35;
  input [7:0] IN36;
  input [7:0] IN37;
  input [7:0] IN38;
  input [7:0] IN39;
  input [7:0] IN40;
  input [7:0] IN41;
  input [7:0] IN42;
  input [7:0] IN43;
  input [7:0] IN44;
  input [6:0] IN45;
  input [5:0] IN46;
  input [4:0] IN47;
  input [3:0] IN48;
  input [2:0] IN49;
  input [1:0] IN50;
  input [0:0] IN51;
  output [51:0] Out1;
  output [43:0] Out2;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w963;
  wire w965;
  wire w967;
  wire w969;
  wire w971;
  wire w973;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w361);
  FullAdder U1 (w361, IN2[0], IN2[1], w362, w363);
  FullAdder U2 (w363, IN3[0], IN3[1], w364, w365);
  FullAdder U3 (w365, IN4[0], IN4[1], w366, w367);
  FullAdder U4 (w367, IN5[0], IN5[1], w368, w369);
  FullAdder U5 (w369, IN6[0], IN6[1], w370, w371);
  FullAdder U6 (w371, IN7[0], IN7[1], w372, w373);
  HalfAdder U7 (w362, IN2[2], Out1[2], w375);
  FullAdder U8 (w375, w364, IN3[2], w376, w377);
  FullAdder U9 (w377, w366, IN4[2], w378, w379);
  FullAdder U10 (w379, w368, IN5[2], w380, w381);
  FullAdder U11 (w381, w370, IN6[2], w382, w383);
  FullAdder U12 (w383, w372, IN7[2], w384, w385);
  FullAdder U13 (w385, w373, IN8[0], w386, w387);
  HalfAdder U14 (w376, IN3[3], Out1[3], w389);
  FullAdder U15 (w389, w378, IN4[3], w390, w391);
  FullAdder U16 (w391, w380, IN5[3], w392, w393);
  FullAdder U17 (w393, w382, IN6[3], w394, w395);
  FullAdder U18 (w395, w384, IN7[3], w396, w397);
  FullAdder U19 (w397, w386, IN8[1], w398, w399);
  FullAdder U20 (w399, w387, IN9[0], w400, w401);
  HalfAdder U21 (w390, IN4[4], Out1[4], w403);
  FullAdder U22 (w403, w392, IN5[4], w404, w405);
  FullAdder U23 (w405, w394, IN6[4], w406, w407);
  FullAdder U24 (w407, w396, IN7[4], w408, w409);
  FullAdder U25 (w409, w398, IN8[2], w410, w411);
  FullAdder U26 (w411, w400, IN9[1], w412, w413);
  FullAdder U27 (w413, w401, IN10[0], w414, w415);
  HalfAdder U28 (w404, IN5[5], Out1[5], w417);
  FullAdder U29 (w417, w406, IN6[5], w418, w419);
  FullAdder U30 (w419, w408, IN7[5], w420, w421);
  FullAdder U31 (w421, w410, IN8[3], w422, w423);
  FullAdder U32 (w423, w412, IN9[2], w424, w425);
  FullAdder U33 (w425, w414, IN10[1], w426, w427);
  FullAdder U34 (w427, w415, IN11[0], w428, w429);
  HalfAdder U35 (w418, IN6[6], Out1[6], w431);
  FullAdder U36 (w431, w420, IN7[6], w432, w433);
  FullAdder U37 (w433, w422, IN8[4], w434, w435);
  FullAdder U38 (w435, w424, IN9[3], w436, w437);
  FullAdder U39 (w437, w426, IN10[2], w438, w439);
  FullAdder U40 (w439, w428, IN11[1], w440, w441);
  FullAdder U41 (w441, w429, IN12[0], w442, w443);
  HalfAdder U42 (w432, IN7[7], Out1[7], w445);
  FullAdder U43 (w445, w434, IN8[5], w446, w447);
  FullAdder U44 (w447, w436, IN9[4], w448, w449);
  FullAdder U45 (w449, w438, IN10[3], w450, w451);
  FullAdder U46 (w451, w440, IN11[2], w452, w453);
  FullAdder U47 (w453, w442, IN12[1], w454, w455);
  FullAdder U48 (w455, w443, IN13[0], w456, w457);
  HalfAdder U49 (w446, IN8[6], Out1[8], w459);
  FullAdder U50 (w459, w448, IN9[5], w460, w461);
  FullAdder U51 (w461, w450, IN10[4], w462, w463);
  FullAdder U52 (w463, w452, IN11[3], w464, w465);
  FullAdder U53 (w465, w454, IN12[2], w466, w467);
  FullAdder U54 (w467, w456, IN13[1], w468, w469);
  FullAdder U55 (w469, w457, IN14[0], w470, w471);
  HalfAdder U56 (w460, IN9[6], Out1[9], w473);
  FullAdder U57 (w473, w462, IN10[5], w474, w475);
  FullAdder U58 (w475, w464, IN11[4], w476, w477);
  FullAdder U59 (w477, w466, IN12[3], w478, w479);
  FullAdder U60 (w479, w468, IN13[2], w480, w481);
  FullAdder U61 (w481, w470, IN14[1], w482, w483);
  FullAdder U62 (w483, w471, IN15[0], w484, w485);
  HalfAdder U63 (w474, IN10[6], Out1[10], w487);
  FullAdder U64 (w487, w476, IN11[5], w488, w489);
  FullAdder U65 (w489, w478, IN12[4], w490, w491);
  FullAdder U66 (w491, w480, IN13[3], w492, w493);
  FullAdder U67 (w493, w482, IN14[2], w494, w495);
  FullAdder U68 (w495, w484, IN15[1], w496, w497);
  FullAdder U69 (w497, w485, IN16[0], w498, w499);
  HalfAdder U70 (w488, IN11[6], Out1[11], w501);
  FullAdder U71 (w501, w490, IN12[5], w502, w503);
  FullAdder U72 (w503, w492, IN13[4], w504, w505);
  FullAdder U73 (w505, w494, IN14[3], w506, w507);
  FullAdder U74 (w507, w496, IN15[2], w508, w509);
  FullAdder U75 (w509, w498, IN16[1], w510, w511);
  FullAdder U76 (w511, w499, IN17[0], w512, w513);
  HalfAdder U77 (w502, IN12[6], Out1[12], w515);
  FullAdder U78 (w515, w504, IN13[5], w516, w517);
  FullAdder U79 (w517, w506, IN14[4], w518, w519);
  FullAdder U80 (w519, w508, IN15[3], w520, w521);
  FullAdder U81 (w521, w510, IN16[2], w522, w523);
  FullAdder U82 (w523, w512, IN17[1], w524, w525);
  FullAdder U83 (w525, w513, IN18[0], w526, w527);
  HalfAdder U84 (w516, IN13[6], Out1[13], w529);
  FullAdder U85 (w529, w518, IN14[5], w530, w531);
  FullAdder U86 (w531, w520, IN15[4], w532, w533);
  FullAdder U87 (w533, w522, IN16[3], w534, w535);
  FullAdder U88 (w535, w524, IN17[2], w536, w537);
  FullAdder U89 (w537, w526, IN18[1], w538, w539);
  FullAdder U90 (w539, w527, IN19[0], w540, w541);
  HalfAdder U91 (w530, IN14[6], Out1[14], w543);
  FullAdder U92 (w543, w532, IN15[5], w544, w545);
  FullAdder U93 (w545, w534, IN16[4], w546, w547);
  FullAdder U94 (w547, w536, IN17[3], w548, w549);
  FullAdder U95 (w549, w538, IN18[2], w550, w551);
  FullAdder U96 (w551, w540, IN19[1], w552, w553);
  FullAdder U97 (w553, w541, IN20[0], w554, w555);
  HalfAdder U98 (w544, IN15[6], Out1[15], w557);
  FullAdder U99 (w557, w546, IN16[5], w558, w559);
  FullAdder U100 (w559, w548, IN17[4], w560, w561);
  FullAdder U101 (w561, w550, IN18[3], w562, w563);
  FullAdder U102 (w563, w552, IN19[2], w564, w565);
  FullAdder U103 (w565, w554, IN20[1], w566, w567);
  FullAdder U104 (w567, w555, IN21[0], w568, w569);
  HalfAdder U105 (w558, IN16[6], Out1[16], w571);
  FullAdder U106 (w571, w560, IN17[5], w572, w573);
  FullAdder U107 (w573, w562, IN18[4], w574, w575);
  FullAdder U108 (w575, w564, IN19[3], w576, w577);
  FullAdder U109 (w577, w566, IN20[2], w578, w579);
  FullAdder U110 (w579, w568, IN21[1], w580, w581);
  FullAdder U111 (w581, w569, IN22[0], w582, w583);
  HalfAdder U112 (w572, IN17[6], Out1[17], w585);
  FullAdder U113 (w585, w574, IN18[5], w586, w587);
  FullAdder U114 (w587, w576, IN19[4], w588, w589);
  FullAdder U115 (w589, w578, IN20[3], w590, w591);
  FullAdder U116 (w591, w580, IN21[2], w592, w593);
  FullAdder U117 (w593, w582, IN22[1], w594, w595);
  FullAdder U118 (w595, w583, IN23[0], w596, w597);
  HalfAdder U119 (w586, IN18[6], Out1[18], w599);
  FullAdder U120 (w599, w588, IN19[5], w600, w601);
  FullAdder U121 (w601, w590, IN20[4], w602, w603);
  FullAdder U122 (w603, w592, IN21[3], w604, w605);
  FullAdder U123 (w605, w594, IN22[2], w606, w607);
  FullAdder U124 (w607, w596, IN23[1], w608, w609);
  FullAdder U125 (w609, w597, IN24[0], w610, w611);
  HalfAdder U126 (w600, IN19[6], Out1[19], w613);
  FullAdder U127 (w613, w602, IN20[5], w614, w615);
  FullAdder U128 (w615, w604, IN21[4], w616, w617);
  FullAdder U129 (w617, w606, IN22[3], w618, w619);
  FullAdder U130 (w619, w608, IN23[2], w620, w621);
  FullAdder U131 (w621, w610, IN24[1], w622, w623);
  FullAdder U132 (w623, w611, IN25[0], w624, w625);
  HalfAdder U133 (w614, IN20[6], Out1[20], w627);
  FullAdder U134 (w627, w616, IN21[5], w628, w629);
  FullAdder U135 (w629, w618, IN22[4], w630, w631);
  FullAdder U136 (w631, w620, IN23[3], w632, w633);
  FullAdder U137 (w633, w622, IN24[2], w634, w635);
  FullAdder U138 (w635, w624, IN25[1], w636, w637);
  FullAdder U139 (w637, w625, IN26[0], w638, w639);
  HalfAdder U140 (w628, IN21[6], Out1[21], w641);
  FullAdder U141 (w641, w630, IN22[5], w642, w643);
  FullAdder U142 (w643, w632, IN23[4], w644, w645);
  FullAdder U143 (w645, w634, IN24[3], w646, w647);
  FullAdder U144 (w647, w636, IN25[2], w648, w649);
  FullAdder U145 (w649, w638, IN26[1], w650, w651);
  FullAdder U146 (w651, w639, IN27[0], w652, w653);
  HalfAdder U147 (w642, IN22[6], Out1[22], w655);
  FullAdder U148 (w655, w644, IN23[5], w656, w657);
  FullAdder U149 (w657, w646, IN24[4], w658, w659);
  FullAdder U150 (w659, w648, IN25[3], w660, w661);
  FullAdder U151 (w661, w650, IN26[2], w662, w663);
  FullAdder U152 (w663, w652, IN27[1], w664, w665);
  FullAdder U153 (w665, w653, IN28[0], w666, w667);
  HalfAdder U154 (w656, IN23[6], Out1[23], w669);
  FullAdder U155 (w669, w658, IN24[5], w670, w671);
  FullAdder U156 (w671, w660, IN25[4], w672, w673);
  FullAdder U157 (w673, w662, IN26[3], w674, w675);
  FullAdder U158 (w675, w664, IN27[2], w676, w677);
  FullAdder U159 (w677, w666, IN28[1], w678, w679);
  FullAdder U160 (w679, w667, IN29[0], w680, w681);
  HalfAdder U161 (w670, IN24[6], Out1[24], w683);
  FullAdder U162 (w683, w672, IN25[5], w684, w685);
  FullAdder U163 (w685, w674, IN26[4], w686, w687);
  FullAdder U164 (w687, w676, IN27[3], w688, w689);
  FullAdder U165 (w689, w678, IN28[2], w690, w691);
  FullAdder U166 (w691, w680, IN29[1], w692, w693);
  FullAdder U167 (w693, w681, IN30[0], w694, w695);
  HalfAdder U168 (w684, IN25[6], Out1[25], w697);
  FullAdder U169 (w697, w686, IN26[5], w698, w699);
  FullAdder U170 (w699, w688, IN27[4], w700, w701);
  FullAdder U171 (w701, w690, IN28[3], w702, w703);
  FullAdder U172 (w703, w692, IN29[2], w704, w705);
  FullAdder U173 (w705, w694, IN30[1], w706, w707);
  FullAdder U174 (w707, w695, IN31[0], w708, w709);
  HalfAdder U175 (w698, IN26[6], Out1[26], w711);
  FullAdder U176 (w711, w700, IN27[5], w712, w713);
  FullAdder U177 (w713, w702, IN28[4], w714, w715);
  FullAdder U178 (w715, w704, IN29[3], w716, w717);
  FullAdder U179 (w717, w706, IN30[2], w718, w719);
  FullAdder U180 (w719, w708, IN31[1], w720, w721);
  FullAdder U181 (w721, w709, IN32[0], w722, w723);
  HalfAdder U182 (w712, IN27[6], Out1[27], w725);
  FullAdder U183 (w725, w714, IN28[5], w726, w727);
  FullAdder U184 (w727, w716, IN29[4], w728, w729);
  FullAdder U185 (w729, w718, IN30[3], w730, w731);
  FullAdder U186 (w731, w720, IN31[2], w732, w733);
  FullAdder U187 (w733, w722, IN32[1], w734, w735);
  FullAdder U188 (w735, w723, IN33[0], w736, w737);
  HalfAdder U189 (w726, IN28[6], Out1[28], w739);
  FullAdder U190 (w739, w728, IN29[5], w740, w741);
  FullAdder U191 (w741, w730, IN30[4], w742, w743);
  FullAdder U192 (w743, w732, IN31[3], w744, w745);
  FullAdder U193 (w745, w734, IN32[2], w746, w747);
  FullAdder U194 (w747, w736, IN33[1], w748, w749);
  FullAdder U195 (w749, w737, IN34[0], w750, w751);
  HalfAdder U196 (w740, IN29[6], Out1[29], w753);
  FullAdder U197 (w753, w742, IN30[5], w754, w755);
  FullAdder U198 (w755, w744, IN31[4], w756, w757);
  FullAdder U199 (w757, w746, IN32[3], w758, w759);
  FullAdder U200 (w759, w748, IN33[2], w760, w761);
  FullAdder U201 (w761, w750, IN34[1], w762, w763);
  FullAdder U202 (w763, w751, IN35[0], w764, w765);
  HalfAdder U203 (w754, IN30[6], Out1[30], w767);
  FullAdder U204 (w767, w756, IN31[5], w768, w769);
  FullAdder U205 (w769, w758, IN32[4], w770, w771);
  FullAdder U206 (w771, w760, IN33[3], w772, w773);
  FullAdder U207 (w773, w762, IN34[2], w774, w775);
  FullAdder U208 (w775, w764, IN35[1], w776, w777);
  FullAdder U209 (w777, w765, IN36[0], w778, w779);
  HalfAdder U210 (w768, IN31[6], Out1[31], w781);
  FullAdder U211 (w781, w770, IN32[5], w782, w783);
  FullAdder U212 (w783, w772, IN33[4], w784, w785);
  FullAdder U213 (w785, w774, IN34[3], w786, w787);
  FullAdder U214 (w787, w776, IN35[2], w788, w789);
  FullAdder U215 (w789, w778, IN36[1], w790, w791);
  FullAdder U216 (w791, w779, IN37[0], w792, w793);
  HalfAdder U217 (w782, IN32[6], Out1[32], w795);
  FullAdder U218 (w795, w784, IN33[5], w796, w797);
  FullAdder U219 (w797, w786, IN34[4], w798, w799);
  FullAdder U220 (w799, w788, IN35[3], w800, w801);
  FullAdder U221 (w801, w790, IN36[2], w802, w803);
  FullAdder U222 (w803, w792, IN37[1], w804, w805);
  FullAdder U223 (w805, w793, IN38[0], w806, w807);
  HalfAdder U224 (w796, IN33[6], Out1[33], w809);
  FullAdder U225 (w809, w798, IN34[5], w810, w811);
  FullAdder U226 (w811, w800, IN35[4], w812, w813);
  FullAdder U227 (w813, w802, IN36[3], w814, w815);
  FullAdder U228 (w815, w804, IN37[2], w816, w817);
  FullAdder U229 (w817, w806, IN38[1], w818, w819);
  FullAdder U230 (w819, w807, IN39[0], w820, w821);
  HalfAdder U231 (w810, IN34[6], Out1[34], w823);
  FullAdder U232 (w823, w812, IN35[5], w824, w825);
  FullAdder U233 (w825, w814, IN36[4], w826, w827);
  FullAdder U234 (w827, w816, IN37[3], w828, w829);
  FullAdder U235 (w829, w818, IN38[2], w830, w831);
  FullAdder U236 (w831, w820, IN39[1], w832, w833);
  FullAdder U237 (w833, w821, IN40[0], w834, w835);
  HalfAdder U238 (w824, IN35[6], Out1[35], w837);
  FullAdder U239 (w837, w826, IN36[5], w838, w839);
  FullAdder U240 (w839, w828, IN37[4], w840, w841);
  FullAdder U241 (w841, w830, IN38[3], w842, w843);
  FullAdder U242 (w843, w832, IN39[2], w844, w845);
  FullAdder U243 (w845, w834, IN40[1], w846, w847);
  FullAdder U244 (w847, w835, IN41[0], w848, w849);
  HalfAdder U245 (w838, IN36[6], Out1[36], w851);
  FullAdder U246 (w851, w840, IN37[5], w852, w853);
  FullAdder U247 (w853, w842, IN38[4], w854, w855);
  FullAdder U248 (w855, w844, IN39[3], w856, w857);
  FullAdder U249 (w857, w846, IN40[2], w858, w859);
  FullAdder U250 (w859, w848, IN41[1], w860, w861);
  FullAdder U251 (w861, w849, IN42[0], w862, w863);
  HalfAdder U252 (w852, IN37[6], Out1[37], w865);
  FullAdder U253 (w865, w854, IN38[5], w866, w867);
  FullAdder U254 (w867, w856, IN39[4], w868, w869);
  FullAdder U255 (w869, w858, IN40[3], w870, w871);
  FullAdder U256 (w871, w860, IN41[2], w872, w873);
  FullAdder U257 (w873, w862, IN42[1], w874, w875);
  FullAdder U258 (w875, w863, IN43[0], w876, w877);
  HalfAdder U259 (w866, IN38[6], Out1[38], w879);
  FullAdder U260 (w879, w868, IN39[5], w880, w881);
  FullAdder U261 (w881, w870, IN40[4], w882, w883);
  FullAdder U262 (w883, w872, IN41[3], w884, w885);
  FullAdder U263 (w885, w874, IN42[2], w886, w887);
  FullAdder U264 (w887, w876, IN43[1], w888, w889);
  FullAdder U265 (w889, w877, IN44[0], w890, w891);
  HalfAdder U266 (w880, IN39[6], Out1[39], w893);
  FullAdder U267 (w893, w882, IN40[5], w894, w895);
  FullAdder U268 (w895, w884, IN41[4], w896, w897);
  FullAdder U269 (w897, w886, IN42[3], w898, w899);
  FullAdder U270 (w899, w888, IN43[2], w900, w901);
  FullAdder U271 (w901, w890, IN44[1], w902, w903);
  FullAdder U272 (w903, w891, IN45[0], w904, w905);
  HalfAdder U273 (w894, IN40[6], Out1[40], w907);
  FullAdder U274 (w907, w896, IN41[5], w908, w909);
  FullAdder U275 (w909, w898, IN42[4], w910, w911);
  FullAdder U276 (w911, w900, IN43[3], w912, w913);
  FullAdder U277 (w913, w902, IN44[2], w914, w915);
  FullAdder U278 (w915, w904, IN45[1], w916, w917);
  FullAdder U279 (w917, w905, IN46[0], w918, w919);
  HalfAdder U280 (w908, IN41[6], Out1[41], w921);
  FullAdder U281 (w921, w910, IN42[5], w922, w923);
  FullAdder U282 (w923, w912, IN43[4], w924, w925);
  FullAdder U283 (w925, w914, IN44[3], w926, w927);
  FullAdder U284 (w927, w916, IN45[2], w928, w929);
  FullAdder U285 (w929, w918, IN46[1], w930, w931);
  FullAdder U286 (w931, w919, IN47[0], w932, w933);
  HalfAdder U287 (w922, IN42[6], Out1[42], w935);
  FullAdder U288 (w935, w924, IN43[5], w936, w937);
  FullAdder U289 (w937, w926, IN44[4], w938, w939);
  FullAdder U290 (w939, w928, IN45[3], w940, w941);
  FullAdder U291 (w941, w930, IN46[2], w942, w943);
  FullAdder U292 (w943, w932, IN47[1], w944, w945);
  FullAdder U293 (w945, w933, IN48[0], w946, w947);
  HalfAdder U294 (w936, IN43[6], Out1[43], w949);
  FullAdder U295 (w949, w938, IN44[5], w950, w951);
  FullAdder U296 (w951, w940, IN45[4], w952, w953);
  FullAdder U297 (w953, w942, IN46[3], w954, w955);
  FullAdder U298 (w955, w944, IN47[2], w956, w957);
  FullAdder U299 (w957, w946, IN48[1], w958, w959);
  FullAdder U300 (w959, w947, IN49[0], w960, w961);
  HalfAdder U301 (w950, IN44[6], Out1[44], w963);
  FullAdder U302 (w963, w952, IN45[5], Out1[45], w965);
  FullAdder U303 (w965, w954, IN46[4], Out1[46], w967);
  FullAdder U304 (w967, w956, IN47[3], Out1[47], w969);
  FullAdder U305 (w969, w958, IN48[2], Out1[48], w971);
  FullAdder U306 (w971, w960, IN49[1], Out1[49], w973);
  FullAdder U307 (w973, w961, IN50[0], Out1[50], Out1[51]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN8[7];
  assign Out2[1] = IN9[7];
  assign Out2[2] = IN10[7];
  assign Out2[3] = IN11[7];
  assign Out2[4] = IN12[7];
  assign Out2[5] = IN13[7];
  assign Out2[6] = IN14[7];
  assign Out2[7] = IN15[7];
  assign Out2[8] = IN16[7];
  assign Out2[9] = IN17[7];
  assign Out2[10] = IN18[7];
  assign Out2[11] = IN19[7];
  assign Out2[12] = IN20[7];
  assign Out2[13] = IN21[7];
  assign Out2[14] = IN22[7];
  assign Out2[15] = IN23[7];
  assign Out2[16] = IN24[7];
  assign Out2[17] = IN25[7];
  assign Out2[18] = IN26[7];
  assign Out2[19] = IN27[7];
  assign Out2[20] = IN28[7];
  assign Out2[21] = IN29[7];
  assign Out2[22] = IN30[7];
  assign Out2[23] = IN31[7];
  assign Out2[24] = IN32[7];
  assign Out2[25] = IN33[7];
  assign Out2[26] = IN34[7];
  assign Out2[27] = IN35[7];
  assign Out2[28] = IN36[7];
  assign Out2[29] = IN37[7];
  assign Out2[30] = IN38[7];
  assign Out2[31] = IN39[7];
  assign Out2[32] = IN40[7];
  assign Out2[33] = IN41[7];
  assign Out2[34] = IN42[7];
  assign Out2[35] = IN43[7];
  assign Out2[36] = IN44[7];
  assign Out2[37] = IN45[6];
  assign Out2[38] = IN46[5];
  assign Out2[39] = IN47[4];
  assign Out2[40] = IN48[3];
  assign Out2[41] = IN49[2];
  assign Out2[42] = IN50[1];
  assign Out2[43] = IN51[0];

endmodule
module RC_44_44(IN1, IN2, Out);
  input [43:0] IN1;
  input [43:0] IN2;
  output [44:0] Out;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w89);
  FullAdder U1 (IN1[1], IN2[1], w89, Out[1], w91);
  FullAdder U2 (IN1[2], IN2[2], w91, Out[2], w93);
  FullAdder U3 (IN1[3], IN2[3], w93, Out[3], w95);
  FullAdder U4 (IN1[4], IN2[4], w95, Out[4], w97);
  FullAdder U5 (IN1[5], IN2[5], w97, Out[5], w99);
  FullAdder U6 (IN1[6], IN2[6], w99, Out[6], w101);
  FullAdder U7 (IN1[7], IN2[7], w101, Out[7], w103);
  FullAdder U8 (IN1[8], IN2[8], w103, Out[8], w105);
  FullAdder U9 (IN1[9], IN2[9], w105, Out[9], w107);
  FullAdder U10 (IN1[10], IN2[10], w107, Out[10], w109);
  FullAdder U11 (IN1[11], IN2[11], w109, Out[11], w111);
  FullAdder U12 (IN1[12], IN2[12], w111, Out[12], w113);
  FullAdder U13 (IN1[13], IN2[13], w113, Out[13], w115);
  FullAdder U14 (IN1[14], IN2[14], w115, Out[14], w117);
  FullAdder U15 (IN1[15], IN2[15], w117, Out[15], w119);
  FullAdder U16 (IN1[16], IN2[16], w119, Out[16], w121);
  FullAdder U17 (IN1[17], IN2[17], w121, Out[17], w123);
  FullAdder U18 (IN1[18], IN2[18], w123, Out[18], w125);
  FullAdder U19 (IN1[19], IN2[19], w125, Out[19], w127);
  FullAdder U20 (IN1[20], IN2[20], w127, Out[20], w129);
  FullAdder U21 (IN1[21], IN2[21], w129, Out[21], w131);
  FullAdder U22 (IN1[22], IN2[22], w131, Out[22], w133);
  FullAdder U23 (IN1[23], IN2[23], w133, Out[23], w135);
  FullAdder U24 (IN1[24], IN2[24], w135, Out[24], w137);
  FullAdder U25 (IN1[25], IN2[25], w137, Out[25], w139);
  FullAdder U26 (IN1[26], IN2[26], w139, Out[26], w141);
  FullAdder U27 (IN1[27], IN2[27], w141, Out[27], w143);
  FullAdder U28 (IN1[28], IN2[28], w143, Out[28], w145);
  FullAdder U29 (IN1[29], IN2[29], w145, Out[29], w147);
  FullAdder U30 (IN1[30], IN2[30], w147, Out[30], w149);
  FullAdder U31 (IN1[31], IN2[31], w149, Out[31], w151);
  FullAdder U32 (IN1[32], IN2[32], w151, Out[32], w153);
  FullAdder U33 (IN1[33], IN2[33], w153, Out[33], w155);
  FullAdder U34 (IN1[34], IN2[34], w155, Out[34], w157);
  FullAdder U35 (IN1[35], IN2[35], w157, Out[35], w159);
  FullAdder U36 (IN1[36], IN2[36], w159, Out[36], w161);
  FullAdder U37 (IN1[37], IN2[37], w161, Out[37], w163);
  FullAdder U38 (IN1[38], IN2[38], w163, Out[38], w165);
  FullAdder U39 (IN1[39], IN2[39], w165, Out[39], w167);
  FullAdder U40 (IN1[40], IN2[40], w167, Out[40], w169);
  FullAdder U41 (IN1[41], IN2[41], w169, Out[41], w171);
  FullAdder U42 (IN1[42], IN2[42], w171, Out[42], w173);
  FullAdder U43 (IN1[43], IN2[43], w173, Out[43], Out[44]);

endmodule
module NR_8_45(IN1, IN2, Out);
  input [7:0] IN1;
  input [44:0] IN2;
  output [52:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [7:0] P8;
  wire [7:0] P9;
  wire [7:0] P10;
  wire [7:0] P11;
  wire [7:0] P12;
  wire [7:0] P13;
  wire [7:0] P14;
  wire [7:0] P15;
  wire [7:0] P16;
  wire [7:0] P17;
  wire [7:0] P18;
  wire [7:0] P19;
  wire [7:0] P20;
  wire [7:0] P21;
  wire [7:0] P22;
  wire [7:0] P23;
  wire [7:0] P24;
  wire [7:0] P25;
  wire [7:0] P26;
  wire [7:0] P27;
  wire [7:0] P28;
  wire [7:0] P29;
  wire [7:0] P30;
  wire [7:0] P31;
  wire [7:0] P32;
  wire [7:0] P33;
  wire [7:0] P34;
  wire [7:0] P35;
  wire [7:0] P36;
  wire [7:0] P37;
  wire [7:0] P38;
  wire [7:0] P39;
  wire [7:0] P40;
  wire [7:0] P41;
  wire [7:0] P42;
  wire [7:0] P43;
  wire [7:0] P44;
  wire [6:0] P45;
  wire [5:0] P46;
  wire [4:0] P47;
  wire [3:0] P48;
  wire [2:0] P49;
  wire [1:0] P50;
  wire [0:0] P51;
  wire [51:0] R1;
  wire [43:0] R2;
  wire [52:0] aOut;
  U_SP_8_45 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, R1, R2);
  RC_44_44 S2 (R1[51:8], R2, aOut[52:8]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign Out = aOut[52:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
