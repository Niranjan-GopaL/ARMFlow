
module customAdder38_0(
    input [37 : 0] A,
    input [37 : 0] B,
    output [38 : 0] Sum
);

    assign Sum = A+B;

endmodule
