
module customAdder36_0(
    input [35 : 0] A,
    input [35 : 0] B,
    output [36 : 0] Sum
);

    assign Sum = A+B;

endmodule
