
module NR_1_47(
    input [0:0]IN1,
    input [46:0]IN2,
    output [46:0]Out
);
    assign Out = IN2;
endmodule
