//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 7
  second input length: 61
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_7_61(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66);
  input [6:0] IN1;
  input [60:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [6:0] P37;
  output [6:0] P38;
  output [6:0] P39;
  output [6:0] P40;
  output [6:0] P41;
  output [6:0] P42;
  output [6:0] P43;
  output [6:0] P44;
  output [6:0] P45;
  output [6:0] P46;
  output [6:0] P47;
  output [6:0] P48;
  output [6:0] P49;
  output [6:0] P50;
  output [6:0] P51;
  output [6:0] P52;
  output [6:0] P53;
  output [6:0] P54;
  output [6:0] P55;
  output [6:0] P56;
  output [6:0] P57;
  output [6:0] P58;
  output [6:0] P59;
  output [6:0] P60;
  output [5:0] P61;
  output [4:0] P62;
  output [3:0] P63;
  output [2:0] P64;
  output [1:0] P65;
  output [0:0] P66;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P59[0] = IN1[0]&IN2[59];
  assign P60[0] = IN1[0]&IN2[60];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[1] = IN1[1]&IN2[58];
  assign P60[1] = IN1[1]&IN2[59];
  assign P61[0] = IN1[1]&IN2[60];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[2] = IN1[2]&IN2[57];
  assign P60[2] = IN1[2]&IN2[58];
  assign P61[1] = IN1[2]&IN2[59];
  assign P62[0] = IN1[2]&IN2[60];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[3] = IN1[3]&IN2[56];
  assign P60[3] = IN1[3]&IN2[57];
  assign P61[2] = IN1[3]&IN2[58];
  assign P62[1] = IN1[3]&IN2[59];
  assign P63[0] = IN1[3]&IN2[60];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[4] = IN1[4]&IN2[55];
  assign P60[4] = IN1[4]&IN2[56];
  assign P61[3] = IN1[4]&IN2[57];
  assign P62[2] = IN1[4]&IN2[58];
  assign P63[1] = IN1[4]&IN2[59];
  assign P64[0] = IN1[4]&IN2[60];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[5] = IN1[5]&IN2[54];
  assign P60[5] = IN1[5]&IN2[55];
  assign P61[4] = IN1[5]&IN2[56];
  assign P62[3] = IN1[5]&IN2[57];
  assign P63[2] = IN1[5]&IN2[58];
  assign P64[1] = IN1[5]&IN2[59];
  assign P65[0] = IN1[5]&IN2[60];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[6] = IN1[6]&IN2[53];
  assign P60[6] = IN1[6]&IN2[54];
  assign P61[5] = IN1[6]&IN2[55];
  assign P62[4] = IN1[6]&IN2[56];
  assign P63[3] = IN1[6]&IN2[57];
  assign P64[2] = IN1[6]&IN2[58];
  assign P65[1] = IN1[6]&IN2[59];
  assign P66[0] = IN1[6]&IN2[60];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [6:0] IN37;
  input [6:0] IN38;
  input [6:0] IN39;
  input [6:0] IN40;
  input [6:0] IN41;
  input [6:0] IN42;
  input [6:0] IN43;
  input [6:0] IN44;
  input [6:0] IN45;
  input [6:0] IN46;
  input [6:0] IN47;
  input [6:0] IN48;
  input [6:0] IN49;
  input [6:0] IN50;
  input [6:0] IN51;
  input [6:0] IN52;
  input [6:0] IN53;
  input [6:0] IN54;
  input [6:0] IN55;
  input [6:0] IN56;
  input [6:0] IN57;
  input [6:0] IN58;
  input [6:0] IN59;
  input [6:0] IN60;
  input [5:0] IN61;
  input [4:0] IN62;
  input [3:0] IN63;
  input [2:0] IN64;
  input [1:0] IN65;
  input [0:0] IN66;
  output [66:0] Out1;
  output [59:0] Out2;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1136;
  wire w1138;
  wire w1140;
  wire w1142;
  wire w1144;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w428);
  FullAdder U1 (w428, IN2[0], IN2[1], w429, w430);
  FullAdder U2 (w430, IN3[0], IN3[1], w431, w432);
  FullAdder U3 (w432, IN4[0], IN4[1], w433, w434);
  FullAdder U4 (w434, IN5[0], IN5[1], w435, w436);
  FullAdder U5 (w436, IN6[0], IN6[1], w437, w438);
  HalfAdder U6 (w429, IN2[2], Out1[2], w440);
  FullAdder U7 (w440, w431, IN3[2], w441, w442);
  FullAdder U8 (w442, w433, IN4[2], w443, w444);
  FullAdder U9 (w444, w435, IN5[2], w445, w446);
  FullAdder U10 (w446, w437, IN6[2], w447, w448);
  FullAdder U11 (w448, w438, IN7[0], w449, w450);
  HalfAdder U12 (w441, IN3[3], Out1[3], w452);
  FullAdder U13 (w452, w443, IN4[3], w453, w454);
  FullAdder U14 (w454, w445, IN5[3], w455, w456);
  FullAdder U15 (w456, w447, IN6[3], w457, w458);
  FullAdder U16 (w458, w449, IN7[1], w459, w460);
  FullAdder U17 (w460, w450, IN8[0], w461, w462);
  HalfAdder U18 (w453, IN4[4], Out1[4], w464);
  FullAdder U19 (w464, w455, IN5[4], w465, w466);
  FullAdder U20 (w466, w457, IN6[4], w467, w468);
  FullAdder U21 (w468, w459, IN7[2], w469, w470);
  FullAdder U22 (w470, w461, IN8[1], w471, w472);
  FullAdder U23 (w472, w462, IN9[0], w473, w474);
  HalfAdder U24 (w465, IN5[5], Out1[5], w476);
  FullAdder U25 (w476, w467, IN6[5], w477, w478);
  FullAdder U26 (w478, w469, IN7[3], w479, w480);
  FullAdder U27 (w480, w471, IN8[2], w481, w482);
  FullAdder U28 (w482, w473, IN9[1], w483, w484);
  FullAdder U29 (w484, w474, IN10[0], w485, w486);
  HalfAdder U30 (w477, IN6[6], Out1[6], w488);
  FullAdder U31 (w488, w479, IN7[4], w489, w490);
  FullAdder U32 (w490, w481, IN8[3], w491, w492);
  FullAdder U33 (w492, w483, IN9[2], w493, w494);
  FullAdder U34 (w494, w485, IN10[1], w495, w496);
  FullAdder U35 (w496, w486, IN11[0], w497, w498);
  HalfAdder U36 (w489, IN7[5], Out1[7], w500);
  FullAdder U37 (w500, w491, IN8[4], w501, w502);
  FullAdder U38 (w502, w493, IN9[3], w503, w504);
  FullAdder U39 (w504, w495, IN10[2], w505, w506);
  FullAdder U40 (w506, w497, IN11[1], w507, w508);
  FullAdder U41 (w508, w498, IN12[0], w509, w510);
  HalfAdder U42 (w501, IN8[5], Out1[8], w512);
  FullAdder U43 (w512, w503, IN9[4], w513, w514);
  FullAdder U44 (w514, w505, IN10[3], w515, w516);
  FullAdder U45 (w516, w507, IN11[2], w517, w518);
  FullAdder U46 (w518, w509, IN12[1], w519, w520);
  FullAdder U47 (w520, w510, IN13[0], w521, w522);
  HalfAdder U48 (w513, IN9[5], Out1[9], w524);
  FullAdder U49 (w524, w515, IN10[4], w525, w526);
  FullAdder U50 (w526, w517, IN11[3], w527, w528);
  FullAdder U51 (w528, w519, IN12[2], w529, w530);
  FullAdder U52 (w530, w521, IN13[1], w531, w532);
  FullAdder U53 (w532, w522, IN14[0], w533, w534);
  HalfAdder U54 (w525, IN10[5], Out1[10], w536);
  FullAdder U55 (w536, w527, IN11[4], w537, w538);
  FullAdder U56 (w538, w529, IN12[3], w539, w540);
  FullAdder U57 (w540, w531, IN13[2], w541, w542);
  FullAdder U58 (w542, w533, IN14[1], w543, w544);
  FullAdder U59 (w544, w534, IN15[0], w545, w546);
  HalfAdder U60 (w537, IN11[5], Out1[11], w548);
  FullAdder U61 (w548, w539, IN12[4], w549, w550);
  FullAdder U62 (w550, w541, IN13[3], w551, w552);
  FullAdder U63 (w552, w543, IN14[2], w553, w554);
  FullAdder U64 (w554, w545, IN15[1], w555, w556);
  FullAdder U65 (w556, w546, IN16[0], w557, w558);
  HalfAdder U66 (w549, IN12[5], Out1[12], w560);
  FullAdder U67 (w560, w551, IN13[4], w561, w562);
  FullAdder U68 (w562, w553, IN14[3], w563, w564);
  FullAdder U69 (w564, w555, IN15[2], w565, w566);
  FullAdder U70 (w566, w557, IN16[1], w567, w568);
  FullAdder U71 (w568, w558, IN17[0], w569, w570);
  HalfAdder U72 (w561, IN13[5], Out1[13], w572);
  FullAdder U73 (w572, w563, IN14[4], w573, w574);
  FullAdder U74 (w574, w565, IN15[3], w575, w576);
  FullAdder U75 (w576, w567, IN16[2], w577, w578);
  FullAdder U76 (w578, w569, IN17[1], w579, w580);
  FullAdder U77 (w580, w570, IN18[0], w581, w582);
  HalfAdder U78 (w573, IN14[5], Out1[14], w584);
  FullAdder U79 (w584, w575, IN15[4], w585, w586);
  FullAdder U80 (w586, w577, IN16[3], w587, w588);
  FullAdder U81 (w588, w579, IN17[2], w589, w590);
  FullAdder U82 (w590, w581, IN18[1], w591, w592);
  FullAdder U83 (w592, w582, IN19[0], w593, w594);
  HalfAdder U84 (w585, IN15[5], Out1[15], w596);
  FullAdder U85 (w596, w587, IN16[4], w597, w598);
  FullAdder U86 (w598, w589, IN17[3], w599, w600);
  FullAdder U87 (w600, w591, IN18[2], w601, w602);
  FullAdder U88 (w602, w593, IN19[1], w603, w604);
  FullAdder U89 (w604, w594, IN20[0], w605, w606);
  HalfAdder U90 (w597, IN16[5], Out1[16], w608);
  FullAdder U91 (w608, w599, IN17[4], w609, w610);
  FullAdder U92 (w610, w601, IN18[3], w611, w612);
  FullAdder U93 (w612, w603, IN19[2], w613, w614);
  FullAdder U94 (w614, w605, IN20[1], w615, w616);
  FullAdder U95 (w616, w606, IN21[0], w617, w618);
  HalfAdder U96 (w609, IN17[5], Out1[17], w620);
  FullAdder U97 (w620, w611, IN18[4], w621, w622);
  FullAdder U98 (w622, w613, IN19[3], w623, w624);
  FullAdder U99 (w624, w615, IN20[2], w625, w626);
  FullAdder U100 (w626, w617, IN21[1], w627, w628);
  FullAdder U101 (w628, w618, IN22[0], w629, w630);
  HalfAdder U102 (w621, IN18[5], Out1[18], w632);
  FullAdder U103 (w632, w623, IN19[4], w633, w634);
  FullAdder U104 (w634, w625, IN20[3], w635, w636);
  FullAdder U105 (w636, w627, IN21[2], w637, w638);
  FullAdder U106 (w638, w629, IN22[1], w639, w640);
  FullAdder U107 (w640, w630, IN23[0], w641, w642);
  HalfAdder U108 (w633, IN19[5], Out1[19], w644);
  FullAdder U109 (w644, w635, IN20[4], w645, w646);
  FullAdder U110 (w646, w637, IN21[3], w647, w648);
  FullAdder U111 (w648, w639, IN22[2], w649, w650);
  FullAdder U112 (w650, w641, IN23[1], w651, w652);
  FullAdder U113 (w652, w642, IN24[0], w653, w654);
  HalfAdder U114 (w645, IN20[5], Out1[20], w656);
  FullAdder U115 (w656, w647, IN21[4], w657, w658);
  FullAdder U116 (w658, w649, IN22[3], w659, w660);
  FullAdder U117 (w660, w651, IN23[2], w661, w662);
  FullAdder U118 (w662, w653, IN24[1], w663, w664);
  FullAdder U119 (w664, w654, IN25[0], w665, w666);
  HalfAdder U120 (w657, IN21[5], Out1[21], w668);
  FullAdder U121 (w668, w659, IN22[4], w669, w670);
  FullAdder U122 (w670, w661, IN23[3], w671, w672);
  FullAdder U123 (w672, w663, IN24[2], w673, w674);
  FullAdder U124 (w674, w665, IN25[1], w675, w676);
  FullAdder U125 (w676, w666, IN26[0], w677, w678);
  HalfAdder U126 (w669, IN22[5], Out1[22], w680);
  FullAdder U127 (w680, w671, IN23[4], w681, w682);
  FullAdder U128 (w682, w673, IN24[3], w683, w684);
  FullAdder U129 (w684, w675, IN25[2], w685, w686);
  FullAdder U130 (w686, w677, IN26[1], w687, w688);
  FullAdder U131 (w688, w678, IN27[0], w689, w690);
  HalfAdder U132 (w681, IN23[5], Out1[23], w692);
  FullAdder U133 (w692, w683, IN24[4], w693, w694);
  FullAdder U134 (w694, w685, IN25[3], w695, w696);
  FullAdder U135 (w696, w687, IN26[2], w697, w698);
  FullAdder U136 (w698, w689, IN27[1], w699, w700);
  FullAdder U137 (w700, w690, IN28[0], w701, w702);
  HalfAdder U138 (w693, IN24[5], Out1[24], w704);
  FullAdder U139 (w704, w695, IN25[4], w705, w706);
  FullAdder U140 (w706, w697, IN26[3], w707, w708);
  FullAdder U141 (w708, w699, IN27[2], w709, w710);
  FullAdder U142 (w710, w701, IN28[1], w711, w712);
  FullAdder U143 (w712, w702, IN29[0], w713, w714);
  HalfAdder U144 (w705, IN25[5], Out1[25], w716);
  FullAdder U145 (w716, w707, IN26[4], w717, w718);
  FullAdder U146 (w718, w709, IN27[3], w719, w720);
  FullAdder U147 (w720, w711, IN28[2], w721, w722);
  FullAdder U148 (w722, w713, IN29[1], w723, w724);
  FullAdder U149 (w724, w714, IN30[0], w725, w726);
  HalfAdder U150 (w717, IN26[5], Out1[26], w728);
  FullAdder U151 (w728, w719, IN27[4], w729, w730);
  FullAdder U152 (w730, w721, IN28[3], w731, w732);
  FullAdder U153 (w732, w723, IN29[2], w733, w734);
  FullAdder U154 (w734, w725, IN30[1], w735, w736);
  FullAdder U155 (w736, w726, IN31[0], w737, w738);
  HalfAdder U156 (w729, IN27[5], Out1[27], w740);
  FullAdder U157 (w740, w731, IN28[4], w741, w742);
  FullAdder U158 (w742, w733, IN29[3], w743, w744);
  FullAdder U159 (w744, w735, IN30[2], w745, w746);
  FullAdder U160 (w746, w737, IN31[1], w747, w748);
  FullAdder U161 (w748, w738, IN32[0], w749, w750);
  HalfAdder U162 (w741, IN28[5], Out1[28], w752);
  FullAdder U163 (w752, w743, IN29[4], w753, w754);
  FullAdder U164 (w754, w745, IN30[3], w755, w756);
  FullAdder U165 (w756, w747, IN31[2], w757, w758);
  FullAdder U166 (w758, w749, IN32[1], w759, w760);
  FullAdder U167 (w760, w750, IN33[0], w761, w762);
  HalfAdder U168 (w753, IN29[5], Out1[29], w764);
  FullAdder U169 (w764, w755, IN30[4], w765, w766);
  FullAdder U170 (w766, w757, IN31[3], w767, w768);
  FullAdder U171 (w768, w759, IN32[2], w769, w770);
  FullAdder U172 (w770, w761, IN33[1], w771, w772);
  FullAdder U173 (w772, w762, IN34[0], w773, w774);
  HalfAdder U174 (w765, IN30[5], Out1[30], w776);
  FullAdder U175 (w776, w767, IN31[4], w777, w778);
  FullAdder U176 (w778, w769, IN32[3], w779, w780);
  FullAdder U177 (w780, w771, IN33[2], w781, w782);
  FullAdder U178 (w782, w773, IN34[1], w783, w784);
  FullAdder U179 (w784, w774, IN35[0], w785, w786);
  HalfAdder U180 (w777, IN31[5], Out1[31], w788);
  FullAdder U181 (w788, w779, IN32[4], w789, w790);
  FullAdder U182 (w790, w781, IN33[3], w791, w792);
  FullAdder U183 (w792, w783, IN34[2], w793, w794);
  FullAdder U184 (w794, w785, IN35[1], w795, w796);
  FullAdder U185 (w796, w786, IN36[0], w797, w798);
  HalfAdder U186 (w789, IN32[5], Out1[32], w800);
  FullAdder U187 (w800, w791, IN33[4], w801, w802);
  FullAdder U188 (w802, w793, IN34[3], w803, w804);
  FullAdder U189 (w804, w795, IN35[2], w805, w806);
  FullAdder U190 (w806, w797, IN36[1], w807, w808);
  FullAdder U191 (w808, w798, IN37[0], w809, w810);
  HalfAdder U192 (w801, IN33[5], Out1[33], w812);
  FullAdder U193 (w812, w803, IN34[4], w813, w814);
  FullAdder U194 (w814, w805, IN35[3], w815, w816);
  FullAdder U195 (w816, w807, IN36[2], w817, w818);
  FullAdder U196 (w818, w809, IN37[1], w819, w820);
  FullAdder U197 (w820, w810, IN38[0], w821, w822);
  HalfAdder U198 (w813, IN34[5], Out1[34], w824);
  FullAdder U199 (w824, w815, IN35[4], w825, w826);
  FullAdder U200 (w826, w817, IN36[3], w827, w828);
  FullAdder U201 (w828, w819, IN37[2], w829, w830);
  FullAdder U202 (w830, w821, IN38[1], w831, w832);
  FullAdder U203 (w832, w822, IN39[0], w833, w834);
  HalfAdder U204 (w825, IN35[5], Out1[35], w836);
  FullAdder U205 (w836, w827, IN36[4], w837, w838);
  FullAdder U206 (w838, w829, IN37[3], w839, w840);
  FullAdder U207 (w840, w831, IN38[2], w841, w842);
  FullAdder U208 (w842, w833, IN39[1], w843, w844);
  FullAdder U209 (w844, w834, IN40[0], w845, w846);
  HalfAdder U210 (w837, IN36[5], Out1[36], w848);
  FullAdder U211 (w848, w839, IN37[4], w849, w850);
  FullAdder U212 (w850, w841, IN38[3], w851, w852);
  FullAdder U213 (w852, w843, IN39[2], w853, w854);
  FullAdder U214 (w854, w845, IN40[1], w855, w856);
  FullAdder U215 (w856, w846, IN41[0], w857, w858);
  HalfAdder U216 (w849, IN37[5], Out1[37], w860);
  FullAdder U217 (w860, w851, IN38[4], w861, w862);
  FullAdder U218 (w862, w853, IN39[3], w863, w864);
  FullAdder U219 (w864, w855, IN40[2], w865, w866);
  FullAdder U220 (w866, w857, IN41[1], w867, w868);
  FullAdder U221 (w868, w858, IN42[0], w869, w870);
  HalfAdder U222 (w861, IN38[5], Out1[38], w872);
  FullAdder U223 (w872, w863, IN39[4], w873, w874);
  FullAdder U224 (w874, w865, IN40[3], w875, w876);
  FullAdder U225 (w876, w867, IN41[2], w877, w878);
  FullAdder U226 (w878, w869, IN42[1], w879, w880);
  FullAdder U227 (w880, w870, IN43[0], w881, w882);
  HalfAdder U228 (w873, IN39[5], Out1[39], w884);
  FullAdder U229 (w884, w875, IN40[4], w885, w886);
  FullAdder U230 (w886, w877, IN41[3], w887, w888);
  FullAdder U231 (w888, w879, IN42[2], w889, w890);
  FullAdder U232 (w890, w881, IN43[1], w891, w892);
  FullAdder U233 (w892, w882, IN44[0], w893, w894);
  HalfAdder U234 (w885, IN40[5], Out1[40], w896);
  FullAdder U235 (w896, w887, IN41[4], w897, w898);
  FullAdder U236 (w898, w889, IN42[3], w899, w900);
  FullAdder U237 (w900, w891, IN43[2], w901, w902);
  FullAdder U238 (w902, w893, IN44[1], w903, w904);
  FullAdder U239 (w904, w894, IN45[0], w905, w906);
  HalfAdder U240 (w897, IN41[5], Out1[41], w908);
  FullAdder U241 (w908, w899, IN42[4], w909, w910);
  FullAdder U242 (w910, w901, IN43[3], w911, w912);
  FullAdder U243 (w912, w903, IN44[2], w913, w914);
  FullAdder U244 (w914, w905, IN45[1], w915, w916);
  FullAdder U245 (w916, w906, IN46[0], w917, w918);
  HalfAdder U246 (w909, IN42[5], Out1[42], w920);
  FullAdder U247 (w920, w911, IN43[4], w921, w922);
  FullAdder U248 (w922, w913, IN44[3], w923, w924);
  FullAdder U249 (w924, w915, IN45[2], w925, w926);
  FullAdder U250 (w926, w917, IN46[1], w927, w928);
  FullAdder U251 (w928, w918, IN47[0], w929, w930);
  HalfAdder U252 (w921, IN43[5], Out1[43], w932);
  FullAdder U253 (w932, w923, IN44[4], w933, w934);
  FullAdder U254 (w934, w925, IN45[3], w935, w936);
  FullAdder U255 (w936, w927, IN46[2], w937, w938);
  FullAdder U256 (w938, w929, IN47[1], w939, w940);
  FullAdder U257 (w940, w930, IN48[0], w941, w942);
  HalfAdder U258 (w933, IN44[5], Out1[44], w944);
  FullAdder U259 (w944, w935, IN45[4], w945, w946);
  FullAdder U260 (w946, w937, IN46[3], w947, w948);
  FullAdder U261 (w948, w939, IN47[2], w949, w950);
  FullAdder U262 (w950, w941, IN48[1], w951, w952);
  FullAdder U263 (w952, w942, IN49[0], w953, w954);
  HalfAdder U264 (w945, IN45[5], Out1[45], w956);
  FullAdder U265 (w956, w947, IN46[4], w957, w958);
  FullAdder U266 (w958, w949, IN47[3], w959, w960);
  FullAdder U267 (w960, w951, IN48[2], w961, w962);
  FullAdder U268 (w962, w953, IN49[1], w963, w964);
  FullAdder U269 (w964, w954, IN50[0], w965, w966);
  HalfAdder U270 (w957, IN46[5], Out1[46], w968);
  FullAdder U271 (w968, w959, IN47[4], w969, w970);
  FullAdder U272 (w970, w961, IN48[3], w971, w972);
  FullAdder U273 (w972, w963, IN49[2], w973, w974);
  FullAdder U274 (w974, w965, IN50[1], w975, w976);
  FullAdder U275 (w976, w966, IN51[0], w977, w978);
  HalfAdder U276 (w969, IN47[5], Out1[47], w980);
  FullAdder U277 (w980, w971, IN48[4], w981, w982);
  FullAdder U278 (w982, w973, IN49[3], w983, w984);
  FullAdder U279 (w984, w975, IN50[2], w985, w986);
  FullAdder U280 (w986, w977, IN51[1], w987, w988);
  FullAdder U281 (w988, w978, IN52[0], w989, w990);
  HalfAdder U282 (w981, IN48[5], Out1[48], w992);
  FullAdder U283 (w992, w983, IN49[4], w993, w994);
  FullAdder U284 (w994, w985, IN50[3], w995, w996);
  FullAdder U285 (w996, w987, IN51[2], w997, w998);
  FullAdder U286 (w998, w989, IN52[1], w999, w1000);
  FullAdder U287 (w1000, w990, IN53[0], w1001, w1002);
  HalfAdder U288 (w993, IN49[5], Out1[49], w1004);
  FullAdder U289 (w1004, w995, IN50[4], w1005, w1006);
  FullAdder U290 (w1006, w997, IN51[3], w1007, w1008);
  FullAdder U291 (w1008, w999, IN52[2], w1009, w1010);
  FullAdder U292 (w1010, w1001, IN53[1], w1011, w1012);
  FullAdder U293 (w1012, w1002, IN54[0], w1013, w1014);
  HalfAdder U294 (w1005, IN50[5], Out1[50], w1016);
  FullAdder U295 (w1016, w1007, IN51[4], w1017, w1018);
  FullAdder U296 (w1018, w1009, IN52[3], w1019, w1020);
  FullAdder U297 (w1020, w1011, IN53[2], w1021, w1022);
  FullAdder U298 (w1022, w1013, IN54[1], w1023, w1024);
  FullAdder U299 (w1024, w1014, IN55[0], w1025, w1026);
  HalfAdder U300 (w1017, IN51[5], Out1[51], w1028);
  FullAdder U301 (w1028, w1019, IN52[4], w1029, w1030);
  FullAdder U302 (w1030, w1021, IN53[3], w1031, w1032);
  FullAdder U303 (w1032, w1023, IN54[2], w1033, w1034);
  FullAdder U304 (w1034, w1025, IN55[1], w1035, w1036);
  FullAdder U305 (w1036, w1026, IN56[0], w1037, w1038);
  HalfAdder U306 (w1029, IN52[5], Out1[52], w1040);
  FullAdder U307 (w1040, w1031, IN53[4], w1041, w1042);
  FullAdder U308 (w1042, w1033, IN54[3], w1043, w1044);
  FullAdder U309 (w1044, w1035, IN55[2], w1045, w1046);
  FullAdder U310 (w1046, w1037, IN56[1], w1047, w1048);
  FullAdder U311 (w1048, w1038, IN57[0], w1049, w1050);
  HalfAdder U312 (w1041, IN53[5], Out1[53], w1052);
  FullAdder U313 (w1052, w1043, IN54[4], w1053, w1054);
  FullAdder U314 (w1054, w1045, IN55[3], w1055, w1056);
  FullAdder U315 (w1056, w1047, IN56[2], w1057, w1058);
  FullAdder U316 (w1058, w1049, IN57[1], w1059, w1060);
  FullAdder U317 (w1060, w1050, IN58[0], w1061, w1062);
  HalfAdder U318 (w1053, IN54[5], Out1[54], w1064);
  FullAdder U319 (w1064, w1055, IN55[4], w1065, w1066);
  FullAdder U320 (w1066, w1057, IN56[3], w1067, w1068);
  FullAdder U321 (w1068, w1059, IN57[2], w1069, w1070);
  FullAdder U322 (w1070, w1061, IN58[1], w1071, w1072);
  FullAdder U323 (w1072, w1062, IN59[0], w1073, w1074);
  HalfAdder U324 (w1065, IN55[5], Out1[55], w1076);
  FullAdder U325 (w1076, w1067, IN56[4], w1077, w1078);
  FullAdder U326 (w1078, w1069, IN57[3], w1079, w1080);
  FullAdder U327 (w1080, w1071, IN58[2], w1081, w1082);
  FullAdder U328 (w1082, w1073, IN59[1], w1083, w1084);
  FullAdder U329 (w1084, w1074, IN60[0], w1085, w1086);
  HalfAdder U330 (w1077, IN56[5], Out1[56], w1088);
  FullAdder U331 (w1088, w1079, IN57[4], w1089, w1090);
  FullAdder U332 (w1090, w1081, IN58[3], w1091, w1092);
  FullAdder U333 (w1092, w1083, IN59[2], w1093, w1094);
  FullAdder U334 (w1094, w1085, IN60[1], w1095, w1096);
  FullAdder U335 (w1096, w1086, IN61[0], w1097, w1098);
  HalfAdder U336 (w1089, IN57[5], Out1[57], w1100);
  FullAdder U337 (w1100, w1091, IN58[4], w1101, w1102);
  FullAdder U338 (w1102, w1093, IN59[3], w1103, w1104);
  FullAdder U339 (w1104, w1095, IN60[2], w1105, w1106);
  FullAdder U340 (w1106, w1097, IN61[1], w1107, w1108);
  FullAdder U341 (w1108, w1098, IN62[0], w1109, w1110);
  HalfAdder U342 (w1101, IN58[5], Out1[58], w1112);
  FullAdder U343 (w1112, w1103, IN59[4], w1113, w1114);
  FullAdder U344 (w1114, w1105, IN60[3], w1115, w1116);
  FullAdder U345 (w1116, w1107, IN61[2], w1117, w1118);
  FullAdder U346 (w1118, w1109, IN62[1], w1119, w1120);
  FullAdder U347 (w1120, w1110, IN63[0], w1121, w1122);
  HalfAdder U348 (w1113, IN59[5], Out1[59], w1124);
  FullAdder U349 (w1124, w1115, IN60[4], w1125, w1126);
  FullAdder U350 (w1126, w1117, IN61[3], w1127, w1128);
  FullAdder U351 (w1128, w1119, IN62[2], w1129, w1130);
  FullAdder U352 (w1130, w1121, IN63[1], w1131, w1132);
  FullAdder U353 (w1132, w1122, IN64[0], w1133, w1134);
  HalfAdder U354 (w1125, IN60[5], Out1[60], w1136);
  FullAdder U355 (w1136, w1127, IN61[4], Out1[61], w1138);
  FullAdder U356 (w1138, w1129, IN62[3], Out1[62], w1140);
  FullAdder U357 (w1140, w1131, IN63[2], Out1[63], w1142);
  FullAdder U358 (w1142, w1133, IN64[1], Out1[64], w1144);
  FullAdder U359 (w1144, w1134, IN65[0], Out1[65], Out1[66]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN7[6];
  assign Out2[1] = IN8[6];
  assign Out2[2] = IN9[6];
  assign Out2[3] = IN10[6];
  assign Out2[4] = IN11[6];
  assign Out2[5] = IN12[6];
  assign Out2[6] = IN13[6];
  assign Out2[7] = IN14[6];
  assign Out2[8] = IN15[6];
  assign Out2[9] = IN16[6];
  assign Out2[10] = IN17[6];
  assign Out2[11] = IN18[6];
  assign Out2[12] = IN19[6];
  assign Out2[13] = IN20[6];
  assign Out2[14] = IN21[6];
  assign Out2[15] = IN22[6];
  assign Out2[16] = IN23[6];
  assign Out2[17] = IN24[6];
  assign Out2[18] = IN25[6];
  assign Out2[19] = IN26[6];
  assign Out2[20] = IN27[6];
  assign Out2[21] = IN28[6];
  assign Out2[22] = IN29[6];
  assign Out2[23] = IN30[6];
  assign Out2[24] = IN31[6];
  assign Out2[25] = IN32[6];
  assign Out2[26] = IN33[6];
  assign Out2[27] = IN34[6];
  assign Out2[28] = IN35[6];
  assign Out2[29] = IN36[6];
  assign Out2[30] = IN37[6];
  assign Out2[31] = IN38[6];
  assign Out2[32] = IN39[6];
  assign Out2[33] = IN40[6];
  assign Out2[34] = IN41[6];
  assign Out2[35] = IN42[6];
  assign Out2[36] = IN43[6];
  assign Out2[37] = IN44[6];
  assign Out2[38] = IN45[6];
  assign Out2[39] = IN46[6];
  assign Out2[40] = IN47[6];
  assign Out2[41] = IN48[6];
  assign Out2[42] = IN49[6];
  assign Out2[43] = IN50[6];
  assign Out2[44] = IN51[6];
  assign Out2[45] = IN52[6];
  assign Out2[46] = IN53[6];
  assign Out2[47] = IN54[6];
  assign Out2[48] = IN55[6];
  assign Out2[49] = IN56[6];
  assign Out2[50] = IN57[6];
  assign Out2[51] = IN58[6];
  assign Out2[52] = IN59[6];
  assign Out2[53] = IN60[6];
  assign Out2[54] = IN61[5];
  assign Out2[55] = IN62[4];
  assign Out2[56] = IN63[3];
  assign Out2[57] = IN64[2];
  assign Out2[58] = IN65[1];
  assign Out2[59] = IN66[0];

endmodule
module RC_60_60(IN1, IN2, Out);
  input [59:0] IN1;
  input [59:0] IN2;
  output [60:0] Out;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  wire w231;
  wire w233;
  wire w235;
  wire w237;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w121);
  FullAdder U1 (IN1[1], IN2[1], w121, Out[1], w123);
  FullAdder U2 (IN1[2], IN2[2], w123, Out[2], w125);
  FullAdder U3 (IN1[3], IN2[3], w125, Out[3], w127);
  FullAdder U4 (IN1[4], IN2[4], w127, Out[4], w129);
  FullAdder U5 (IN1[5], IN2[5], w129, Out[5], w131);
  FullAdder U6 (IN1[6], IN2[6], w131, Out[6], w133);
  FullAdder U7 (IN1[7], IN2[7], w133, Out[7], w135);
  FullAdder U8 (IN1[8], IN2[8], w135, Out[8], w137);
  FullAdder U9 (IN1[9], IN2[9], w137, Out[9], w139);
  FullAdder U10 (IN1[10], IN2[10], w139, Out[10], w141);
  FullAdder U11 (IN1[11], IN2[11], w141, Out[11], w143);
  FullAdder U12 (IN1[12], IN2[12], w143, Out[12], w145);
  FullAdder U13 (IN1[13], IN2[13], w145, Out[13], w147);
  FullAdder U14 (IN1[14], IN2[14], w147, Out[14], w149);
  FullAdder U15 (IN1[15], IN2[15], w149, Out[15], w151);
  FullAdder U16 (IN1[16], IN2[16], w151, Out[16], w153);
  FullAdder U17 (IN1[17], IN2[17], w153, Out[17], w155);
  FullAdder U18 (IN1[18], IN2[18], w155, Out[18], w157);
  FullAdder U19 (IN1[19], IN2[19], w157, Out[19], w159);
  FullAdder U20 (IN1[20], IN2[20], w159, Out[20], w161);
  FullAdder U21 (IN1[21], IN2[21], w161, Out[21], w163);
  FullAdder U22 (IN1[22], IN2[22], w163, Out[22], w165);
  FullAdder U23 (IN1[23], IN2[23], w165, Out[23], w167);
  FullAdder U24 (IN1[24], IN2[24], w167, Out[24], w169);
  FullAdder U25 (IN1[25], IN2[25], w169, Out[25], w171);
  FullAdder U26 (IN1[26], IN2[26], w171, Out[26], w173);
  FullAdder U27 (IN1[27], IN2[27], w173, Out[27], w175);
  FullAdder U28 (IN1[28], IN2[28], w175, Out[28], w177);
  FullAdder U29 (IN1[29], IN2[29], w177, Out[29], w179);
  FullAdder U30 (IN1[30], IN2[30], w179, Out[30], w181);
  FullAdder U31 (IN1[31], IN2[31], w181, Out[31], w183);
  FullAdder U32 (IN1[32], IN2[32], w183, Out[32], w185);
  FullAdder U33 (IN1[33], IN2[33], w185, Out[33], w187);
  FullAdder U34 (IN1[34], IN2[34], w187, Out[34], w189);
  FullAdder U35 (IN1[35], IN2[35], w189, Out[35], w191);
  FullAdder U36 (IN1[36], IN2[36], w191, Out[36], w193);
  FullAdder U37 (IN1[37], IN2[37], w193, Out[37], w195);
  FullAdder U38 (IN1[38], IN2[38], w195, Out[38], w197);
  FullAdder U39 (IN1[39], IN2[39], w197, Out[39], w199);
  FullAdder U40 (IN1[40], IN2[40], w199, Out[40], w201);
  FullAdder U41 (IN1[41], IN2[41], w201, Out[41], w203);
  FullAdder U42 (IN1[42], IN2[42], w203, Out[42], w205);
  FullAdder U43 (IN1[43], IN2[43], w205, Out[43], w207);
  FullAdder U44 (IN1[44], IN2[44], w207, Out[44], w209);
  FullAdder U45 (IN1[45], IN2[45], w209, Out[45], w211);
  FullAdder U46 (IN1[46], IN2[46], w211, Out[46], w213);
  FullAdder U47 (IN1[47], IN2[47], w213, Out[47], w215);
  FullAdder U48 (IN1[48], IN2[48], w215, Out[48], w217);
  FullAdder U49 (IN1[49], IN2[49], w217, Out[49], w219);
  FullAdder U50 (IN1[50], IN2[50], w219, Out[50], w221);
  FullAdder U51 (IN1[51], IN2[51], w221, Out[51], w223);
  FullAdder U52 (IN1[52], IN2[52], w223, Out[52], w225);
  FullAdder U53 (IN1[53], IN2[53], w225, Out[53], w227);
  FullAdder U54 (IN1[54], IN2[54], w227, Out[54], w229);
  FullAdder U55 (IN1[55], IN2[55], w229, Out[55], w231);
  FullAdder U56 (IN1[56], IN2[56], w231, Out[56], w233);
  FullAdder U57 (IN1[57], IN2[57], w233, Out[57], w235);
  FullAdder U58 (IN1[58], IN2[58], w235, Out[58], w237);
  FullAdder U59 (IN1[59], IN2[59], w237, Out[59], Out[60]);

endmodule
module NR_7_61(IN1, IN2, Out);
  input [6:0] IN1;
  input [60:0] IN2;
  output [67:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [6:0] P37;
  wire [6:0] P38;
  wire [6:0] P39;
  wire [6:0] P40;
  wire [6:0] P41;
  wire [6:0] P42;
  wire [6:0] P43;
  wire [6:0] P44;
  wire [6:0] P45;
  wire [6:0] P46;
  wire [6:0] P47;
  wire [6:0] P48;
  wire [6:0] P49;
  wire [6:0] P50;
  wire [6:0] P51;
  wire [6:0] P52;
  wire [6:0] P53;
  wire [6:0] P54;
  wire [6:0] P55;
  wire [6:0] P56;
  wire [6:0] P57;
  wire [6:0] P58;
  wire [6:0] P59;
  wire [6:0] P60;
  wire [5:0] P61;
  wire [4:0] P62;
  wire [3:0] P63;
  wire [2:0] P64;
  wire [1:0] P65;
  wire [0:0] P66;
  wire [66:0] R1;
  wire [59:0] R2;
  wire [67:0] aOut;
  U_SP_7_61 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, R1, R2);
  RC_60_60 S2 (R1[66:7], R2, aOut[67:7]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign Out = aOut[67:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
