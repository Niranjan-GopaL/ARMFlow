//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 14
  second input length: 49
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_14_49(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61);
  input [13:0] IN1;
  input [48:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [13:0] P14;
  output [13:0] P15;
  output [13:0] P16;
  output [13:0] P17;
  output [13:0] P18;
  output [13:0] P19;
  output [13:0] P20;
  output [13:0] P21;
  output [13:0] P22;
  output [13:0] P23;
  output [13:0] P24;
  output [13:0] P25;
  output [13:0] P26;
  output [13:0] P27;
  output [13:0] P28;
  output [13:0] P29;
  output [13:0] P30;
  output [13:0] P31;
  output [13:0] P32;
  output [13:0] P33;
  output [13:0] P34;
  output [13:0] P35;
  output [13:0] P36;
  output [13:0] P37;
  output [13:0] P38;
  output [13:0] P39;
  output [13:0] P40;
  output [13:0] P41;
  output [13:0] P42;
  output [13:0] P43;
  output [13:0] P44;
  output [13:0] P45;
  output [13:0] P46;
  output [13:0] P47;
  output [13:0] P48;
  output [12:0] P49;
  output [11:0] P50;
  output [10:0] P51;
  output [9:0] P52;
  output [8:0] P53;
  output [7:0] P54;
  output [6:0] P55;
  output [5:0] P56;
  output [4:0] P57;
  output [3:0] P58;
  output [2:0] P59;
  output [1:0] P60;
  output [0:0] P61;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[0] = IN1[1]&IN2[48];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[1] = IN1[2]&IN2[47];
  assign P50[0] = IN1[2]&IN2[48];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[2] = IN1[3]&IN2[46];
  assign P50[1] = IN1[3]&IN2[47];
  assign P51[0] = IN1[3]&IN2[48];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[3] = IN1[4]&IN2[45];
  assign P50[2] = IN1[4]&IN2[46];
  assign P51[1] = IN1[4]&IN2[47];
  assign P52[0] = IN1[4]&IN2[48];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[4] = IN1[5]&IN2[44];
  assign P50[3] = IN1[5]&IN2[45];
  assign P51[2] = IN1[5]&IN2[46];
  assign P52[1] = IN1[5]&IN2[47];
  assign P53[0] = IN1[5]&IN2[48];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[5] = IN1[6]&IN2[43];
  assign P50[4] = IN1[6]&IN2[44];
  assign P51[3] = IN1[6]&IN2[45];
  assign P52[2] = IN1[6]&IN2[46];
  assign P53[1] = IN1[6]&IN2[47];
  assign P54[0] = IN1[6]&IN2[48];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[6] = IN1[7]&IN2[42];
  assign P50[5] = IN1[7]&IN2[43];
  assign P51[4] = IN1[7]&IN2[44];
  assign P52[3] = IN1[7]&IN2[45];
  assign P53[2] = IN1[7]&IN2[46];
  assign P54[1] = IN1[7]&IN2[47];
  assign P55[0] = IN1[7]&IN2[48];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[7] = IN1[8]&IN2[41];
  assign P50[6] = IN1[8]&IN2[42];
  assign P51[5] = IN1[8]&IN2[43];
  assign P52[4] = IN1[8]&IN2[44];
  assign P53[3] = IN1[8]&IN2[45];
  assign P54[2] = IN1[8]&IN2[46];
  assign P55[1] = IN1[8]&IN2[47];
  assign P56[0] = IN1[8]&IN2[48];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[8] = IN1[9]&IN2[40];
  assign P50[7] = IN1[9]&IN2[41];
  assign P51[6] = IN1[9]&IN2[42];
  assign P52[5] = IN1[9]&IN2[43];
  assign P53[4] = IN1[9]&IN2[44];
  assign P54[3] = IN1[9]&IN2[45];
  assign P55[2] = IN1[9]&IN2[46];
  assign P56[1] = IN1[9]&IN2[47];
  assign P57[0] = IN1[9]&IN2[48];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[9] = IN1[10]&IN2[39];
  assign P50[8] = IN1[10]&IN2[40];
  assign P51[7] = IN1[10]&IN2[41];
  assign P52[6] = IN1[10]&IN2[42];
  assign P53[5] = IN1[10]&IN2[43];
  assign P54[4] = IN1[10]&IN2[44];
  assign P55[3] = IN1[10]&IN2[45];
  assign P56[2] = IN1[10]&IN2[46];
  assign P57[1] = IN1[10]&IN2[47];
  assign P58[0] = IN1[10]&IN2[48];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[10] = IN1[11]&IN2[38];
  assign P50[9] = IN1[11]&IN2[39];
  assign P51[8] = IN1[11]&IN2[40];
  assign P52[7] = IN1[11]&IN2[41];
  assign P53[6] = IN1[11]&IN2[42];
  assign P54[5] = IN1[11]&IN2[43];
  assign P55[4] = IN1[11]&IN2[44];
  assign P56[3] = IN1[11]&IN2[45];
  assign P57[2] = IN1[11]&IN2[46];
  assign P58[1] = IN1[11]&IN2[47];
  assign P59[0] = IN1[11]&IN2[48];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[11] = IN1[12]&IN2[37];
  assign P50[10] = IN1[12]&IN2[38];
  assign P51[9] = IN1[12]&IN2[39];
  assign P52[8] = IN1[12]&IN2[40];
  assign P53[7] = IN1[12]&IN2[41];
  assign P54[6] = IN1[12]&IN2[42];
  assign P55[5] = IN1[12]&IN2[43];
  assign P56[4] = IN1[12]&IN2[44];
  assign P57[3] = IN1[12]&IN2[45];
  assign P58[2] = IN1[12]&IN2[46];
  assign P59[1] = IN1[12]&IN2[47];
  assign P60[0] = IN1[12]&IN2[48];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[12] = IN1[13]&IN2[36];
  assign P50[11] = IN1[13]&IN2[37];
  assign P51[10] = IN1[13]&IN2[38];
  assign P52[9] = IN1[13]&IN2[39];
  assign P53[8] = IN1[13]&IN2[40];
  assign P54[7] = IN1[13]&IN2[41];
  assign P55[6] = IN1[13]&IN2[42];
  assign P56[5] = IN1[13]&IN2[43];
  assign P57[4] = IN1[13]&IN2[44];
  assign P58[3] = IN1[13]&IN2[45];
  assign P59[2] = IN1[13]&IN2[46];
  assign P60[1] = IN1[13]&IN2[47];
  assign P61[0] = IN1[13]&IN2[48];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [13:0] IN14;
  input [13:0] IN15;
  input [13:0] IN16;
  input [13:0] IN17;
  input [13:0] IN18;
  input [13:0] IN19;
  input [13:0] IN20;
  input [13:0] IN21;
  input [13:0] IN22;
  input [13:0] IN23;
  input [13:0] IN24;
  input [13:0] IN25;
  input [13:0] IN26;
  input [13:0] IN27;
  input [13:0] IN28;
  input [13:0] IN29;
  input [13:0] IN30;
  input [13:0] IN31;
  input [13:0] IN32;
  input [13:0] IN33;
  input [13:0] IN34;
  input [13:0] IN35;
  input [13:0] IN36;
  input [13:0] IN37;
  input [13:0] IN38;
  input [13:0] IN39;
  input [13:0] IN40;
  input [13:0] IN41;
  input [13:0] IN42;
  input [13:0] IN43;
  input [13:0] IN44;
  input [13:0] IN45;
  input [13:0] IN46;
  input [13:0] IN47;
  input [13:0] IN48;
  input [12:0] IN49;
  input [11:0] IN50;
  input [10:0] IN51;
  input [9:0] IN52;
  input [8:0] IN53;
  input [7:0] IN54;
  input [6:0] IN55;
  input [5:0] IN56;
  input [4:0] IN57;
  input [3:0] IN58;
  input [2:0] IN59;
  input [1:0] IN60;
  input [0:0] IN61;
  output [61:0] Out1;
  output [47:0] Out2;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1126;
  wire w1127;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1192;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1214;
  wire w1215;
  wire w1216;
  wire w1217;
  wire w1218;
  wire w1219;
  wire w1220;
  wire w1221;
  wire w1222;
  wire w1223;
  wire w1224;
  wire w1225;
  wire w1226;
  wire w1227;
  wire w1228;
  wire w1229;
  wire w1230;
  wire w1231;
  wire w1233;
  wire w1234;
  wire w1235;
  wire w1236;
  wire w1237;
  wire w1238;
  wire w1239;
  wire w1240;
  wire w1241;
  wire w1242;
  wire w1243;
  wire w1244;
  wire w1245;
  wire w1246;
  wire w1247;
  wire w1248;
  wire w1249;
  wire w1250;
  wire w1251;
  wire w1252;
  wire w1253;
  wire w1254;
  wire w1255;
  wire w1256;
  wire w1257;
  wire w1259;
  wire w1260;
  wire w1261;
  wire w1262;
  wire w1263;
  wire w1264;
  wire w1265;
  wire w1266;
  wire w1267;
  wire w1268;
  wire w1269;
  wire w1270;
  wire w1271;
  wire w1272;
  wire w1273;
  wire w1274;
  wire w1275;
  wire w1276;
  wire w1277;
  wire w1278;
  wire w1279;
  wire w1280;
  wire w1281;
  wire w1282;
  wire w1283;
  wire w1285;
  wire w1286;
  wire w1287;
  wire w1288;
  wire w1289;
  wire w1290;
  wire w1291;
  wire w1292;
  wire w1293;
  wire w1294;
  wire w1295;
  wire w1296;
  wire w1297;
  wire w1298;
  wire w1299;
  wire w1300;
  wire w1301;
  wire w1302;
  wire w1303;
  wire w1304;
  wire w1305;
  wire w1306;
  wire w1307;
  wire w1308;
  wire w1309;
  wire w1311;
  wire w1312;
  wire w1313;
  wire w1314;
  wire w1315;
  wire w1316;
  wire w1317;
  wire w1318;
  wire w1319;
  wire w1320;
  wire w1321;
  wire w1322;
  wire w1323;
  wire w1324;
  wire w1325;
  wire w1326;
  wire w1327;
  wire w1328;
  wire w1329;
  wire w1330;
  wire w1331;
  wire w1332;
  wire w1333;
  wire w1334;
  wire w1335;
  wire w1337;
  wire w1338;
  wire w1339;
  wire w1340;
  wire w1341;
  wire w1342;
  wire w1343;
  wire w1344;
  wire w1345;
  wire w1346;
  wire w1347;
  wire w1348;
  wire w1349;
  wire w1350;
  wire w1351;
  wire w1352;
  wire w1353;
  wire w1354;
  wire w1355;
  wire w1356;
  wire w1357;
  wire w1358;
  wire w1359;
  wire w1360;
  wire w1361;
  wire w1363;
  wire w1364;
  wire w1365;
  wire w1366;
  wire w1367;
  wire w1368;
  wire w1369;
  wire w1370;
  wire w1371;
  wire w1372;
  wire w1373;
  wire w1374;
  wire w1375;
  wire w1376;
  wire w1377;
  wire w1378;
  wire w1379;
  wire w1380;
  wire w1381;
  wire w1382;
  wire w1383;
  wire w1384;
  wire w1385;
  wire w1386;
  wire w1387;
  wire w1389;
  wire w1390;
  wire w1391;
  wire w1392;
  wire w1393;
  wire w1394;
  wire w1395;
  wire w1396;
  wire w1397;
  wire w1398;
  wire w1399;
  wire w1400;
  wire w1401;
  wire w1402;
  wire w1403;
  wire w1404;
  wire w1405;
  wire w1406;
  wire w1407;
  wire w1408;
  wire w1409;
  wire w1410;
  wire w1411;
  wire w1412;
  wire w1413;
  wire w1415;
  wire w1416;
  wire w1417;
  wire w1418;
  wire w1419;
  wire w1420;
  wire w1421;
  wire w1422;
  wire w1423;
  wire w1424;
  wire w1425;
  wire w1426;
  wire w1427;
  wire w1428;
  wire w1429;
  wire w1430;
  wire w1431;
  wire w1432;
  wire w1433;
  wire w1434;
  wire w1435;
  wire w1436;
  wire w1437;
  wire w1438;
  wire w1439;
  wire w1441;
  wire w1442;
  wire w1443;
  wire w1444;
  wire w1445;
  wire w1446;
  wire w1447;
  wire w1448;
  wire w1449;
  wire w1450;
  wire w1451;
  wire w1452;
  wire w1453;
  wire w1454;
  wire w1455;
  wire w1456;
  wire w1457;
  wire w1458;
  wire w1459;
  wire w1460;
  wire w1461;
  wire w1462;
  wire w1463;
  wire w1464;
  wire w1465;
  wire w1467;
  wire w1468;
  wire w1469;
  wire w1470;
  wire w1471;
  wire w1472;
  wire w1473;
  wire w1474;
  wire w1475;
  wire w1476;
  wire w1477;
  wire w1478;
  wire w1479;
  wire w1480;
  wire w1481;
  wire w1482;
  wire w1483;
  wire w1484;
  wire w1485;
  wire w1486;
  wire w1487;
  wire w1488;
  wire w1489;
  wire w1490;
  wire w1491;
  wire w1493;
  wire w1494;
  wire w1495;
  wire w1496;
  wire w1497;
  wire w1498;
  wire w1499;
  wire w1500;
  wire w1501;
  wire w1502;
  wire w1503;
  wire w1504;
  wire w1505;
  wire w1506;
  wire w1507;
  wire w1508;
  wire w1509;
  wire w1510;
  wire w1511;
  wire w1512;
  wire w1513;
  wire w1514;
  wire w1515;
  wire w1516;
  wire w1517;
  wire w1519;
  wire w1520;
  wire w1521;
  wire w1522;
  wire w1523;
  wire w1524;
  wire w1525;
  wire w1526;
  wire w1527;
  wire w1528;
  wire w1529;
  wire w1530;
  wire w1531;
  wire w1532;
  wire w1533;
  wire w1534;
  wire w1535;
  wire w1536;
  wire w1537;
  wire w1538;
  wire w1539;
  wire w1540;
  wire w1541;
  wire w1542;
  wire w1543;
  wire w1545;
  wire w1546;
  wire w1547;
  wire w1548;
  wire w1549;
  wire w1550;
  wire w1551;
  wire w1552;
  wire w1553;
  wire w1554;
  wire w1555;
  wire w1556;
  wire w1557;
  wire w1558;
  wire w1559;
  wire w1560;
  wire w1561;
  wire w1562;
  wire w1563;
  wire w1564;
  wire w1565;
  wire w1566;
  wire w1567;
  wire w1568;
  wire w1569;
  wire w1571;
  wire w1572;
  wire w1573;
  wire w1574;
  wire w1575;
  wire w1576;
  wire w1577;
  wire w1578;
  wire w1579;
  wire w1580;
  wire w1581;
  wire w1582;
  wire w1583;
  wire w1584;
  wire w1585;
  wire w1586;
  wire w1587;
  wire w1588;
  wire w1589;
  wire w1590;
  wire w1591;
  wire w1592;
  wire w1593;
  wire w1594;
  wire w1595;
  wire w1597;
  wire w1598;
  wire w1599;
  wire w1600;
  wire w1601;
  wire w1602;
  wire w1603;
  wire w1604;
  wire w1605;
  wire w1606;
  wire w1607;
  wire w1608;
  wire w1609;
  wire w1610;
  wire w1611;
  wire w1612;
  wire w1613;
  wire w1614;
  wire w1615;
  wire w1616;
  wire w1617;
  wire w1618;
  wire w1619;
  wire w1620;
  wire w1621;
  wire w1623;
  wire w1624;
  wire w1625;
  wire w1626;
  wire w1627;
  wire w1628;
  wire w1629;
  wire w1630;
  wire w1631;
  wire w1632;
  wire w1633;
  wire w1634;
  wire w1635;
  wire w1636;
  wire w1637;
  wire w1638;
  wire w1639;
  wire w1640;
  wire w1641;
  wire w1642;
  wire w1643;
  wire w1644;
  wire w1645;
  wire w1646;
  wire w1647;
  wire w1649;
  wire w1650;
  wire w1651;
  wire w1652;
  wire w1653;
  wire w1654;
  wire w1655;
  wire w1656;
  wire w1657;
  wire w1658;
  wire w1659;
  wire w1660;
  wire w1661;
  wire w1662;
  wire w1663;
  wire w1664;
  wire w1665;
  wire w1666;
  wire w1667;
  wire w1668;
  wire w1669;
  wire w1670;
  wire w1671;
  wire w1672;
  wire w1673;
  wire w1675;
  wire w1676;
  wire w1677;
  wire w1678;
  wire w1679;
  wire w1680;
  wire w1681;
  wire w1682;
  wire w1683;
  wire w1684;
  wire w1685;
  wire w1686;
  wire w1687;
  wire w1688;
  wire w1689;
  wire w1690;
  wire w1691;
  wire w1692;
  wire w1693;
  wire w1694;
  wire w1695;
  wire w1696;
  wire w1697;
  wire w1698;
  wire w1699;
  wire w1701;
  wire w1702;
  wire w1703;
  wire w1704;
  wire w1705;
  wire w1706;
  wire w1707;
  wire w1708;
  wire w1709;
  wire w1710;
  wire w1711;
  wire w1712;
  wire w1713;
  wire w1714;
  wire w1715;
  wire w1716;
  wire w1717;
  wire w1718;
  wire w1719;
  wire w1720;
  wire w1721;
  wire w1722;
  wire w1723;
  wire w1724;
  wire w1725;
  wire w1727;
  wire w1728;
  wire w1729;
  wire w1730;
  wire w1731;
  wire w1732;
  wire w1733;
  wire w1734;
  wire w1735;
  wire w1736;
  wire w1737;
  wire w1738;
  wire w1739;
  wire w1740;
  wire w1741;
  wire w1742;
  wire w1743;
  wire w1744;
  wire w1745;
  wire w1746;
  wire w1747;
  wire w1748;
  wire w1749;
  wire w1750;
  wire w1751;
  wire w1753;
  wire w1754;
  wire w1755;
  wire w1756;
  wire w1757;
  wire w1758;
  wire w1759;
  wire w1760;
  wire w1761;
  wire w1762;
  wire w1763;
  wire w1764;
  wire w1765;
  wire w1766;
  wire w1767;
  wire w1768;
  wire w1769;
  wire w1770;
  wire w1771;
  wire w1772;
  wire w1773;
  wire w1774;
  wire w1775;
  wire w1776;
  wire w1777;
  wire w1779;
  wire w1780;
  wire w1781;
  wire w1782;
  wire w1783;
  wire w1784;
  wire w1785;
  wire w1786;
  wire w1787;
  wire w1788;
  wire w1789;
  wire w1790;
  wire w1791;
  wire w1792;
  wire w1793;
  wire w1794;
  wire w1795;
  wire w1796;
  wire w1797;
  wire w1798;
  wire w1799;
  wire w1800;
  wire w1801;
  wire w1802;
  wire w1803;
  wire w1805;
  wire w1806;
  wire w1807;
  wire w1808;
  wire w1809;
  wire w1810;
  wire w1811;
  wire w1812;
  wire w1813;
  wire w1814;
  wire w1815;
  wire w1816;
  wire w1817;
  wire w1818;
  wire w1819;
  wire w1820;
  wire w1821;
  wire w1822;
  wire w1823;
  wire w1824;
  wire w1825;
  wire w1826;
  wire w1827;
  wire w1828;
  wire w1829;
  wire w1831;
  wire w1832;
  wire w1833;
  wire w1834;
  wire w1835;
  wire w1836;
  wire w1837;
  wire w1838;
  wire w1839;
  wire w1840;
  wire w1841;
  wire w1842;
  wire w1843;
  wire w1844;
  wire w1845;
  wire w1846;
  wire w1847;
  wire w1848;
  wire w1849;
  wire w1850;
  wire w1851;
  wire w1852;
  wire w1853;
  wire w1854;
  wire w1855;
  wire w1857;
  wire w1858;
  wire w1859;
  wire w1860;
  wire w1861;
  wire w1862;
  wire w1863;
  wire w1864;
  wire w1865;
  wire w1866;
  wire w1867;
  wire w1868;
  wire w1869;
  wire w1870;
  wire w1871;
  wire w1872;
  wire w1873;
  wire w1874;
  wire w1875;
  wire w1876;
  wire w1877;
  wire w1878;
  wire w1879;
  wire w1880;
  wire w1881;
  wire w1883;
  wire w1884;
  wire w1885;
  wire w1886;
  wire w1887;
  wire w1888;
  wire w1889;
  wire w1890;
  wire w1891;
  wire w1892;
  wire w1893;
  wire w1894;
  wire w1895;
  wire w1896;
  wire w1897;
  wire w1898;
  wire w1899;
  wire w1900;
  wire w1901;
  wire w1902;
  wire w1903;
  wire w1904;
  wire w1905;
  wire w1906;
  wire w1907;
  wire w1909;
  wire w1911;
  wire w1913;
  wire w1915;
  wire w1917;
  wire w1919;
  wire w1921;
  wire w1923;
  wire w1925;
  wire w1927;
  wire w1929;
  wire w1931;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w687);
  FullAdder U1 (w687, IN2[0], IN2[1], w688, w689);
  FullAdder U2 (w689, IN3[0], IN3[1], w690, w691);
  FullAdder U3 (w691, IN4[0], IN4[1], w692, w693);
  FullAdder U4 (w693, IN5[0], IN5[1], w694, w695);
  FullAdder U5 (w695, IN6[0], IN6[1], w696, w697);
  FullAdder U6 (w697, IN7[0], IN7[1], w698, w699);
  FullAdder U7 (w699, IN8[0], IN8[1], w700, w701);
  FullAdder U8 (w701, IN9[0], IN9[1], w702, w703);
  FullAdder U9 (w703, IN10[0], IN10[1], w704, w705);
  FullAdder U10 (w705, IN11[0], IN11[1], w706, w707);
  FullAdder U11 (w707, IN12[0], IN12[1], w708, w709);
  FullAdder U12 (w709, IN13[0], IN13[1], w710, w711);
  HalfAdder U13 (w688, IN2[2], Out1[2], w713);
  FullAdder U14 (w713, w690, IN3[2], w714, w715);
  FullAdder U15 (w715, w692, IN4[2], w716, w717);
  FullAdder U16 (w717, w694, IN5[2], w718, w719);
  FullAdder U17 (w719, w696, IN6[2], w720, w721);
  FullAdder U18 (w721, w698, IN7[2], w722, w723);
  FullAdder U19 (w723, w700, IN8[2], w724, w725);
  FullAdder U20 (w725, w702, IN9[2], w726, w727);
  FullAdder U21 (w727, w704, IN10[2], w728, w729);
  FullAdder U22 (w729, w706, IN11[2], w730, w731);
  FullAdder U23 (w731, w708, IN12[2], w732, w733);
  FullAdder U24 (w733, w710, IN13[2], w734, w735);
  FullAdder U25 (w735, w711, IN14[0], w736, w737);
  HalfAdder U26 (w714, IN3[3], Out1[3], w739);
  FullAdder U27 (w739, w716, IN4[3], w740, w741);
  FullAdder U28 (w741, w718, IN5[3], w742, w743);
  FullAdder U29 (w743, w720, IN6[3], w744, w745);
  FullAdder U30 (w745, w722, IN7[3], w746, w747);
  FullAdder U31 (w747, w724, IN8[3], w748, w749);
  FullAdder U32 (w749, w726, IN9[3], w750, w751);
  FullAdder U33 (w751, w728, IN10[3], w752, w753);
  FullAdder U34 (w753, w730, IN11[3], w754, w755);
  FullAdder U35 (w755, w732, IN12[3], w756, w757);
  FullAdder U36 (w757, w734, IN13[3], w758, w759);
  FullAdder U37 (w759, w736, IN14[1], w760, w761);
  FullAdder U38 (w761, w737, IN15[0], w762, w763);
  HalfAdder U39 (w740, IN4[4], Out1[4], w765);
  FullAdder U40 (w765, w742, IN5[4], w766, w767);
  FullAdder U41 (w767, w744, IN6[4], w768, w769);
  FullAdder U42 (w769, w746, IN7[4], w770, w771);
  FullAdder U43 (w771, w748, IN8[4], w772, w773);
  FullAdder U44 (w773, w750, IN9[4], w774, w775);
  FullAdder U45 (w775, w752, IN10[4], w776, w777);
  FullAdder U46 (w777, w754, IN11[4], w778, w779);
  FullAdder U47 (w779, w756, IN12[4], w780, w781);
  FullAdder U48 (w781, w758, IN13[4], w782, w783);
  FullAdder U49 (w783, w760, IN14[2], w784, w785);
  FullAdder U50 (w785, w762, IN15[1], w786, w787);
  FullAdder U51 (w787, w763, IN16[0], w788, w789);
  HalfAdder U52 (w766, IN5[5], Out1[5], w791);
  FullAdder U53 (w791, w768, IN6[5], w792, w793);
  FullAdder U54 (w793, w770, IN7[5], w794, w795);
  FullAdder U55 (w795, w772, IN8[5], w796, w797);
  FullAdder U56 (w797, w774, IN9[5], w798, w799);
  FullAdder U57 (w799, w776, IN10[5], w800, w801);
  FullAdder U58 (w801, w778, IN11[5], w802, w803);
  FullAdder U59 (w803, w780, IN12[5], w804, w805);
  FullAdder U60 (w805, w782, IN13[5], w806, w807);
  FullAdder U61 (w807, w784, IN14[3], w808, w809);
  FullAdder U62 (w809, w786, IN15[2], w810, w811);
  FullAdder U63 (w811, w788, IN16[1], w812, w813);
  FullAdder U64 (w813, w789, IN17[0], w814, w815);
  HalfAdder U65 (w792, IN6[6], Out1[6], w817);
  FullAdder U66 (w817, w794, IN7[6], w818, w819);
  FullAdder U67 (w819, w796, IN8[6], w820, w821);
  FullAdder U68 (w821, w798, IN9[6], w822, w823);
  FullAdder U69 (w823, w800, IN10[6], w824, w825);
  FullAdder U70 (w825, w802, IN11[6], w826, w827);
  FullAdder U71 (w827, w804, IN12[6], w828, w829);
  FullAdder U72 (w829, w806, IN13[6], w830, w831);
  FullAdder U73 (w831, w808, IN14[4], w832, w833);
  FullAdder U74 (w833, w810, IN15[3], w834, w835);
  FullAdder U75 (w835, w812, IN16[2], w836, w837);
  FullAdder U76 (w837, w814, IN17[1], w838, w839);
  FullAdder U77 (w839, w815, IN18[0], w840, w841);
  HalfAdder U78 (w818, IN7[7], Out1[7], w843);
  FullAdder U79 (w843, w820, IN8[7], w844, w845);
  FullAdder U80 (w845, w822, IN9[7], w846, w847);
  FullAdder U81 (w847, w824, IN10[7], w848, w849);
  FullAdder U82 (w849, w826, IN11[7], w850, w851);
  FullAdder U83 (w851, w828, IN12[7], w852, w853);
  FullAdder U84 (w853, w830, IN13[7], w854, w855);
  FullAdder U85 (w855, w832, IN14[5], w856, w857);
  FullAdder U86 (w857, w834, IN15[4], w858, w859);
  FullAdder U87 (w859, w836, IN16[3], w860, w861);
  FullAdder U88 (w861, w838, IN17[2], w862, w863);
  FullAdder U89 (w863, w840, IN18[1], w864, w865);
  FullAdder U90 (w865, w841, IN19[0], w866, w867);
  HalfAdder U91 (w844, IN8[8], Out1[8], w869);
  FullAdder U92 (w869, w846, IN9[8], w870, w871);
  FullAdder U93 (w871, w848, IN10[8], w872, w873);
  FullAdder U94 (w873, w850, IN11[8], w874, w875);
  FullAdder U95 (w875, w852, IN12[8], w876, w877);
  FullAdder U96 (w877, w854, IN13[8], w878, w879);
  FullAdder U97 (w879, w856, IN14[6], w880, w881);
  FullAdder U98 (w881, w858, IN15[5], w882, w883);
  FullAdder U99 (w883, w860, IN16[4], w884, w885);
  FullAdder U100 (w885, w862, IN17[3], w886, w887);
  FullAdder U101 (w887, w864, IN18[2], w888, w889);
  FullAdder U102 (w889, w866, IN19[1], w890, w891);
  FullAdder U103 (w891, w867, IN20[0], w892, w893);
  HalfAdder U104 (w870, IN9[9], Out1[9], w895);
  FullAdder U105 (w895, w872, IN10[9], w896, w897);
  FullAdder U106 (w897, w874, IN11[9], w898, w899);
  FullAdder U107 (w899, w876, IN12[9], w900, w901);
  FullAdder U108 (w901, w878, IN13[9], w902, w903);
  FullAdder U109 (w903, w880, IN14[7], w904, w905);
  FullAdder U110 (w905, w882, IN15[6], w906, w907);
  FullAdder U111 (w907, w884, IN16[5], w908, w909);
  FullAdder U112 (w909, w886, IN17[4], w910, w911);
  FullAdder U113 (w911, w888, IN18[3], w912, w913);
  FullAdder U114 (w913, w890, IN19[2], w914, w915);
  FullAdder U115 (w915, w892, IN20[1], w916, w917);
  FullAdder U116 (w917, w893, IN21[0], w918, w919);
  HalfAdder U117 (w896, IN10[10], Out1[10], w921);
  FullAdder U118 (w921, w898, IN11[10], w922, w923);
  FullAdder U119 (w923, w900, IN12[10], w924, w925);
  FullAdder U120 (w925, w902, IN13[10], w926, w927);
  FullAdder U121 (w927, w904, IN14[8], w928, w929);
  FullAdder U122 (w929, w906, IN15[7], w930, w931);
  FullAdder U123 (w931, w908, IN16[6], w932, w933);
  FullAdder U124 (w933, w910, IN17[5], w934, w935);
  FullAdder U125 (w935, w912, IN18[4], w936, w937);
  FullAdder U126 (w937, w914, IN19[3], w938, w939);
  FullAdder U127 (w939, w916, IN20[2], w940, w941);
  FullAdder U128 (w941, w918, IN21[1], w942, w943);
  FullAdder U129 (w943, w919, IN22[0], w944, w945);
  HalfAdder U130 (w922, IN11[11], Out1[11], w947);
  FullAdder U131 (w947, w924, IN12[11], w948, w949);
  FullAdder U132 (w949, w926, IN13[11], w950, w951);
  FullAdder U133 (w951, w928, IN14[9], w952, w953);
  FullAdder U134 (w953, w930, IN15[8], w954, w955);
  FullAdder U135 (w955, w932, IN16[7], w956, w957);
  FullAdder U136 (w957, w934, IN17[6], w958, w959);
  FullAdder U137 (w959, w936, IN18[5], w960, w961);
  FullAdder U138 (w961, w938, IN19[4], w962, w963);
  FullAdder U139 (w963, w940, IN20[3], w964, w965);
  FullAdder U140 (w965, w942, IN21[2], w966, w967);
  FullAdder U141 (w967, w944, IN22[1], w968, w969);
  FullAdder U142 (w969, w945, IN23[0], w970, w971);
  HalfAdder U143 (w948, IN12[12], Out1[12], w973);
  FullAdder U144 (w973, w950, IN13[12], w974, w975);
  FullAdder U145 (w975, w952, IN14[10], w976, w977);
  FullAdder U146 (w977, w954, IN15[9], w978, w979);
  FullAdder U147 (w979, w956, IN16[8], w980, w981);
  FullAdder U148 (w981, w958, IN17[7], w982, w983);
  FullAdder U149 (w983, w960, IN18[6], w984, w985);
  FullAdder U150 (w985, w962, IN19[5], w986, w987);
  FullAdder U151 (w987, w964, IN20[4], w988, w989);
  FullAdder U152 (w989, w966, IN21[3], w990, w991);
  FullAdder U153 (w991, w968, IN22[2], w992, w993);
  FullAdder U154 (w993, w970, IN23[1], w994, w995);
  FullAdder U155 (w995, w971, IN24[0], w996, w997);
  HalfAdder U156 (w974, IN13[13], Out1[13], w999);
  FullAdder U157 (w999, w976, IN14[11], w1000, w1001);
  FullAdder U158 (w1001, w978, IN15[10], w1002, w1003);
  FullAdder U159 (w1003, w980, IN16[9], w1004, w1005);
  FullAdder U160 (w1005, w982, IN17[8], w1006, w1007);
  FullAdder U161 (w1007, w984, IN18[7], w1008, w1009);
  FullAdder U162 (w1009, w986, IN19[6], w1010, w1011);
  FullAdder U163 (w1011, w988, IN20[5], w1012, w1013);
  FullAdder U164 (w1013, w990, IN21[4], w1014, w1015);
  FullAdder U165 (w1015, w992, IN22[3], w1016, w1017);
  FullAdder U166 (w1017, w994, IN23[2], w1018, w1019);
  FullAdder U167 (w1019, w996, IN24[1], w1020, w1021);
  FullAdder U168 (w1021, w997, IN25[0], w1022, w1023);
  HalfAdder U169 (w1000, IN14[12], Out1[14], w1025);
  FullAdder U170 (w1025, w1002, IN15[11], w1026, w1027);
  FullAdder U171 (w1027, w1004, IN16[10], w1028, w1029);
  FullAdder U172 (w1029, w1006, IN17[9], w1030, w1031);
  FullAdder U173 (w1031, w1008, IN18[8], w1032, w1033);
  FullAdder U174 (w1033, w1010, IN19[7], w1034, w1035);
  FullAdder U175 (w1035, w1012, IN20[6], w1036, w1037);
  FullAdder U176 (w1037, w1014, IN21[5], w1038, w1039);
  FullAdder U177 (w1039, w1016, IN22[4], w1040, w1041);
  FullAdder U178 (w1041, w1018, IN23[3], w1042, w1043);
  FullAdder U179 (w1043, w1020, IN24[2], w1044, w1045);
  FullAdder U180 (w1045, w1022, IN25[1], w1046, w1047);
  FullAdder U181 (w1047, w1023, IN26[0], w1048, w1049);
  HalfAdder U182 (w1026, IN15[12], Out1[15], w1051);
  FullAdder U183 (w1051, w1028, IN16[11], w1052, w1053);
  FullAdder U184 (w1053, w1030, IN17[10], w1054, w1055);
  FullAdder U185 (w1055, w1032, IN18[9], w1056, w1057);
  FullAdder U186 (w1057, w1034, IN19[8], w1058, w1059);
  FullAdder U187 (w1059, w1036, IN20[7], w1060, w1061);
  FullAdder U188 (w1061, w1038, IN21[6], w1062, w1063);
  FullAdder U189 (w1063, w1040, IN22[5], w1064, w1065);
  FullAdder U190 (w1065, w1042, IN23[4], w1066, w1067);
  FullAdder U191 (w1067, w1044, IN24[3], w1068, w1069);
  FullAdder U192 (w1069, w1046, IN25[2], w1070, w1071);
  FullAdder U193 (w1071, w1048, IN26[1], w1072, w1073);
  FullAdder U194 (w1073, w1049, IN27[0], w1074, w1075);
  HalfAdder U195 (w1052, IN16[12], Out1[16], w1077);
  FullAdder U196 (w1077, w1054, IN17[11], w1078, w1079);
  FullAdder U197 (w1079, w1056, IN18[10], w1080, w1081);
  FullAdder U198 (w1081, w1058, IN19[9], w1082, w1083);
  FullAdder U199 (w1083, w1060, IN20[8], w1084, w1085);
  FullAdder U200 (w1085, w1062, IN21[7], w1086, w1087);
  FullAdder U201 (w1087, w1064, IN22[6], w1088, w1089);
  FullAdder U202 (w1089, w1066, IN23[5], w1090, w1091);
  FullAdder U203 (w1091, w1068, IN24[4], w1092, w1093);
  FullAdder U204 (w1093, w1070, IN25[3], w1094, w1095);
  FullAdder U205 (w1095, w1072, IN26[2], w1096, w1097);
  FullAdder U206 (w1097, w1074, IN27[1], w1098, w1099);
  FullAdder U207 (w1099, w1075, IN28[0], w1100, w1101);
  HalfAdder U208 (w1078, IN17[12], Out1[17], w1103);
  FullAdder U209 (w1103, w1080, IN18[11], w1104, w1105);
  FullAdder U210 (w1105, w1082, IN19[10], w1106, w1107);
  FullAdder U211 (w1107, w1084, IN20[9], w1108, w1109);
  FullAdder U212 (w1109, w1086, IN21[8], w1110, w1111);
  FullAdder U213 (w1111, w1088, IN22[7], w1112, w1113);
  FullAdder U214 (w1113, w1090, IN23[6], w1114, w1115);
  FullAdder U215 (w1115, w1092, IN24[5], w1116, w1117);
  FullAdder U216 (w1117, w1094, IN25[4], w1118, w1119);
  FullAdder U217 (w1119, w1096, IN26[3], w1120, w1121);
  FullAdder U218 (w1121, w1098, IN27[2], w1122, w1123);
  FullAdder U219 (w1123, w1100, IN28[1], w1124, w1125);
  FullAdder U220 (w1125, w1101, IN29[0], w1126, w1127);
  HalfAdder U221 (w1104, IN18[12], Out1[18], w1129);
  FullAdder U222 (w1129, w1106, IN19[11], w1130, w1131);
  FullAdder U223 (w1131, w1108, IN20[10], w1132, w1133);
  FullAdder U224 (w1133, w1110, IN21[9], w1134, w1135);
  FullAdder U225 (w1135, w1112, IN22[8], w1136, w1137);
  FullAdder U226 (w1137, w1114, IN23[7], w1138, w1139);
  FullAdder U227 (w1139, w1116, IN24[6], w1140, w1141);
  FullAdder U228 (w1141, w1118, IN25[5], w1142, w1143);
  FullAdder U229 (w1143, w1120, IN26[4], w1144, w1145);
  FullAdder U230 (w1145, w1122, IN27[3], w1146, w1147);
  FullAdder U231 (w1147, w1124, IN28[2], w1148, w1149);
  FullAdder U232 (w1149, w1126, IN29[1], w1150, w1151);
  FullAdder U233 (w1151, w1127, IN30[0], w1152, w1153);
  HalfAdder U234 (w1130, IN19[12], Out1[19], w1155);
  FullAdder U235 (w1155, w1132, IN20[11], w1156, w1157);
  FullAdder U236 (w1157, w1134, IN21[10], w1158, w1159);
  FullAdder U237 (w1159, w1136, IN22[9], w1160, w1161);
  FullAdder U238 (w1161, w1138, IN23[8], w1162, w1163);
  FullAdder U239 (w1163, w1140, IN24[7], w1164, w1165);
  FullAdder U240 (w1165, w1142, IN25[6], w1166, w1167);
  FullAdder U241 (w1167, w1144, IN26[5], w1168, w1169);
  FullAdder U242 (w1169, w1146, IN27[4], w1170, w1171);
  FullAdder U243 (w1171, w1148, IN28[3], w1172, w1173);
  FullAdder U244 (w1173, w1150, IN29[2], w1174, w1175);
  FullAdder U245 (w1175, w1152, IN30[1], w1176, w1177);
  FullAdder U246 (w1177, w1153, IN31[0], w1178, w1179);
  HalfAdder U247 (w1156, IN20[12], Out1[20], w1181);
  FullAdder U248 (w1181, w1158, IN21[11], w1182, w1183);
  FullAdder U249 (w1183, w1160, IN22[10], w1184, w1185);
  FullAdder U250 (w1185, w1162, IN23[9], w1186, w1187);
  FullAdder U251 (w1187, w1164, IN24[8], w1188, w1189);
  FullAdder U252 (w1189, w1166, IN25[7], w1190, w1191);
  FullAdder U253 (w1191, w1168, IN26[6], w1192, w1193);
  FullAdder U254 (w1193, w1170, IN27[5], w1194, w1195);
  FullAdder U255 (w1195, w1172, IN28[4], w1196, w1197);
  FullAdder U256 (w1197, w1174, IN29[3], w1198, w1199);
  FullAdder U257 (w1199, w1176, IN30[2], w1200, w1201);
  FullAdder U258 (w1201, w1178, IN31[1], w1202, w1203);
  FullAdder U259 (w1203, w1179, IN32[0], w1204, w1205);
  HalfAdder U260 (w1182, IN21[12], Out1[21], w1207);
  FullAdder U261 (w1207, w1184, IN22[11], w1208, w1209);
  FullAdder U262 (w1209, w1186, IN23[10], w1210, w1211);
  FullAdder U263 (w1211, w1188, IN24[9], w1212, w1213);
  FullAdder U264 (w1213, w1190, IN25[8], w1214, w1215);
  FullAdder U265 (w1215, w1192, IN26[7], w1216, w1217);
  FullAdder U266 (w1217, w1194, IN27[6], w1218, w1219);
  FullAdder U267 (w1219, w1196, IN28[5], w1220, w1221);
  FullAdder U268 (w1221, w1198, IN29[4], w1222, w1223);
  FullAdder U269 (w1223, w1200, IN30[3], w1224, w1225);
  FullAdder U270 (w1225, w1202, IN31[2], w1226, w1227);
  FullAdder U271 (w1227, w1204, IN32[1], w1228, w1229);
  FullAdder U272 (w1229, w1205, IN33[0], w1230, w1231);
  HalfAdder U273 (w1208, IN22[12], Out1[22], w1233);
  FullAdder U274 (w1233, w1210, IN23[11], w1234, w1235);
  FullAdder U275 (w1235, w1212, IN24[10], w1236, w1237);
  FullAdder U276 (w1237, w1214, IN25[9], w1238, w1239);
  FullAdder U277 (w1239, w1216, IN26[8], w1240, w1241);
  FullAdder U278 (w1241, w1218, IN27[7], w1242, w1243);
  FullAdder U279 (w1243, w1220, IN28[6], w1244, w1245);
  FullAdder U280 (w1245, w1222, IN29[5], w1246, w1247);
  FullAdder U281 (w1247, w1224, IN30[4], w1248, w1249);
  FullAdder U282 (w1249, w1226, IN31[3], w1250, w1251);
  FullAdder U283 (w1251, w1228, IN32[2], w1252, w1253);
  FullAdder U284 (w1253, w1230, IN33[1], w1254, w1255);
  FullAdder U285 (w1255, w1231, IN34[0], w1256, w1257);
  HalfAdder U286 (w1234, IN23[12], Out1[23], w1259);
  FullAdder U287 (w1259, w1236, IN24[11], w1260, w1261);
  FullAdder U288 (w1261, w1238, IN25[10], w1262, w1263);
  FullAdder U289 (w1263, w1240, IN26[9], w1264, w1265);
  FullAdder U290 (w1265, w1242, IN27[8], w1266, w1267);
  FullAdder U291 (w1267, w1244, IN28[7], w1268, w1269);
  FullAdder U292 (w1269, w1246, IN29[6], w1270, w1271);
  FullAdder U293 (w1271, w1248, IN30[5], w1272, w1273);
  FullAdder U294 (w1273, w1250, IN31[4], w1274, w1275);
  FullAdder U295 (w1275, w1252, IN32[3], w1276, w1277);
  FullAdder U296 (w1277, w1254, IN33[2], w1278, w1279);
  FullAdder U297 (w1279, w1256, IN34[1], w1280, w1281);
  FullAdder U298 (w1281, w1257, IN35[0], w1282, w1283);
  HalfAdder U299 (w1260, IN24[12], Out1[24], w1285);
  FullAdder U300 (w1285, w1262, IN25[11], w1286, w1287);
  FullAdder U301 (w1287, w1264, IN26[10], w1288, w1289);
  FullAdder U302 (w1289, w1266, IN27[9], w1290, w1291);
  FullAdder U303 (w1291, w1268, IN28[8], w1292, w1293);
  FullAdder U304 (w1293, w1270, IN29[7], w1294, w1295);
  FullAdder U305 (w1295, w1272, IN30[6], w1296, w1297);
  FullAdder U306 (w1297, w1274, IN31[5], w1298, w1299);
  FullAdder U307 (w1299, w1276, IN32[4], w1300, w1301);
  FullAdder U308 (w1301, w1278, IN33[3], w1302, w1303);
  FullAdder U309 (w1303, w1280, IN34[2], w1304, w1305);
  FullAdder U310 (w1305, w1282, IN35[1], w1306, w1307);
  FullAdder U311 (w1307, w1283, IN36[0], w1308, w1309);
  HalfAdder U312 (w1286, IN25[12], Out1[25], w1311);
  FullAdder U313 (w1311, w1288, IN26[11], w1312, w1313);
  FullAdder U314 (w1313, w1290, IN27[10], w1314, w1315);
  FullAdder U315 (w1315, w1292, IN28[9], w1316, w1317);
  FullAdder U316 (w1317, w1294, IN29[8], w1318, w1319);
  FullAdder U317 (w1319, w1296, IN30[7], w1320, w1321);
  FullAdder U318 (w1321, w1298, IN31[6], w1322, w1323);
  FullAdder U319 (w1323, w1300, IN32[5], w1324, w1325);
  FullAdder U320 (w1325, w1302, IN33[4], w1326, w1327);
  FullAdder U321 (w1327, w1304, IN34[3], w1328, w1329);
  FullAdder U322 (w1329, w1306, IN35[2], w1330, w1331);
  FullAdder U323 (w1331, w1308, IN36[1], w1332, w1333);
  FullAdder U324 (w1333, w1309, IN37[0], w1334, w1335);
  HalfAdder U325 (w1312, IN26[12], Out1[26], w1337);
  FullAdder U326 (w1337, w1314, IN27[11], w1338, w1339);
  FullAdder U327 (w1339, w1316, IN28[10], w1340, w1341);
  FullAdder U328 (w1341, w1318, IN29[9], w1342, w1343);
  FullAdder U329 (w1343, w1320, IN30[8], w1344, w1345);
  FullAdder U330 (w1345, w1322, IN31[7], w1346, w1347);
  FullAdder U331 (w1347, w1324, IN32[6], w1348, w1349);
  FullAdder U332 (w1349, w1326, IN33[5], w1350, w1351);
  FullAdder U333 (w1351, w1328, IN34[4], w1352, w1353);
  FullAdder U334 (w1353, w1330, IN35[3], w1354, w1355);
  FullAdder U335 (w1355, w1332, IN36[2], w1356, w1357);
  FullAdder U336 (w1357, w1334, IN37[1], w1358, w1359);
  FullAdder U337 (w1359, w1335, IN38[0], w1360, w1361);
  HalfAdder U338 (w1338, IN27[12], Out1[27], w1363);
  FullAdder U339 (w1363, w1340, IN28[11], w1364, w1365);
  FullAdder U340 (w1365, w1342, IN29[10], w1366, w1367);
  FullAdder U341 (w1367, w1344, IN30[9], w1368, w1369);
  FullAdder U342 (w1369, w1346, IN31[8], w1370, w1371);
  FullAdder U343 (w1371, w1348, IN32[7], w1372, w1373);
  FullAdder U344 (w1373, w1350, IN33[6], w1374, w1375);
  FullAdder U345 (w1375, w1352, IN34[5], w1376, w1377);
  FullAdder U346 (w1377, w1354, IN35[4], w1378, w1379);
  FullAdder U347 (w1379, w1356, IN36[3], w1380, w1381);
  FullAdder U348 (w1381, w1358, IN37[2], w1382, w1383);
  FullAdder U349 (w1383, w1360, IN38[1], w1384, w1385);
  FullAdder U350 (w1385, w1361, IN39[0], w1386, w1387);
  HalfAdder U351 (w1364, IN28[12], Out1[28], w1389);
  FullAdder U352 (w1389, w1366, IN29[11], w1390, w1391);
  FullAdder U353 (w1391, w1368, IN30[10], w1392, w1393);
  FullAdder U354 (w1393, w1370, IN31[9], w1394, w1395);
  FullAdder U355 (w1395, w1372, IN32[8], w1396, w1397);
  FullAdder U356 (w1397, w1374, IN33[7], w1398, w1399);
  FullAdder U357 (w1399, w1376, IN34[6], w1400, w1401);
  FullAdder U358 (w1401, w1378, IN35[5], w1402, w1403);
  FullAdder U359 (w1403, w1380, IN36[4], w1404, w1405);
  FullAdder U360 (w1405, w1382, IN37[3], w1406, w1407);
  FullAdder U361 (w1407, w1384, IN38[2], w1408, w1409);
  FullAdder U362 (w1409, w1386, IN39[1], w1410, w1411);
  FullAdder U363 (w1411, w1387, IN40[0], w1412, w1413);
  HalfAdder U364 (w1390, IN29[12], Out1[29], w1415);
  FullAdder U365 (w1415, w1392, IN30[11], w1416, w1417);
  FullAdder U366 (w1417, w1394, IN31[10], w1418, w1419);
  FullAdder U367 (w1419, w1396, IN32[9], w1420, w1421);
  FullAdder U368 (w1421, w1398, IN33[8], w1422, w1423);
  FullAdder U369 (w1423, w1400, IN34[7], w1424, w1425);
  FullAdder U370 (w1425, w1402, IN35[6], w1426, w1427);
  FullAdder U371 (w1427, w1404, IN36[5], w1428, w1429);
  FullAdder U372 (w1429, w1406, IN37[4], w1430, w1431);
  FullAdder U373 (w1431, w1408, IN38[3], w1432, w1433);
  FullAdder U374 (w1433, w1410, IN39[2], w1434, w1435);
  FullAdder U375 (w1435, w1412, IN40[1], w1436, w1437);
  FullAdder U376 (w1437, w1413, IN41[0], w1438, w1439);
  HalfAdder U377 (w1416, IN30[12], Out1[30], w1441);
  FullAdder U378 (w1441, w1418, IN31[11], w1442, w1443);
  FullAdder U379 (w1443, w1420, IN32[10], w1444, w1445);
  FullAdder U380 (w1445, w1422, IN33[9], w1446, w1447);
  FullAdder U381 (w1447, w1424, IN34[8], w1448, w1449);
  FullAdder U382 (w1449, w1426, IN35[7], w1450, w1451);
  FullAdder U383 (w1451, w1428, IN36[6], w1452, w1453);
  FullAdder U384 (w1453, w1430, IN37[5], w1454, w1455);
  FullAdder U385 (w1455, w1432, IN38[4], w1456, w1457);
  FullAdder U386 (w1457, w1434, IN39[3], w1458, w1459);
  FullAdder U387 (w1459, w1436, IN40[2], w1460, w1461);
  FullAdder U388 (w1461, w1438, IN41[1], w1462, w1463);
  FullAdder U389 (w1463, w1439, IN42[0], w1464, w1465);
  HalfAdder U390 (w1442, IN31[12], Out1[31], w1467);
  FullAdder U391 (w1467, w1444, IN32[11], w1468, w1469);
  FullAdder U392 (w1469, w1446, IN33[10], w1470, w1471);
  FullAdder U393 (w1471, w1448, IN34[9], w1472, w1473);
  FullAdder U394 (w1473, w1450, IN35[8], w1474, w1475);
  FullAdder U395 (w1475, w1452, IN36[7], w1476, w1477);
  FullAdder U396 (w1477, w1454, IN37[6], w1478, w1479);
  FullAdder U397 (w1479, w1456, IN38[5], w1480, w1481);
  FullAdder U398 (w1481, w1458, IN39[4], w1482, w1483);
  FullAdder U399 (w1483, w1460, IN40[3], w1484, w1485);
  FullAdder U400 (w1485, w1462, IN41[2], w1486, w1487);
  FullAdder U401 (w1487, w1464, IN42[1], w1488, w1489);
  FullAdder U402 (w1489, w1465, IN43[0], w1490, w1491);
  HalfAdder U403 (w1468, IN32[12], Out1[32], w1493);
  FullAdder U404 (w1493, w1470, IN33[11], w1494, w1495);
  FullAdder U405 (w1495, w1472, IN34[10], w1496, w1497);
  FullAdder U406 (w1497, w1474, IN35[9], w1498, w1499);
  FullAdder U407 (w1499, w1476, IN36[8], w1500, w1501);
  FullAdder U408 (w1501, w1478, IN37[7], w1502, w1503);
  FullAdder U409 (w1503, w1480, IN38[6], w1504, w1505);
  FullAdder U410 (w1505, w1482, IN39[5], w1506, w1507);
  FullAdder U411 (w1507, w1484, IN40[4], w1508, w1509);
  FullAdder U412 (w1509, w1486, IN41[3], w1510, w1511);
  FullAdder U413 (w1511, w1488, IN42[2], w1512, w1513);
  FullAdder U414 (w1513, w1490, IN43[1], w1514, w1515);
  FullAdder U415 (w1515, w1491, IN44[0], w1516, w1517);
  HalfAdder U416 (w1494, IN33[12], Out1[33], w1519);
  FullAdder U417 (w1519, w1496, IN34[11], w1520, w1521);
  FullAdder U418 (w1521, w1498, IN35[10], w1522, w1523);
  FullAdder U419 (w1523, w1500, IN36[9], w1524, w1525);
  FullAdder U420 (w1525, w1502, IN37[8], w1526, w1527);
  FullAdder U421 (w1527, w1504, IN38[7], w1528, w1529);
  FullAdder U422 (w1529, w1506, IN39[6], w1530, w1531);
  FullAdder U423 (w1531, w1508, IN40[5], w1532, w1533);
  FullAdder U424 (w1533, w1510, IN41[4], w1534, w1535);
  FullAdder U425 (w1535, w1512, IN42[3], w1536, w1537);
  FullAdder U426 (w1537, w1514, IN43[2], w1538, w1539);
  FullAdder U427 (w1539, w1516, IN44[1], w1540, w1541);
  FullAdder U428 (w1541, w1517, IN45[0], w1542, w1543);
  HalfAdder U429 (w1520, IN34[12], Out1[34], w1545);
  FullAdder U430 (w1545, w1522, IN35[11], w1546, w1547);
  FullAdder U431 (w1547, w1524, IN36[10], w1548, w1549);
  FullAdder U432 (w1549, w1526, IN37[9], w1550, w1551);
  FullAdder U433 (w1551, w1528, IN38[8], w1552, w1553);
  FullAdder U434 (w1553, w1530, IN39[7], w1554, w1555);
  FullAdder U435 (w1555, w1532, IN40[6], w1556, w1557);
  FullAdder U436 (w1557, w1534, IN41[5], w1558, w1559);
  FullAdder U437 (w1559, w1536, IN42[4], w1560, w1561);
  FullAdder U438 (w1561, w1538, IN43[3], w1562, w1563);
  FullAdder U439 (w1563, w1540, IN44[2], w1564, w1565);
  FullAdder U440 (w1565, w1542, IN45[1], w1566, w1567);
  FullAdder U441 (w1567, w1543, IN46[0], w1568, w1569);
  HalfAdder U442 (w1546, IN35[12], Out1[35], w1571);
  FullAdder U443 (w1571, w1548, IN36[11], w1572, w1573);
  FullAdder U444 (w1573, w1550, IN37[10], w1574, w1575);
  FullAdder U445 (w1575, w1552, IN38[9], w1576, w1577);
  FullAdder U446 (w1577, w1554, IN39[8], w1578, w1579);
  FullAdder U447 (w1579, w1556, IN40[7], w1580, w1581);
  FullAdder U448 (w1581, w1558, IN41[6], w1582, w1583);
  FullAdder U449 (w1583, w1560, IN42[5], w1584, w1585);
  FullAdder U450 (w1585, w1562, IN43[4], w1586, w1587);
  FullAdder U451 (w1587, w1564, IN44[3], w1588, w1589);
  FullAdder U452 (w1589, w1566, IN45[2], w1590, w1591);
  FullAdder U453 (w1591, w1568, IN46[1], w1592, w1593);
  FullAdder U454 (w1593, w1569, IN47[0], w1594, w1595);
  HalfAdder U455 (w1572, IN36[12], Out1[36], w1597);
  FullAdder U456 (w1597, w1574, IN37[11], w1598, w1599);
  FullAdder U457 (w1599, w1576, IN38[10], w1600, w1601);
  FullAdder U458 (w1601, w1578, IN39[9], w1602, w1603);
  FullAdder U459 (w1603, w1580, IN40[8], w1604, w1605);
  FullAdder U460 (w1605, w1582, IN41[7], w1606, w1607);
  FullAdder U461 (w1607, w1584, IN42[6], w1608, w1609);
  FullAdder U462 (w1609, w1586, IN43[5], w1610, w1611);
  FullAdder U463 (w1611, w1588, IN44[4], w1612, w1613);
  FullAdder U464 (w1613, w1590, IN45[3], w1614, w1615);
  FullAdder U465 (w1615, w1592, IN46[2], w1616, w1617);
  FullAdder U466 (w1617, w1594, IN47[1], w1618, w1619);
  FullAdder U467 (w1619, w1595, IN48[0], w1620, w1621);
  HalfAdder U468 (w1598, IN37[12], Out1[37], w1623);
  FullAdder U469 (w1623, w1600, IN38[11], w1624, w1625);
  FullAdder U470 (w1625, w1602, IN39[10], w1626, w1627);
  FullAdder U471 (w1627, w1604, IN40[9], w1628, w1629);
  FullAdder U472 (w1629, w1606, IN41[8], w1630, w1631);
  FullAdder U473 (w1631, w1608, IN42[7], w1632, w1633);
  FullAdder U474 (w1633, w1610, IN43[6], w1634, w1635);
  FullAdder U475 (w1635, w1612, IN44[5], w1636, w1637);
  FullAdder U476 (w1637, w1614, IN45[4], w1638, w1639);
  FullAdder U477 (w1639, w1616, IN46[3], w1640, w1641);
  FullAdder U478 (w1641, w1618, IN47[2], w1642, w1643);
  FullAdder U479 (w1643, w1620, IN48[1], w1644, w1645);
  FullAdder U480 (w1645, w1621, IN49[0], w1646, w1647);
  HalfAdder U481 (w1624, IN38[12], Out1[38], w1649);
  FullAdder U482 (w1649, w1626, IN39[11], w1650, w1651);
  FullAdder U483 (w1651, w1628, IN40[10], w1652, w1653);
  FullAdder U484 (w1653, w1630, IN41[9], w1654, w1655);
  FullAdder U485 (w1655, w1632, IN42[8], w1656, w1657);
  FullAdder U486 (w1657, w1634, IN43[7], w1658, w1659);
  FullAdder U487 (w1659, w1636, IN44[6], w1660, w1661);
  FullAdder U488 (w1661, w1638, IN45[5], w1662, w1663);
  FullAdder U489 (w1663, w1640, IN46[4], w1664, w1665);
  FullAdder U490 (w1665, w1642, IN47[3], w1666, w1667);
  FullAdder U491 (w1667, w1644, IN48[2], w1668, w1669);
  FullAdder U492 (w1669, w1646, IN49[1], w1670, w1671);
  FullAdder U493 (w1671, w1647, IN50[0], w1672, w1673);
  HalfAdder U494 (w1650, IN39[12], Out1[39], w1675);
  FullAdder U495 (w1675, w1652, IN40[11], w1676, w1677);
  FullAdder U496 (w1677, w1654, IN41[10], w1678, w1679);
  FullAdder U497 (w1679, w1656, IN42[9], w1680, w1681);
  FullAdder U498 (w1681, w1658, IN43[8], w1682, w1683);
  FullAdder U499 (w1683, w1660, IN44[7], w1684, w1685);
  FullAdder U500 (w1685, w1662, IN45[6], w1686, w1687);
  FullAdder U501 (w1687, w1664, IN46[5], w1688, w1689);
  FullAdder U502 (w1689, w1666, IN47[4], w1690, w1691);
  FullAdder U503 (w1691, w1668, IN48[3], w1692, w1693);
  FullAdder U504 (w1693, w1670, IN49[2], w1694, w1695);
  FullAdder U505 (w1695, w1672, IN50[1], w1696, w1697);
  FullAdder U506 (w1697, w1673, IN51[0], w1698, w1699);
  HalfAdder U507 (w1676, IN40[12], Out1[40], w1701);
  FullAdder U508 (w1701, w1678, IN41[11], w1702, w1703);
  FullAdder U509 (w1703, w1680, IN42[10], w1704, w1705);
  FullAdder U510 (w1705, w1682, IN43[9], w1706, w1707);
  FullAdder U511 (w1707, w1684, IN44[8], w1708, w1709);
  FullAdder U512 (w1709, w1686, IN45[7], w1710, w1711);
  FullAdder U513 (w1711, w1688, IN46[6], w1712, w1713);
  FullAdder U514 (w1713, w1690, IN47[5], w1714, w1715);
  FullAdder U515 (w1715, w1692, IN48[4], w1716, w1717);
  FullAdder U516 (w1717, w1694, IN49[3], w1718, w1719);
  FullAdder U517 (w1719, w1696, IN50[2], w1720, w1721);
  FullAdder U518 (w1721, w1698, IN51[1], w1722, w1723);
  FullAdder U519 (w1723, w1699, IN52[0], w1724, w1725);
  HalfAdder U520 (w1702, IN41[12], Out1[41], w1727);
  FullAdder U521 (w1727, w1704, IN42[11], w1728, w1729);
  FullAdder U522 (w1729, w1706, IN43[10], w1730, w1731);
  FullAdder U523 (w1731, w1708, IN44[9], w1732, w1733);
  FullAdder U524 (w1733, w1710, IN45[8], w1734, w1735);
  FullAdder U525 (w1735, w1712, IN46[7], w1736, w1737);
  FullAdder U526 (w1737, w1714, IN47[6], w1738, w1739);
  FullAdder U527 (w1739, w1716, IN48[5], w1740, w1741);
  FullAdder U528 (w1741, w1718, IN49[4], w1742, w1743);
  FullAdder U529 (w1743, w1720, IN50[3], w1744, w1745);
  FullAdder U530 (w1745, w1722, IN51[2], w1746, w1747);
  FullAdder U531 (w1747, w1724, IN52[1], w1748, w1749);
  FullAdder U532 (w1749, w1725, IN53[0], w1750, w1751);
  HalfAdder U533 (w1728, IN42[12], Out1[42], w1753);
  FullAdder U534 (w1753, w1730, IN43[11], w1754, w1755);
  FullAdder U535 (w1755, w1732, IN44[10], w1756, w1757);
  FullAdder U536 (w1757, w1734, IN45[9], w1758, w1759);
  FullAdder U537 (w1759, w1736, IN46[8], w1760, w1761);
  FullAdder U538 (w1761, w1738, IN47[7], w1762, w1763);
  FullAdder U539 (w1763, w1740, IN48[6], w1764, w1765);
  FullAdder U540 (w1765, w1742, IN49[5], w1766, w1767);
  FullAdder U541 (w1767, w1744, IN50[4], w1768, w1769);
  FullAdder U542 (w1769, w1746, IN51[3], w1770, w1771);
  FullAdder U543 (w1771, w1748, IN52[2], w1772, w1773);
  FullAdder U544 (w1773, w1750, IN53[1], w1774, w1775);
  FullAdder U545 (w1775, w1751, IN54[0], w1776, w1777);
  HalfAdder U546 (w1754, IN43[12], Out1[43], w1779);
  FullAdder U547 (w1779, w1756, IN44[11], w1780, w1781);
  FullAdder U548 (w1781, w1758, IN45[10], w1782, w1783);
  FullAdder U549 (w1783, w1760, IN46[9], w1784, w1785);
  FullAdder U550 (w1785, w1762, IN47[8], w1786, w1787);
  FullAdder U551 (w1787, w1764, IN48[7], w1788, w1789);
  FullAdder U552 (w1789, w1766, IN49[6], w1790, w1791);
  FullAdder U553 (w1791, w1768, IN50[5], w1792, w1793);
  FullAdder U554 (w1793, w1770, IN51[4], w1794, w1795);
  FullAdder U555 (w1795, w1772, IN52[3], w1796, w1797);
  FullAdder U556 (w1797, w1774, IN53[2], w1798, w1799);
  FullAdder U557 (w1799, w1776, IN54[1], w1800, w1801);
  FullAdder U558 (w1801, w1777, IN55[0], w1802, w1803);
  HalfAdder U559 (w1780, IN44[12], Out1[44], w1805);
  FullAdder U560 (w1805, w1782, IN45[11], w1806, w1807);
  FullAdder U561 (w1807, w1784, IN46[10], w1808, w1809);
  FullAdder U562 (w1809, w1786, IN47[9], w1810, w1811);
  FullAdder U563 (w1811, w1788, IN48[8], w1812, w1813);
  FullAdder U564 (w1813, w1790, IN49[7], w1814, w1815);
  FullAdder U565 (w1815, w1792, IN50[6], w1816, w1817);
  FullAdder U566 (w1817, w1794, IN51[5], w1818, w1819);
  FullAdder U567 (w1819, w1796, IN52[4], w1820, w1821);
  FullAdder U568 (w1821, w1798, IN53[3], w1822, w1823);
  FullAdder U569 (w1823, w1800, IN54[2], w1824, w1825);
  FullAdder U570 (w1825, w1802, IN55[1], w1826, w1827);
  FullAdder U571 (w1827, w1803, IN56[0], w1828, w1829);
  HalfAdder U572 (w1806, IN45[12], Out1[45], w1831);
  FullAdder U573 (w1831, w1808, IN46[11], w1832, w1833);
  FullAdder U574 (w1833, w1810, IN47[10], w1834, w1835);
  FullAdder U575 (w1835, w1812, IN48[9], w1836, w1837);
  FullAdder U576 (w1837, w1814, IN49[8], w1838, w1839);
  FullAdder U577 (w1839, w1816, IN50[7], w1840, w1841);
  FullAdder U578 (w1841, w1818, IN51[6], w1842, w1843);
  FullAdder U579 (w1843, w1820, IN52[5], w1844, w1845);
  FullAdder U580 (w1845, w1822, IN53[4], w1846, w1847);
  FullAdder U581 (w1847, w1824, IN54[3], w1848, w1849);
  FullAdder U582 (w1849, w1826, IN55[2], w1850, w1851);
  FullAdder U583 (w1851, w1828, IN56[1], w1852, w1853);
  FullAdder U584 (w1853, w1829, IN57[0], w1854, w1855);
  HalfAdder U585 (w1832, IN46[12], Out1[46], w1857);
  FullAdder U586 (w1857, w1834, IN47[11], w1858, w1859);
  FullAdder U587 (w1859, w1836, IN48[10], w1860, w1861);
  FullAdder U588 (w1861, w1838, IN49[9], w1862, w1863);
  FullAdder U589 (w1863, w1840, IN50[8], w1864, w1865);
  FullAdder U590 (w1865, w1842, IN51[7], w1866, w1867);
  FullAdder U591 (w1867, w1844, IN52[6], w1868, w1869);
  FullAdder U592 (w1869, w1846, IN53[5], w1870, w1871);
  FullAdder U593 (w1871, w1848, IN54[4], w1872, w1873);
  FullAdder U594 (w1873, w1850, IN55[3], w1874, w1875);
  FullAdder U595 (w1875, w1852, IN56[2], w1876, w1877);
  FullAdder U596 (w1877, w1854, IN57[1], w1878, w1879);
  FullAdder U597 (w1879, w1855, IN58[0], w1880, w1881);
  HalfAdder U598 (w1858, IN47[12], Out1[47], w1883);
  FullAdder U599 (w1883, w1860, IN48[11], w1884, w1885);
  FullAdder U600 (w1885, w1862, IN49[10], w1886, w1887);
  FullAdder U601 (w1887, w1864, IN50[9], w1888, w1889);
  FullAdder U602 (w1889, w1866, IN51[8], w1890, w1891);
  FullAdder U603 (w1891, w1868, IN52[7], w1892, w1893);
  FullAdder U604 (w1893, w1870, IN53[6], w1894, w1895);
  FullAdder U605 (w1895, w1872, IN54[5], w1896, w1897);
  FullAdder U606 (w1897, w1874, IN55[4], w1898, w1899);
  FullAdder U607 (w1899, w1876, IN56[3], w1900, w1901);
  FullAdder U608 (w1901, w1878, IN57[2], w1902, w1903);
  FullAdder U609 (w1903, w1880, IN58[1], w1904, w1905);
  FullAdder U610 (w1905, w1881, IN59[0], w1906, w1907);
  HalfAdder U611 (w1884, IN48[12], Out1[48], w1909);
  FullAdder U612 (w1909, w1886, IN49[11], Out1[49], w1911);
  FullAdder U613 (w1911, w1888, IN50[10], Out1[50], w1913);
  FullAdder U614 (w1913, w1890, IN51[9], Out1[51], w1915);
  FullAdder U615 (w1915, w1892, IN52[8], Out1[52], w1917);
  FullAdder U616 (w1917, w1894, IN53[7], Out1[53], w1919);
  FullAdder U617 (w1919, w1896, IN54[6], Out1[54], w1921);
  FullAdder U618 (w1921, w1898, IN55[5], Out1[55], w1923);
  FullAdder U619 (w1923, w1900, IN56[4], Out1[56], w1925);
  FullAdder U620 (w1925, w1902, IN57[3], Out1[57], w1927);
  FullAdder U621 (w1927, w1904, IN58[2], Out1[58], w1929);
  FullAdder U622 (w1929, w1906, IN59[1], Out1[59], w1931);
  FullAdder U623 (w1931, w1907, IN60[0], Out1[60], Out1[61]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN14[13];
  assign Out2[1] = IN15[13];
  assign Out2[2] = IN16[13];
  assign Out2[3] = IN17[13];
  assign Out2[4] = IN18[13];
  assign Out2[5] = IN19[13];
  assign Out2[6] = IN20[13];
  assign Out2[7] = IN21[13];
  assign Out2[8] = IN22[13];
  assign Out2[9] = IN23[13];
  assign Out2[10] = IN24[13];
  assign Out2[11] = IN25[13];
  assign Out2[12] = IN26[13];
  assign Out2[13] = IN27[13];
  assign Out2[14] = IN28[13];
  assign Out2[15] = IN29[13];
  assign Out2[16] = IN30[13];
  assign Out2[17] = IN31[13];
  assign Out2[18] = IN32[13];
  assign Out2[19] = IN33[13];
  assign Out2[20] = IN34[13];
  assign Out2[21] = IN35[13];
  assign Out2[22] = IN36[13];
  assign Out2[23] = IN37[13];
  assign Out2[24] = IN38[13];
  assign Out2[25] = IN39[13];
  assign Out2[26] = IN40[13];
  assign Out2[27] = IN41[13];
  assign Out2[28] = IN42[13];
  assign Out2[29] = IN43[13];
  assign Out2[30] = IN44[13];
  assign Out2[31] = IN45[13];
  assign Out2[32] = IN46[13];
  assign Out2[33] = IN47[13];
  assign Out2[34] = IN48[13];
  assign Out2[35] = IN49[12];
  assign Out2[36] = IN50[11];
  assign Out2[37] = IN51[10];
  assign Out2[38] = IN52[9];
  assign Out2[39] = IN53[8];
  assign Out2[40] = IN54[7];
  assign Out2[41] = IN55[6];
  assign Out2[42] = IN56[5];
  assign Out2[43] = IN57[4];
  assign Out2[44] = IN58[3];
  assign Out2[45] = IN59[2];
  assign Out2[46] = IN60[1];
  assign Out2[47] = IN61[0];

endmodule
module RC_48_48(IN1, IN2, Out);
  input [47:0] IN1;
  input [47:0] IN2;
  output [48:0] Out;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w97);
  FullAdder U1 (IN1[1], IN2[1], w97, Out[1], w99);
  FullAdder U2 (IN1[2], IN2[2], w99, Out[2], w101);
  FullAdder U3 (IN1[3], IN2[3], w101, Out[3], w103);
  FullAdder U4 (IN1[4], IN2[4], w103, Out[4], w105);
  FullAdder U5 (IN1[5], IN2[5], w105, Out[5], w107);
  FullAdder U6 (IN1[6], IN2[6], w107, Out[6], w109);
  FullAdder U7 (IN1[7], IN2[7], w109, Out[7], w111);
  FullAdder U8 (IN1[8], IN2[8], w111, Out[8], w113);
  FullAdder U9 (IN1[9], IN2[9], w113, Out[9], w115);
  FullAdder U10 (IN1[10], IN2[10], w115, Out[10], w117);
  FullAdder U11 (IN1[11], IN2[11], w117, Out[11], w119);
  FullAdder U12 (IN1[12], IN2[12], w119, Out[12], w121);
  FullAdder U13 (IN1[13], IN2[13], w121, Out[13], w123);
  FullAdder U14 (IN1[14], IN2[14], w123, Out[14], w125);
  FullAdder U15 (IN1[15], IN2[15], w125, Out[15], w127);
  FullAdder U16 (IN1[16], IN2[16], w127, Out[16], w129);
  FullAdder U17 (IN1[17], IN2[17], w129, Out[17], w131);
  FullAdder U18 (IN1[18], IN2[18], w131, Out[18], w133);
  FullAdder U19 (IN1[19], IN2[19], w133, Out[19], w135);
  FullAdder U20 (IN1[20], IN2[20], w135, Out[20], w137);
  FullAdder U21 (IN1[21], IN2[21], w137, Out[21], w139);
  FullAdder U22 (IN1[22], IN2[22], w139, Out[22], w141);
  FullAdder U23 (IN1[23], IN2[23], w141, Out[23], w143);
  FullAdder U24 (IN1[24], IN2[24], w143, Out[24], w145);
  FullAdder U25 (IN1[25], IN2[25], w145, Out[25], w147);
  FullAdder U26 (IN1[26], IN2[26], w147, Out[26], w149);
  FullAdder U27 (IN1[27], IN2[27], w149, Out[27], w151);
  FullAdder U28 (IN1[28], IN2[28], w151, Out[28], w153);
  FullAdder U29 (IN1[29], IN2[29], w153, Out[29], w155);
  FullAdder U30 (IN1[30], IN2[30], w155, Out[30], w157);
  FullAdder U31 (IN1[31], IN2[31], w157, Out[31], w159);
  FullAdder U32 (IN1[32], IN2[32], w159, Out[32], w161);
  FullAdder U33 (IN1[33], IN2[33], w161, Out[33], w163);
  FullAdder U34 (IN1[34], IN2[34], w163, Out[34], w165);
  FullAdder U35 (IN1[35], IN2[35], w165, Out[35], w167);
  FullAdder U36 (IN1[36], IN2[36], w167, Out[36], w169);
  FullAdder U37 (IN1[37], IN2[37], w169, Out[37], w171);
  FullAdder U38 (IN1[38], IN2[38], w171, Out[38], w173);
  FullAdder U39 (IN1[39], IN2[39], w173, Out[39], w175);
  FullAdder U40 (IN1[40], IN2[40], w175, Out[40], w177);
  FullAdder U41 (IN1[41], IN2[41], w177, Out[41], w179);
  FullAdder U42 (IN1[42], IN2[42], w179, Out[42], w181);
  FullAdder U43 (IN1[43], IN2[43], w181, Out[43], w183);
  FullAdder U44 (IN1[44], IN2[44], w183, Out[44], w185);
  FullAdder U45 (IN1[45], IN2[45], w185, Out[45], w187);
  FullAdder U46 (IN1[46], IN2[46], w187, Out[46], w189);
  FullAdder U47 (IN1[47], IN2[47], w189, Out[47], Out[48]);

endmodule
module NR_14_49(IN1, IN2, Out);
  input [13:0] IN1;
  input [48:0] IN2;
  output [62:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [13:0] P14;
  wire [13:0] P15;
  wire [13:0] P16;
  wire [13:0] P17;
  wire [13:0] P18;
  wire [13:0] P19;
  wire [13:0] P20;
  wire [13:0] P21;
  wire [13:0] P22;
  wire [13:0] P23;
  wire [13:0] P24;
  wire [13:0] P25;
  wire [13:0] P26;
  wire [13:0] P27;
  wire [13:0] P28;
  wire [13:0] P29;
  wire [13:0] P30;
  wire [13:0] P31;
  wire [13:0] P32;
  wire [13:0] P33;
  wire [13:0] P34;
  wire [13:0] P35;
  wire [13:0] P36;
  wire [13:0] P37;
  wire [13:0] P38;
  wire [13:0] P39;
  wire [13:0] P40;
  wire [13:0] P41;
  wire [13:0] P42;
  wire [13:0] P43;
  wire [13:0] P44;
  wire [13:0] P45;
  wire [13:0] P46;
  wire [13:0] P47;
  wire [13:0] P48;
  wire [12:0] P49;
  wire [11:0] P50;
  wire [10:0] P51;
  wire [9:0] P52;
  wire [8:0] P53;
  wire [7:0] P54;
  wire [6:0] P55;
  wire [5:0] P56;
  wire [4:0] P57;
  wire [3:0] P58;
  wire [2:0] P59;
  wire [1:0] P60;
  wire [0:0] P61;
  wire [61:0] R1;
  wire [47:0] R2;
  wire [62:0] aOut;
  U_SP_14_49 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, R1, R2);
  RC_48_48 S2 (R1[61:14], R2, aOut[62:14]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign Out = aOut[62:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
