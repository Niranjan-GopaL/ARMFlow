
module NR_60_1(
    input [59:0]IN1,
    input [0:0]IN2,
    output [59:0]Out
);
    assign Out = IN2;
endmodule
