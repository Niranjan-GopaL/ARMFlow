//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 12
  second input length: 37
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_12_37(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47);
  input [11:0] IN1;
  input [36:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [11:0] P12;
  output [11:0] P13;
  output [11:0] P14;
  output [11:0] P15;
  output [11:0] P16;
  output [11:0] P17;
  output [11:0] P18;
  output [11:0] P19;
  output [11:0] P20;
  output [11:0] P21;
  output [11:0] P22;
  output [11:0] P23;
  output [11:0] P24;
  output [11:0] P25;
  output [11:0] P26;
  output [11:0] P27;
  output [11:0] P28;
  output [11:0] P29;
  output [11:0] P30;
  output [11:0] P31;
  output [11:0] P32;
  output [11:0] P33;
  output [11:0] P34;
  output [11:0] P35;
  output [11:0] P36;
  output [10:0] P37;
  output [9:0] P38;
  output [8:0] P39;
  output [7:0] P40;
  output [6:0] P41;
  output [5:0] P42;
  output [4:0] P43;
  output [3:0] P44;
  output [2:0] P45;
  output [1:0] P46;
  output [0:0] P47;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[0] = IN1[1]&IN2[36];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[1] = IN1[2]&IN2[35];
  assign P38[0] = IN1[2]&IN2[36];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[2] = IN1[3]&IN2[34];
  assign P38[1] = IN1[3]&IN2[35];
  assign P39[0] = IN1[3]&IN2[36];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[3] = IN1[4]&IN2[33];
  assign P38[2] = IN1[4]&IN2[34];
  assign P39[1] = IN1[4]&IN2[35];
  assign P40[0] = IN1[4]&IN2[36];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[4] = IN1[5]&IN2[32];
  assign P38[3] = IN1[5]&IN2[33];
  assign P39[2] = IN1[5]&IN2[34];
  assign P40[1] = IN1[5]&IN2[35];
  assign P41[0] = IN1[5]&IN2[36];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[5] = IN1[6]&IN2[31];
  assign P38[4] = IN1[6]&IN2[32];
  assign P39[3] = IN1[6]&IN2[33];
  assign P40[2] = IN1[6]&IN2[34];
  assign P41[1] = IN1[6]&IN2[35];
  assign P42[0] = IN1[6]&IN2[36];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[6] = IN1[7]&IN2[30];
  assign P38[5] = IN1[7]&IN2[31];
  assign P39[4] = IN1[7]&IN2[32];
  assign P40[3] = IN1[7]&IN2[33];
  assign P41[2] = IN1[7]&IN2[34];
  assign P42[1] = IN1[7]&IN2[35];
  assign P43[0] = IN1[7]&IN2[36];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[7] = IN1[8]&IN2[29];
  assign P38[6] = IN1[8]&IN2[30];
  assign P39[5] = IN1[8]&IN2[31];
  assign P40[4] = IN1[8]&IN2[32];
  assign P41[3] = IN1[8]&IN2[33];
  assign P42[2] = IN1[8]&IN2[34];
  assign P43[1] = IN1[8]&IN2[35];
  assign P44[0] = IN1[8]&IN2[36];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[8] = IN1[9]&IN2[28];
  assign P38[7] = IN1[9]&IN2[29];
  assign P39[6] = IN1[9]&IN2[30];
  assign P40[5] = IN1[9]&IN2[31];
  assign P41[4] = IN1[9]&IN2[32];
  assign P42[3] = IN1[9]&IN2[33];
  assign P43[2] = IN1[9]&IN2[34];
  assign P44[1] = IN1[9]&IN2[35];
  assign P45[0] = IN1[9]&IN2[36];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[9] = IN1[10]&IN2[27];
  assign P38[8] = IN1[10]&IN2[28];
  assign P39[7] = IN1[10]&IN2[29];
  assign P40[6] = IN1[10]&IN2[30];
  assign P41[5] = IN1[10]&IN2[31];
  assign P42[4] = IN1[10]&IN2[32];
  assign P43[3] = IN1[10]&IN2[33];
  assign P44[2] = IN1[10]&IN2[34];
  assign P45[1] = IN1[10]&IN2[35];
  assign P46[0] = IN1[10]&IN2[36];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[10] = IN1[11]&IN2[26];
  assign P38[9] = IN1[11]&IN2[27];
  assign P39[8] = IN1[11]&IN2[28];
  assign P40[7] = IN1[11]&IN2[29];
  assign P41[6] = IN1[11]&IN2[30];
  assign P42[5] = IN1[11]&IN2[31];
  assign P43[4] = IN1[11]&IN2[32];
  assign P44[3] = IN1[11]&IN2[33];
  assign P45[2] = IN1[11]&IN2[34];
  assign P46[1] = IN1[11]&IN2[35];
  assign P47[0] = IN1[11]&IN2[36];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [11:0] IN12;
  input [11:0] IN13;
  input [11:0] IN14;
  input [11:0] IN15;
  input [11:0] IN16;
  input [11:0] IN17;
  input [11:0] IN18;
  input [11:0] IN19;
  input [11:0] IN20;
  input [11:0] IN21;
  input [11:0] IN22;
  input [11:0] IN23;
  input [11:0] IN24;
  input [11:0] IN25;
  input [11:0] IN26;
  input [11:0] IN27;
  input [11:0] IN28;
  input [11:0] IN29;
  input [11:0] IN30;
  input [11:0] IN31;
  input [11:0] IN32;
  input [11:0] IN33;
  input [11:0] IN34;
  input [11:0] IN35;
  input [11:0] IN36;
  input [10:0] IN37;
  input [9:0] IN38;
  input [8:0] IN39;
  input [7:0] IN40;
  input [6:0] IN41;
  input [5:0] IN42;
  input [4:0] IN43;
  input [3:0] IN44;
  input [2:0] IN45;
  input [1:0] IN46;
  input [0:0] IN47;
  output [47:0] Out1;
  output [35:0] Out2;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1005;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1029;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1053;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1077;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1101;
  wire w1102;
  wire w1103;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1125;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1149;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1171;
  wire w1172;
  wire w1173;
  wire w1174;
  wire w1175;
  wire w1176;
  wire w1177;
  wire w1178;
  wire w1179;
  wire w1180;
  wire w1181;
  wire w1182;
  wire w1183;
  wire w1184;
  wire w1185;
  wire w1186;
  wire w1187;
  wire w1188;
  wire w1189;
  wire w1190;
  wire w1191;
  wire w1193;
  wire w1194;
  wire w1195;
  wire w1196;
  wire w1197;
  wire w1198;
  wire w1199;
  wire w1200;
  wire w1201;
  wire w1202;
  wire w1203;
  wire w1204;
  wire w1205;
  wire w1206;
  wire w1207;
  wire w1208;
  wire w1209;
  wire w1210;
  wire w1211;
  wire w1212;
  wire w1213;
  wire w1215;
  wire w1217;
  wire w1219;
  wire w1221;
  wire w1223;
  wire w1225;
  wire w1227;
  wire w1229;
  wire w1231;
  wire w1233;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w445);
  FullAdder U1 (w445, IN2[0], IN2[1], w446, w447);
  FullAdder U2 (w447, IN3[0], IN3[1], w448, w449);
  FullAdder U3 (w449, IN4[0], IN4[1], w450, w451);
  FullAdder U4 (w451, IN5[0], IN5[1], w452, w453);
  FullAdder U5 (w453, IN6[0], IN6[1], w454, w455);
  FullAdder U6 (w455, IN7[0], IN7[1], w456, w457);
  FullAdder U7 (w457, IN8[0], IN8[1], w458, w459);
  FullAdder U8 (w459, IN9[0], IN9[1], w460, w461);
  FullAdder U9 (w461, IN10[0], IN10[1], w462, w463);
  FullAdder U10 (w463, IN11[0], IN11[1], w464, w465);
  HalfAdder U11 (w446, IN2[2], Out1[2], w467);
  FullAdder U12 (w467, w448, IN3[2], w468, w469);
  FullAdder U13 (w469, w450, IN4[2], w470, w471);
  FullAdder U14 (w471, w452, IN5[2], w472, w473);
  FullAdder U15 (w473, w454, IN6[2], w474, w475);
  FullAdder U16 (w475, w456, IN7[2], w476, w477);
  FullAdder U17 (w477, w458, IN8[2], w478, w479);
  FullAdder U18 (w479, w460, IN9[2], w480, w481);
  FullAdder U19 (w481, w462, IN10[2], w482, w483);
  FullAdder U20 (w483, w464, IN11[2], w484, w485);
  FullAdder U21 (w485, w465, IN12[0], w486, w487);
  HalfAdder U22 (w468, IN3[3], Out1[3], w489);
  FullAdder U23 (w489, w470, IN4[3], w490, w491);
  FullAdder U24 (w491, w472, IN5[3], w492, w493);
  FullAdder U25 (w493, w474, IN6[3], w494, w495);
  FullAdder U26 (w495, w476, IN7[3], w496, w497);
  FullAdder U27 (w497, w478, IN8[3], w498, w499);
  FullAdder U28 (w499, w480, IN9[3], w500, w501);
  FullAdder U29 (w501, w482, IN10[3], w502, w503);
  FullAdder U30 (w503, w484, IN11[3], w504, w505);
  FullAdder U31 (w505, w486, IN12[1], w506, w507);
  FullAdder U32 (w507, w487, IN13[0], w508, w509);
  HalfAdder U33 (w490, IN4[4], Out1[4], w511);
  FullAdder U34 (w511, w492, IN5[4], w512, w513);
  FullAdder U35 (w513, w494, IN6[4], w514, w515);
  FullAdder U36 (w515, w496, IN7[4], w516, w517);
  FullAdder U37 (w517, w498, IN8[4], w518, w519);
  FullAdder U38 (w519, w500, IN9[4], w520, w521);
  FullAdder U39 (w521, w502, IN10[4], w522, w523);
  FullAdder U40 (w523, w504, IN11[4], w524, w525);
  FullAdder U41 (w525, w506, IN12[2], w526, w527);
  FullAdder U42 (w527, w508, IN13[1], w528, w529);
  FullAdder U43 (w529, w509, IN14[0], w530, w531);
  HalfAdder U44 (w512, IN5[5], Out1[5], w533);
  FullAdder U45 (w533, w514, IN6[5], w534, w535);
  FullAdder U46 (w535, w516, IN7[5], w536, w537);
  FullAdder U47 (w537, w518, IN8[5], w538, w539);
  FullAdder U48 (w539, w520, IN9[5], w540, w541);
  FullAdder U49 (w541, w522, IN10[5], w542, w543);
  FullAdder U50 (w543, w524, IN11[5], w544, w545);
  FullAdder U51 (w545, w526, IN12[3], w546, w547);
  FullAdder U52 (w547, w528, IN13[2], w548, w549);
  FullAdder U53 (w549, w530, IN14[1], w550, w551);
  FullAdder U54 (w551, w531, IN15[0], w552, w553);
  HalfAdder U55 (w534, IN6[6], Out1[6], w555);
  FullAdder U56 (w555, w536, IN7[6], w556, w557);
  FullAdder U57 (w557, w538, IN8[6], w558, w559);
  FullAdder U58 (w559, w540, IN9[6], w560, w561);
  FullAdder U59 (w561, w542, IN10[6], w562, w563);
  FullAdder U60 (w563, w544, IN11[6], w564, w565);
  FullAdder U61 (w565, w546, IN12[4], w566, w567);
  FullAdder U62 (w567, w548, IN13[3], w568, w569);
  FullAdder U63 (w569, w550, IN14[2], w570, w571);
  FullAdder U64 (w571, w552, IN15[1], w572, w573);
  FullAdder U65 (w573, w553, IN16[0], w574, w575);
  HalfAdder U66 (w556, IN7[7], Out1[7], w577);
  FullAdder U67 (w577, w558, IN8[7], w578, w579);
  FullAdder U68 (w579, w560, IN9[7], w580, w581);
  FullAdder U69 (w581, w562, IN10[7], w582, w583);
  FullAdder U70 (w583, w564, IN11[7], w584, w585);
  FullAdder U71 (w585, w566, IN12[5], w586, w587);
  FullAdder U72 (w587, w568, IN13[4], w588, w589);
  FullAdder U73 (w589, w570, IN14[3], w590, w591);
  FullAdder U74 (w591, w572, IN15[2], w592, w593);
  FullAdder U75 (w593, w574, IN16[1], w594, w595);
  FullAdder U76 (w595, w575, IN17[0], w596, w597);
  HalfAdder U77 (w578, IN8[8], Out1[8], w599);
  FullAdder U78 (w599, w580, IN9[8], w600, w601);
  FullAdder U79 (w601, w582, IN10[8], w602, w603);
  FullAdder U80 (w603, w584, IN11[8], w604, w605);
  FullAdder U81 (w605, w586, IN12[6], w606, w607);
  FullAdder U82 (w607, w588, IN13[5], w608, w609);
  FullAdder U83 (w609, w590, IN14[4], w610, w611);
  FullAdder U84 (w611, w592, IN15[3], w612, w613);
  FullAdder U85 (w613, w594, IN16[2], w614, w615);
  FullAdder U86 (w615, w596, IN17[1], w616, w617);
  FullAdder U87 (w617, w597, IN18[0], w618, w619);
  HalfAdder U88 (w600, IN9[9], Out1[9], w621);
  FullAdder U89 (w621, w602, IN10[9], w622, w623);
  FullAdder U90 (w623, w604, IN11[9], w624, w625);
  FullAdder U91 (w625, w606, IN12[7], w626, w627);
  FullAdder U92 (w627, w608, IN13[6], w628, w629);
  FullAdder U93 (w629, w610, IN14[5], w630, w631);
  FullAdder U94 (w631, w612, IN15[4], w632, w633);
  FullAdder U95 (w633, w614, IN16[3], w634, w635);
  FullAdder U96 (w635, w616, IN17[2], w636, w637);
  FullAdder U97 (w637, w618, IN18[1], w638, w639);
  FullAdder U98 (w639, w619, IN19[0], w640, w641);
  HalfAdder U99 (w622, IN10[10], Out1[10], w643);
  FullAdder U100 (w643, w624, IN11[10], w644, w645);
  FullAdder U101 (w645, w626, IN12[8], w646, w647);
  FullAdder U102 (w647, w628, IN13[7], w648, w649);
  FullAdder U103 (w649, w630, IN14[6], w650, w651);
  FullAdder U104 (w651, w632, IN15[5], w652, w653);
  FullAdder U105 (w653, w634, IN16[4], w654, w655);
  FullAdder U106 (w655, w636, IN17[3], w656, w657);
  FullAdder U107 (w657, w638, IN18[2], w658, w659);
  FullAdder U108 (w659, w640, IN19[1], w660, w661);
  FullAdder U109 (w661, w641, IN20[0], w662, w663);
  HalfAdder U110 (w644, IN11[11], Out1[11], w665);
  FullAdder U111 (w665, w646, IN12[9], w666, w667);
  FullAdder U112 (w667, w648, IN13[8], w668, w669);
  FullAdder U113 (w669, w650, IN14[7], w670, w671);
  FullAdder U114 (w671, w652, IN15[6], w672, w673);
  FullAdder U115 (w673, w654, IN16[5], w674, w675);
  FullAdder U116 (w675, w656, IN17[4], w676, w677);
  FullAdder U117 (w677, w658, IN18[3], w678, w679);
  FullAdder U118 (w679, w660, IN19[2], w680, w681);
  FullAdder U119 (w681, w662, IN20[1], w682, w683);
  FullAdder U120 (w683, w663, IN21[0], w684, w685);
  HalfAdder U121 (w666, IN12[10], Out1[12], w687);
  FullAdder U122 (w687, w668, IN13[9], w688, w689);
  FullAdder U123 (w689, w670, IN14[8], w690, w691);
  FullAdder U124 (w691, w672, IN15[7], w692, w693);
  FullAdder U125 (w693, w674, IN16[6], w694, w695);
  FullAdder U126 (w695, w676, IN17[5], w696, w697);
  FullAdder U127 (w697, w678, IN18[4], w698, w699);
  FullAdder U128 (w699, w680, IN19[3], w700, w701);
  FullAdder U129 (w701, w682, IN20[2], w702, w703);
  FullAdder U130 (w703, w684, IN21[1], w704, w705);
  FullAdder U131 (w705, w685, IN22[0], w706, w707);
  HalfAdder U132 (w688, IN13[10], Out1[13], w709);
  FullAdder U133 (w709, w690, IN14[9], w710, w711);
  FullAdder U134 (w711, w692, IN15[8], w712, w713);
  FullAdder U135 (w713, w694, IN16[7], w714, w715);
  FullAdder U136 (w715, w696, IN17[6], w716, w717);
  FullAdder U137 (w717, w698, IN18[5], w718, w719);
  FullAdder U138 (w719, w700, IN19[4], w720, w721);
  FullAdder U139 (w721, w702, IN20[3], w722, w723);
  FullAdder U140 (w723, w704, IN21[2], w724, w725);
  FullAdder U141 (w725, w706, IN22[1], w726, w727);
  FullAdder U142 (w727, w707, IN23[0], w728, w729);
  HalfAdder U143 (w710, IN14[10], Out1[14], w731);
  FullAdder U144 (w731, w712, IN15[9], w732, w733);
  FullAdder U145 (w733, w714, IN16[8], w734, w735);
  FullAdder U146 (w735, w716, IN17[7], w736, w737);
  FullAdder U147 (w737, w718, IN18[6], w738, w739);
  FullAdder U148 (w739, w720, IN19[5], w740, w741);
  FullAdder U149 (w741, w722, IN20[4], w742, w743);
  FullAdder U150 (w743, w724, IN21[3], w744, w745);
  FullAdder U151 (w745, w726, IN22[2], w746, w747);
  FullAdder U152 (w747, w728, IN23[1], w748, w749);
  FullAdder U153 (w749, w729, IN24[0], w750, w751);
  HalfAdder U154 (w732, IN15[10], Out1[15], w753);
  FullAdder U155 (w753, w734, IN16[9], w754, w755);
  FullAdder U156 (w755, w736, IN17[8], w756, w757);
  FullAdder U157 (w757, w738, IN18[7], w758, w759);
  FullAdder U158 (w759, w740, IN19[6], w760, w761);
  FullAdder U159 (w761, w742, IN20[5], w762, w763);
  FullAdder U160 (w763, w744, IN21[4], w764, w765);
  FullAdder U161 (w765, w746, IN22[3], w766, w767);
  FullAdder U162 (w767, w748, IN23[2], w768, w769);
  FullAdder U163 (w769, w750, IN24[1], w770, w771);
  FullAdder U164 (w771, w751, IN25[0], w772, w773);
  HalfAdder U165 (w754, IN16[10], Out1[16], w775);
  FullAdder U166 (w775, w756, IN17[9], w776, w777);
  FullAdder U167 (w777, w758, IN18[8], w778, w779);
  FullAdder U168 (w779, w760, IN19[7], w780, w781);
  FullAdder U169 (w781, w762, IN20[6], w782, w783);
  FullAdder U170 (w783, w764, IN21[5], w784, w785);
  FullAdder U171 (w785, w766, IN22[4], w786, w787);
  FullAdder U172 (w787, w768, IN23[3], w788, w789);
  FullAdder U173 (w789, w770, IN24[2], w790, w791);
  FullAdder U174 (w791, w772, IN25[1], w792, w793);
  FullAdder U175 (w793, w773, IN26[0], w794, w795);
  HalfAdder U176 (w776, IN17[10], Out1[17], w797);
  FullAdder U177 (w797, w778, IN18[9], w798, w799);
  FullAdder U178 (w799, w780, IN19[8], w800, w801);
  FullAdder U179 (w801, w782, IN20[7], w802, w803);
  FullAdder U180 (w803, w784, IN21[6], w804, w805);
  FullAdder U181 (w805, w786, IN22[5], w806, w807);
  FullAdder U182 (w807, w788, IN23[4], w808, w809);
  FullAdder U183 (w809, w790, IN24[3], w810, w811);
  FullAdder U184 (w811, w792, IN25[2], w812, w813);
  FullAdder U185 (w813, w794, IN26[1], w814, w815);
  FullAdder U186 (w815, w795, IN27[0], w816, w817);
  HalfAdder U187 (w798, IN18[10], Out1[18], w819);
  FullAdder U188 (w819, w800, IN19[9], w820, w821);
  FullAdder U189 (w821, w802, IN20[8], w822, w823);
  FullAdder U190 (w823, w804, IN21[7], w824, w825);
  FullAdder U191 (w825, w806, IN22[6], w826, w827);
  FullAdder U192 (w827, w808, IN23[5], w828, w829);
  FullAdder U193 (w829, w810, IN24[4], w830, w831);
  FullAdder U194 (w831, w812, IN25[3], w832, w833);
  FullAdder U195 (w833, w814, IN26[2], w834, w835);
  FullAdder U196 (w835, w816, IN27[1], w836, w837);
  FullAdder U197 (w837, w817, IN28[0], w838, w839);
  HalfAdder U198 (w820, IN19[10], Out1[19], w841);
  FullAdder U199 (w841, w822, IN20[9], w842, w843);
  FullAdder U200 (w843, w824, IN21[8], w844, w845);
  FullAdder U201 (w845, w826, IN22[7], w846, w847);
  FullAdder U202 (w847, w828, IN23[6], w848, w849);
  FullAdder U203 (w849, w830, IN24[5], w850, w851);
  FullAdder U204 (w851, w832, IN25[4], w852, w853);
  FullAdder U205 (w853, w834, IN26[3], w854, w855);
  FullAdder U206 (w855, w836, IN27[2], w856, w857);
  FullAdder U207 (w857, w838, IN28[1], w858, w859);
  FullAdder U208 (w859, w839, IN29[0], w860, w861);
  HalfAdder U209 (w842, IN20[10], Out1[20], w863);
  FullAdder U210 (w863, w844, IN21[9], w864, w865);
  FullAdder U211 (w865, w846, IN22[8], w866, w867);
  FullAdder U212 (w867, w848, IN23[7], w868, w869);
  FullAdder U213 (w869, w850, IN24[6], w870, w871);
  FullAdder U214 (w871, w852, IN25[5], w872, w873);
  FullAdder U215 (w873, w854, IN26[4], w874, w875);
  FullAdder U216 (w875, w856, IN27[3], w876, w877);
  FullAdder U217 (w877, w858, IN28[2], w878, w879);
  FullAdder U218 (w879, w860, IN29[1], w880, w881);
  FullAdder U219 (w881, w861, IN30[0], w882, w883);
  HalfAdder U220 (w864, IN21[10], Out1[21], w885);
  FullAdder U221 (w885, w866, IN22[9], w886, w887);
  FullAdder U222 (w887, w868, IN23[8], w888, w889);
  FullAdder U223 (w889, w870, IN24[7], w890, w891);
  FullAdder U224 (w891, w872, IN25[6], w892, w893);
  FullAdder U225 (w893, w874, IN26[5], w894, w895);
  FullAdder U226 (w895, w876, IN27[4], w896, w897);
  FullAdder U227 (w897, w878, IN28[3], w898, w899);
  FullAdder U228 (w899, w880, IN29[2], w900, w901);
  FullAdder U229 (w901, w882, IN30[1], w902, w903);
  FullAdder U230 (w903, w883, IN31[0], w904, w905);
  HalfAdder U231 (w886, IN22[10], Out1[22], w907);
  FullAdder U232 (w907, w888, IN23[9], w908, w909);
  FullAdder U233 (w909, w890, IN24[8], w910, w911);
  FullAdder U234 (w911, w892, IN25[7], w912, w913);
  FullAdder U235 (w913, w894, IN26[6], w914, w915);
  FullAdder U236 (w915, w896, IN27[5], w916, w917);
  FullAdder U237 (w917, w898, IN28[4], w918, w919);
  FullAdder U238 (w919, w900, IN29[3], w920, w921);
  FullAdder U239 (w921, w902, IN30[2], w922, w923);
  FullAdder U240 (w923, w904, IN31[1], w924, w925);
  FullAdder U241 (w925, w905, IN32[0], w926, w927);
  HalfAdder U242 (w908, IN23[10], Out1[23], w929);
  FullAdder U243 (w929, w910, IN24[9], w930, w931);
  FullAdder U244 (w931, w912, IN25[8], w932, w933);
  FullAdder U245 (w933, w914, IN26[7], w934, w935);
  FullAdder U246 (w935, w916, IN27[6], w936, w937);
  FullAdder U247 (w937, w918, IN28[5], w938, w939);
  FullAdder U248 (w939, w920, IN29[4], w940, w941);
  FullAdder U249 (w941, w922, IN30[3], w942, w943);
  FullAdder U250 (w943, w924, IN31[2], w944, w945);
  FullAdder U251 (w945, w926, IN32[1], w946, w947);
  FullAdder U252 (w947, w927, IN33[0], w948, w949);
  HalfAdder U253 (w930, IN24[10], Out1[24], w951);
  FullAdder U254 (w951, w932, IN25[9], w952, w953);
  FullAdder U255 (w953, w934, IN26[8], w954, w955);
  FullAdder U256 (w955, w936, IN27[7], w956, w957);
  FullAdder U257 (w957, w938, IN28[6], w958, w959);
  FullAdder U258 (w959, w940, IN29[5], w960, w961);
  FullAdder U259 (w961, w942, IN30[4], w962, w963);
  FullAdder U260 (w963, w944, IN31[3], w964, w965);
  FullAdder U261 (w965, w946, IN32[2], w966, w967);
  FullAdder U262 (w967, w948, IN33[1], w968, w969);
  FullAdder U263 (w969, w949, IN34[0], w970, w971);
  HalfAdder U264 (w952, IN25[10], Out1[25], w973);
  FullAdder U265 (w973, w954, IN26[9], w974, w975);
  FullAdder U266 (w975, w956, IN27[8], w976, w977);
  FullAdder U267 (w977, w958, IN28[7], w978, w979);
  FullAdder U268 (w979, w960, IN29[6], w980, w981);
  FullAdder U269 (w981, w962, IN30[5], w982, w983);
  FullAdder U270 (w983, w964, IN31[4], w984, w985);
  FullAdder U271 (w985, w966, IN32[3], w986, w987);
  FullAdder U272 (w987, w968, IN33[2], w988, w989);
  FullAdder U273 (w989, w970, IN34[1], w990, w991);
  FullAdder U274 (w991, w971, IN35[0], w992, w993);
  HalfAdder U275 (w974, IN26[10], Out1[26], w995);
  FullAdder U276 (w995, w976, IN27[9], w996, w997);
  FullAdder U277 (w997, w978, IN28[8], w998, w999);
  FullAdder U278 (w999, w980, IN29[7], w1000, w1001);
  FullAdder U279 (w1001, w982, IN30[6], w1002, w1003);
  FullAdder U280 (w1003, w984, IN31[5], w1004, w1005);
  FullAdder U281 (w1005, w986, IN32[4], w1006, w1007);
  FullAdder U282 (w1007, w988, IN33[3], w1008, w1009);
  FullAdder U283 (w1009, w990, IN34[2], w1010, w1011);
  FullAdder U284 (w1011, w992, IN35[1], w1012, w1013);
  FullAdder U285 (w1013, w993, IN36[0], w1014, w1015);
  HalfAdder U286 (w996, IN27[10], Out1[27], w1017);
  FullAdder U287 (w1017, w998, IN28[9], w1018, w1019);
  FullAdder U288 (w1019, w1000, IN29[8], w1020, w1021);
  FullAdder U289 (w1021, w1002, IN30[7], w1022, w1023);
  FullAdder U290 (w1023, w1004, IN31[6], w1024, w1025);
  FullAdder U291 (w1025, w1006, IN32[5], w1026, w1027);
  FullAdder U292 (w1027, w1008, IN33[4], w1028, w1029);
  FullAdder U293 (w1029, w1010, IN34[3], w1030, w1031);
  FullAdder U294 (w1031, w1012, IN35[2], w1032, w1033);
  FullAdder U295 (w1033, w1014, IN36[1], w1034, w1035);
  FullAdder U296 (w1035, w1015, IN37[0], w1036, w1037);
  HalfAdder U297 (w1018, IN28[10], Out1[28], w1039);
  FullAdder U298 (w1039, w1020, IN29[9], w1040, w1041);
  FullAdder U299 (w1041, w1022, IN30[8], w1042, w1043);
  FullAdder U300 (w1043, w1024, IN31[7], w1044, w1045);
  FullAdder U301 (w1045, w1026, IN32[6], w1046, w1047);
  FullAdder U302 (w1047, w1028, IN33[5], w1048, w1049);
  FullAdder U303 (w1049, w1030, IN34[4], w1050, w1051);
  FullAdder U304 (w1051, w1032, IN35[3], w1052, w1053);
  FullAdder U305 (w1053, w1034, IN36[2], w1054, w1055);
  FullAdder U306 (w1055, w1036, IN37[1], w1056, w1057);
  FullAdder U307 (w1057, w1037, IN38[0], w1058, w1059);
  HalfAdder U308 (w1040, IN29[10], Out1[29], w1061);
  FullAdder U309 (w1061, w1042, IN30[9], w1062, w1063);
  FullAdder U310 (w1063, w1044, IN31[8], w1064, w1065);
  FullAdder U311 (w1065, w1046, IN32[7], w1066, w1067);
  FullAdder U312 (w1067, w1048, IN33[6], w1068, w1069);
  FullAdder U313 (w1069, w1050, IN34[5], w1070, w1071);
  FullAdder U314 (w1071, w1052, IN35[4], w1072, w1073);
  FullAdder U315 (w1073, w1054, IN36[3], w1074, w1075);
  FullAdder U316 (w1075, w1056, IN37[2], w1076, w1077);
  FullAdder U317 (w1077, w1058, IN38[1], w1078, w1079);
  FullAdder U318 (w1079, w1059, IN39[0], w1080, w1081);
  HalfAdder U319 (w1062, IN30[10], Out1[30], w1083);
  FullAdder U320 (w1083, w1064, IN31[9], w1084, w1085);
  FullAdder U321 (w1085, w1066, IN32[8], w1086, w1087);
  FullAdder U322 (w1087, w1068, IN33[7], w1088, w1089);
  FullAdder U323 (w1089, w1070, IN34[6], w1090, w1091);
  FullAdder U324 (w1091, w1072, IN35[5], w1092, w1093);
  FullAdder U325 (w1093, w1074, IN36[4], w1094, w1095);
  FullAdder U326 (w1095, w1076, IN37[3], w1096, w1097);
  FullAdder U327 (w1097, w1078, IN38[2], w1098, w1099);
  FullAdder U328 (w1099, w1080, IN39[1], w1100, w1101);
  FullAdder U329 (w1101, w1081, IN40[0], w1102, w1103);
  HalfAdder U330 (w1084, IN31[10], Out1[31], w1105);
  FullAdder U331 (w1105, w1086, IN32[9], w1106, w1107);
  FullAdder U332 (w1107, w1088, IN33[8], w1108, w1109);
  FullAdder U333 (w1109, w1090, IN34[7], w1110, w1111);
  FullAdder U334 (w1111, w1092, IN35[6], w1112, w1113);
  FullAdder U335 (w1113, w1094, IN36[5], w1114, w1115);
  FullAdder U336 (w1115, w1096, IN37[4], w1116, w1117);
  FullAdder U337 (w1117, w1098, IN38[3], w1118, w1119);
  FullAdder U338 (w1119, w1100, IN39[2], w1120, w1121);
  FullAdder U339 (w1121, w1102, IN40[1], w1122, w1123);
  FullAdder U340 (w1123, w1103, IN41[0], w1124, w1125);
  HalfAdder U341 (w1106, IN32[10], Out1[32], w1127);
  FullAdder U342 (w1127, w1108, IN33[9], w1128, w1129);
  FullAdder U343 (w1129, w1110, IN34[8], w1130, w1131);
  FullAdder U344 (w1131, w1112, IN35[7], w1132, w1133);
  FullAdder U345 (w1133, w1114, IN36[6], w1134, w1135);
  FullAdder U346 (w1135, w1116, IN37[5], w1136, w1137);
  FullAdder U347 (w1137, w1118, IN38[4], w1138, w1139);
  FullAdder U348 (w1139, w1120, IN39[3], w1140, w1141);
  FullAdder U349 (w1141, w1122, IN40[2], w1142, w1143);
  FullAdder U350 (w1143, w1124, IN41[1], w1144, w1145);
  FullAdder U351 (w1145, w1125, IN42[0], w1146, w1147);
  HalfAdder U352 (w1128, IN33[10], Out1[33], w1149);
  FullAdder U353 (w1149, w1130, IN34[9], w1150, w1151);
  FullAdder U354 (w1151, w1132, IN35[8], w1152, w1153);
  FullAdder U355 (w1153, w1134, IN36[7], w1154, w1155);
  FullAdder U356 (w1155, w1136, IN37[6], w1156, w1157);
  FullAdder U357 (w1157, w1138, IN38[5], w1158, w1159);
  FullAdder U358 (w1159, w1140, IN39[4], w1160, w1161);
  FullAdder U359 (w1161, w1142, IN40[3], w1162, w1163);
  FullAdder U360 (w1163, w1144, IN41[2], w1164, w1165);
  FullAdder U361 (w1165, w1146, IN42[1], w1166, w1167);
  FullAdder U362 (w1167, w1147, IN43[0], w1168, w1169);
  HalfAdder U363 (w1150, IN34[10], Out1[34], w1171);
  FullAdder U364 (w1171, w1152, IN35[9], w1172, w1173);
  FullAdder U365 (w1173, w1154, IN36[8], w1174, w1175);
  FullAdder U366 (w1175, w1156, IN37[7], w1176, w1177);
  FullAdder U367 (w1177, w1158, IN38[6], w1178, w1179);
  FullAdder U368 (w1179, w1160, IN39[5], w1180, w1181);
  FullAdder U369 (w1181, w1162, IN40[4], w1182, w1183);
  FullAdder U370 (w1183, w1164, IN41[3], w1184, w1185);
  FullAdder U371 (w1185, w1166, IN42[2], w1186, w1187);
  FullAdder U372 (w1187, w1168, IN43[1], w1188, w1189);
  FullAdder U373 (w1189, w1169, IN44[0], w1190, w1191);
  HalfAdder U374 (w1172, IN35[10], Out1[35], w1193);
  FullAdder U375 (w1193, w1174, IN36[9], w1194, w1195);
  FullAdder U376 (w1195, w1176, IN37[8], w1196, w1197);
  FullAdder U377 (w1197, w1178, IN38[7], w1198, w1199);
  FullAdder U378 (w1199, w1180, IN39[6], w1200, w1201);
  FullAdder U379 (w1201, w1182, IN40[5], w1202, w1203);
  FullAdder U380 (w1203, w1184, IN41[4], w1204, w1205);
  FullAdder U381 (w1205, w1186, IN42[3], w1206, w1207);
  FullAdder U382 (w1207, w1188, IN43[2], w1208, w1209);
  FullAdder U383 (w1209, w1190, IN44[1], w1210, w1211);
  FullAdder U384 (w1211, w1191, IN45[0], w1212, w1213);
  HalfAdder U385 (w1194, IN36[10], Out1[36], w1215);
  FullAdder U386 (w1215, w1196, IN37[9], Out1[37], w1217);
  FullAdder U387 (w1217, w1198, IN38[8], Out1[38], w1219);
  FullAdder U388 (w1219, w1200, IN39[7], Out1[39], w1221);
  FullAdder U389 (w1221, w1202, IN40[6], Out1[40], w1223);
  FullAdder U390 (w1223, w1204, IN41[5], Out1[41], w1225);
  FullAdder U391 (w1225, w1206, IN42[4], Out1[42], w1227);
  FullAdder U392 (w1227, w1208, IN43[3], Out1[43], w1229);
  FullAdder U393 (w1229, w1210, IN44[2], Out1[44], w1231);
  FullAdder U394 (w1231, w1212, IN45[1], Out1[45], w1233);
  FullAdder U395 (w1233, w1213, IN46[0], Out1[46], Out1[47]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN12[11];
  assign Out2[1] = IN13[11];
  assign Out2[2] = IN14[11];
  assign Out2[3] = IN15[11];
  assign Out2[4] = IN16[11];
  assign Out2[5] = IN17[11];
  assign Out2[6] = IN18[11];
  assign Out2[7] = IN19[11];
  assign Out2[8] = IN20[11];
  assign Out2[9] = IN21[11];
  assign Out2[10] = IN22[11];
  assign Out2[11] = IN23[11];
  assign Out2[12] = IN24[11];
  assign Out2[13] = IN25[11];
  assign Out2[14] = IN26[11];
  assign Out2[15] = IN27[11];
  assign Out2[16] = IN28[11];
  assign Out2[17] = IN29[11];
  assign Out2[18] = IN30[11];
  assign Out2[19] = IN31[11];
  assign Out2[20] = IN32[11];
  assign Out2[21] = IN33[11];
  assign Out2[22] = IN34[11];
  assign Out2[23] = IN35[11];
  assign Out2[24] = IN36[11];
  assign Out2[25] = IN37[10];
  assign Out2[26] = IN38[9];
  assign Out2[27] = IN39[8];
  assign Out2[28] = IN40[7];
  assign Out2[29] = IN41[6];
  assign Out2[30] = IN42[5];
  assign Out2[31] = IN43[4];
  assign Out2[32] = IN44[3];
  assign Out2[33] = IN45[2];
  assign Out2[34] = IN46[1];
  assign Out2[35] = IN47[0];

endmodule
module RC_36_36(IN1, IN2, Out);
  input [35:0] IN1;
  input [35:0] IN2;
  output [36:0] Out;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w73);
  FullAdder U1 (IN1[1], IN2[1], w73, Out[1], w75);
  FullAdder U2 (IN1[2], IN2[2], w75, Out[2], w77);
  FullAdder U3 (IN1[3], IN2[3], w77, Out[3], w79);
  FullAdder U4 (IN1[4], IN2[4], w79, Out[4], w81);
  FullAdder U5 (IN1[5], IN2[5], w81, Out[5], w83);
  FullAdder U6 (IN1[6], IN2[6], w83, Out[6], w85);
  FullAdder U7 (IN1[7], IN2[7], w85, Out[7], w87);
  FullAdder U8 (IN1[8], IN2[8], w87, Out[8], w89);
  FullAdder U9 (IN1[9], IN2[9], w89, Out[9], w91);
  FullAdder U10 (IN1[10], IN2[10], w91, Out[10], w93);
  FullAdder U11 (IN1[11], IN2[11], w93, Out[11], w95);
  FullAdder U12 (IN1[12], IN2[12], w95, Out[12], w97);
  FullAdder U13 (IN1[13], IN2[13], w97, Out[13], w99);
  FullAdder U14 (IN1[14], IN2[14], w99, Out[14], w101);
  FullAdder U15 (IN1[15], IN2[15], w101, Out[15], w103);
  FullAdder U16 (IN1[16], IN2[16], w103, Out[16], w105);
  FullAdder U17 (IN1[17], IN2[17], w105, Out[17], w107);
  FullAdder U18 (IN1[18], IN2[18], w107, Out[18], w109);
  FullAdder U19 (IN1[19], IN2[19], w109, Out[19], w111);
  FullAdder U20 (IN1[20], IN2[20], w111, Out[20], w113);
  FullAdder U21 (IN1[21], IN2[21], w113, Out[21], w115);
  FullAdder U22 (IN1[22], IN2[22], w115, Out[22], w117);
  FullAdder U23 (IN1[23], IN2[23], w117, Out[23], w119);
  FullAdder U24 (IN1[24], IN2[24], w119, Out[24], w121);
  FullAdder U25 (IN1[25], IN2[25], w121, Out[25], w123);
  FullAdder U26 (IN1[26], IN2[26], w123, Out[26], w125);
  FullAdder U27 (IN1[27], IN2[27], w125, Out[27], w127);
  FullAdder U28 (IN1[28], IN2[28], w127, Out[28], w129);
  FullAdder U29 (IN1[29], IN2[29], w129, Out[29], w131);
  FullAdder U30 (IN1[30], IN2[30], w131, Out[30], w133);
  FullAdder U31 (IN1[31], IN2[31], w133, Out[31], w135);
  FullAdder U32 (IN1[32], IN2[32], w135, Out[32], w137);
  FullAdder U33 (IN1[33], IN2[33], w137, Out[33], w139);
  FullAdder U34 (IN1[34], IN2[34], w139, Out[34], w141);
  FullAdder U35 (IN1[35], IN2[35], w141, Out[35], Out[36]);

endmodule
module NR_12_37(IN1, IN2, Out);
  input [11:0] IN1;
  input [36:0] IN2;
  output [48:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [11:0] P12;
  wire [11:0] P13;
  wire [11:0] P14;
  wire [11:0] P15;
  wire [11:0] P16;
  wire [11:0] P17;
  wire [11:0] P18;
  wire [11:0] P19;
  wire [11:0] P20;
  wire [11:0] P21;
  wire [11:0] P22;
  wire [11:0] P23;
  wire [11:0] P24;
  wire [11:0] P25;
  wire [11:0] P26;
  wire [11:0] P27;
  wire [11:0] P28;
  wire [11:0] P29;
  wire [11:0] P30;
  wire [11:0] P31;
  wire [11:0] P32;
  wire [11:0] P33;
  wire [11:0] P34;
  wire [11:0] P35;
  wire [11:0] P36;
  wire [10:0] P37;
  wire [9:0] P38;
  wire [8:0] P39;
  wire [7:0] P40;
  wire [6:0] P41;
  wire [5:0] P42;
  wire [4:0] P43;
  wire [3:0] P44;
  wire [2:0] P45;
  wire [1:0] P46;
  wire [0:0] P47;
  wire [47:0] R1;
  wire [35:0] R2;
  wire [48:0] aOut;
  U_SP_12_37 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, R1, R2);
  RC_36_36 S2 (R1[47:12], R2, aOut[48:12]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign Out = aOut[48:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
