//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 8
  second input length: 37
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_8_37(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43);
  input [7:0] IN1;
  input [36:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [7:0] P8;
  output [7:0] P9;
  output [7:0] P10;
  output [7:0] P11;
  output [7:0] P12;
  output [7:0] P13;
  output [7:0] P14;
  output [7:0] P15;
  output [7:0] P16;
  output [7:0] P17;
  output [7:0] P18;
  output [7:0] P19;
  output [7:0] P20;
  output [7:0] P21;
  output [7:0] P22;
  output [7:0] P23;
  output [7:0] P24;
  output [7:0] P25;
  output [7:0] P26;
  output [7:0] P27;
  output [7:0] P28;
  output [7:0] P29;
  output [7:0] P30;
  output [7:0] P31;
  output [7:0] P32;
  output [7:0] P33;
  output [7:0] P34;
  output [7:0] P35;
  output [7:0] P36;
  output [6:0] P37;
  output [5:0] P38;
  output [4:0] P39;
  output [3:0] P40;
  output [2:0] P41;
  output [1:0] P42;
  output [0:0] P43;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[0] = IN1[1]&IN2[36];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[1] = IN1[2]&IN2[35];
  assign P38[0] = IN1[2]&IN2[36];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[2] = IN1[3]&IN2[34];
  assign P38[1] = IN1[3]&IN2[35];
  assign P39[0] = IN1[3]&IN2[36];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[3] = IN1[4]&IN2[33];
  assign P38[2] = IN1[4]&IN2[34];
  assign P39[1] = IN1[4]&IN2[35];
  assign P40[0] = IN1[4]&IN2[36];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[4] = IN1[5]&IN2[32];
  assign P38[3] = IN1[5]&IN2[33];
  assign P39[2] = IN1[5]&IN2[34];
  assign P40[1] = IN1[5]&IN2[35];
  assign P41[0] = IN1[5]&IN2[36];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[5] = IN1[6]&IN2[31];
  assign P38[4] = IN1[6]&IN2[32];
  assign P39[3] = IN1[6]&IN2[33];
  assign P40[2] = IN1[6]&IN2[34];
  assign P41[1] = IN1[6]&IN2[35];
  assign P42[0] = IN1[6]&IN2[36];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[6] = IN1[7]&IN2[30];
  assign P38[5] = IN1[7]&IN2[31];
  assign P39[4] = IN1[7]&IN2[32];
  assign P40[3] = IN1[7]&IN2[33];
  assign P41[2] = IN1[7]&IN2[34];
  assign P42[1] = IN1[7]&IN2[35];
  assign P43[0] = IN1[7]&IN2[36];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [7:0] IN8;
  input [7:0] IN9;
  input [7:0] IN10;
  input [7:0] IN11;
  input [7:0] IN12;
  input [7:0] IN13;
  input [7:0] IN14;
  input [7:0] IN15;
  input [7:0] IN16;
  input [7:0] IN17;
  input [7:0] IN18;
  input [7:0] IN19;
  input [7:0] IN20;
  input [7:0] IN21;
  input [7:0] IN22;
  input [7:0] IN23;
  input [7:0] IN24;
  input [7:0] IN25;
  input [7:0] IN26;
  input [7:0] IN27;
  input [7:0] IN28;
  input [7:0] IN29;
  input [7:0] IN30;
  input [7:0] IN31;
  input [7:0] IN32;
  input [7:0] IN33;
  input [7:0] IN34;
  input [7:0] IN35;
  input [7:0] IN36;
  input [6:0] IN37;
  input [5:0] IN38;
  input [4:0] IN39;
  input [3:0] IN40;
  input [2:0] IN41;
  input [1:0] IN42;
  input [0:0] IN43;
  output [43:0] Out1;
  output [35:0] Out2;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w787;
  wire w789;
  wire w791;
  wire w793;
  wire w795;
  wire w797;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w297);
  FullAdder U1 (w297, IN2[0], IN2[1], w298, w299);
  FullAdder U2 (w299, IN3[0], IN3[1], w300, w301);
  FullAdder U3 (w301, IN4[0], IN4[1], w302, w303);
  FullAdder U4 (w303, IN5[0], IN5[1], w304, w305);
  FullAdder U5 (w305, IN6[0], IN6[1], w306, w307);
  FullAdder U6 (w307, IN7[0], IN7[1], w308, w309);
  HalfAdder U7 (w298, IN2[2], Out1[2], w311);
  FullAdder U8 (w311, w300, IN3[2], w312, w313);
  FullAdder U9 (w313, w302, IN4[2], w314, w315);
  FullAdder U10 (w315, w304, IN5[2], w316, w317);
  FullAdder U11 (w317, w306, IN6[2], w318, w319);
  FullAdder U12 (w319, w308, IN7[2], w320, w321);
  FullAdder U13 (w321, w309, IN8[0], w322, w323);
  HalfAdder U14 (w312, IN3[3], Out1[3], w325);
  FullAdder U15 (w325, w314, IN4[3], w326, w327);
  FullAdder U16 (w327, w316, IN5[3], w328, w329);
  FullAdder U17 (w329, w318, IN6[3], w330, w331);
  FullAdder U18 (w331, w320, IN7[3], w332, w333);
  FullAdder U19 (w333, w322, IN8[1], w334, w335);
  FullAdder U20 (w335, w323, IN9[0], w336, w337);
  HalfAdder U21 (w326, IN4[4], Out1[4], w339);
  FullAdder U22 (w339, w328, IN5[4], w340, w341);
  FullAdder U23 (w341, w330, IN6[4], w342, w343);
  FullAdder U24 (w343, w332, IN7[4], w344, w345);
  FullAdder U25 (w345, w334, IN8[2], w346, w347);
  FullAdder U26 (w347, w336, IN9[1], w348, w349);
  FullAdder U27 (w349, w337, IN10[0], w350, w351);
  HalfAdder U28 (w340, IN5[5], Out1[5], w353);
  FullAdder U29 (w353, w342, IN6[5], w354, w355);
  FullAdder U30 (w355, w344, IN7[5], w356, w357);
  FullAdder U31 (w357, w346, IN8[3], w358, w359);
  FullAdder U32 (w359, w348, IN9[2], w360, w361);
  FullAdder U33 (w361, w350, IN10[1], w362, w363);
  FullAdder U34 (w363, w351, IN11[0], w364, w365);
  HalfAdder U35 (w354, IN6[6], Out1[6], w367);
  FullAdder U36 (w367, w356, IN7[6], w368, w369);
  FullAdder U37 (w369, w358, IN8[4], w370, w371);
  FullAdder U38 (w371, w360, IN9[3], w372, w373);
  FullAdder U39 (w373, w362, IN10[2], w374, w375);
  FullAdder U40 (w375, w364, IN11[1], w376, w377);
  FullAdder U41 (w377, w365, IN12[0], w378, w379);
  HalfAdder U42 (w368, IN7[7], Out1[7], w381);
  FullAdder U43 (w381, w370, IN8[5], w382, w383);
  FullAdder U44 (w383, w372, IN9[4], w384, w385);
  FullAdder U45 (w385, w374, IN10[3], w386, w387);
  FullAdder U46 (w387, w376, IN11[2], w388, w389);
  FullAdder U47 (w389, w378, IN12[1], w390, w391);
  FullAdder U48 (w391, w379, IN13[0], w392, w393);
  HalfAdder U49 (w382, IN8[6], Out1[8], w395);
  FullAdder U50 (w395, w384, IN9[5], w396, w397);
  FullAdder U51 (w397, w386, IN10[4], w398, w399);
  FullAdder U52 (w399, w388, IN11[3], w400, w401);
  FullAdder U53 (w401, w390, IN12[2], w402, w403);
  FullAdder U54 (w403, w392, IN13[1], w404, w405);
  FullAdder U55 (w405, w393, IN14[0], w406, w407);
  HalfAdder U56 (w396, IN9[6], Out1[9], w409);
  FullAdder U57 (w409, w398, IN10[5], w410, w411);
  FullAdder U58 (w411, w400, IN11[4], w412, w413);
  FullAdder U59 (w413, w402, IN12[3], w414, w415);
  FullAdder U60 (w415, w404, IN13[2], w416, w417);
  FullAdder U61 (w417, w406, IN14[1], w418, w419);
  FullAdder U62 (w419, w407, IN15[0], w420, w421);
  HalfAdder U63 (w410, IN10[6], Out1[10], w423);
  FullAdder U64 (w423, w412, IN11[5], w424, w425);
  FullAdder U65 (w425, w414, IN12[4], w426, w427);
  FullAdder U66 (w427, w416, IN13[3], w428, w429);
  FullAdder U67 (w429, w418, IN14[2], w430, w431);
  FullAdder U68 (w431, w420, IN15[1], w432, w433);
  FullAdder U69 (w433, w421, IN16[0], w434, w435);
  HalfAdder U70 (w424, IN11[6], Out1[11], w437);
  FullAdder U71 (w437, w426, IN12[5], w438, w439);
  FullAdder U72 (w439, w428, IN13[4], w440, w441);
  FullAdder U73 (w441, w430, IN14[3], w442, w443);
  FullAdder U74 (w443, w432, IN15[2], w444, w445);
  FullAdder U75 (w445, w434, IN16[1], w446, w447);
  FullAdder U76 (w447, w435, IN17[0], w448, w449);
  HalfAdder U77 (w438, IN12[6], Out1[12], w451);
  FullAdder U78 (w451, w440, IN13[5], w452, w453);
  FullAdder U79 (w453, w442, IN14[4], w454, w455);
  FullAdder U80 (w455, w444, IN15[3], w456, w457);
  FullAdder U81 (w457, w446, IN16[2], w458, w459);
  FullAdder U82 (w459, w448, IN17[1], w460, w461);
  FullAdder U83 (w461, w449, IN18[0], w462, w463);
  HalfAdder U84 (w452, IN13[6], Out1[13], w465);
  FullAdder U85 (w465, w454, IN14[5], w466, w467);
  FullAdder U86 (w467, w456, IN15[4], w468, w469);
  FullAdder U87 (w469, w458, IN16[3], w470, w471);
  FullAdder U88 (w471, w460, IN17[2], w472, w473);
  FullAdder U89 (w473, w462, IN18[1], w474, w475);
  FullAdder U90 (w475, w463, IN19[0], w476, w477);
  HalfAdder U91 (w466, IN14[6], Out1[14], w479);
  FullAdder U92 (w479, w468, IN15[5], w480, w481);
  FullAdder U93 (w481, w470, IN16[4], w482, w483);
  FullAdder U94 (w483, w472, IN17[3], w484, w485);
  FullAdder U95 (w485, w474, IN18[2], w486, w487);
  FullAdder U96 (w487, w476, IN19[1], w488, w489);
  FullAdder U97 (w489, w477, IN20[0], w490, w491);
  HalfAdder U98 (w480, IN15[6], Out1[15], w493);
  FullAdder U99 (w493, w482, IN16[5], w494, w495);
  FullAdder U100 (w495, w484, IN17[4], w496, w497);
  FullAdder U101 (w497, w486, IN18[3], w498, w499);
  FullAdder U102 (w499, w488, IN19[2], w500, w501);
  FullAdder U103 (w501, w490, IN20[1], w502, w503);
  FullAdder U104 (w503, w491, IN21[0], w504, w505);
  HalfAdder U105 (w494, IN16[6], Out1[16], w507);
  FullAdder U106 (w507, w496, IN17[5], w508, w509);
  FullAdder U107 (w509, w498, IN18[4], w510, w511);
  FullAdder U108 (w511, w500, IN19[3], w512, w513);
  FullAdder U109 (w513, w502, IN20[2], w514, w515);
  FullAdder U110 (w515, w504, IN21[1], w516, w517);
  FullAdder U111 (w517, w505, IN22[0], w518, w519);
  HalfAdder U112 (w508, IN17[6], Out1[17], w521);
  FullAdder U113 (w521, w510, IN18[5], w522, w523);
  FullAdder U114 (w523, w512, IN19[4], w524, w525);
  FullAdder U115 (w525, w514, IN20[3], w526, w527);
  FullAdder U116 (w527, w516, IN21[2], w528, w529);
  FullAdder U117 (w529, w518, IN22[1], w530, w531);
  FullAdder U118 (w531, w519, IN23[0], w532, w533);
  HalfAdder U119 (w522, IN18[6], Out1[18], w535);
  FullAdder U120 (w535, w524, IN19[5], w536, w537);
  FullAdder U121 (w537, w526, IN20[4], w538, w539);
  FullAdder U122 (w539, w528, IN21[3], w540, w541);
  FullAdder U123 (w541, w530, IN22[2], w542, w543);
  FullAdder U124 (w543, w532, IN23[1], w544, w545);
  FullAdder U125 (w545, w533, IN24[0], w546, w547);
  HalfAdder U126 (w536, IN19[6], Out1[19], w549);
  FullAdder U127 (w549, w538, IN20[5], w550, w551);
  FullAdder U128 (w551, w540, IN21[4], w552, w553);
  FullAdder U129 (w553, w542, IN22[3], w554, w555);
  FullAdder U130 (w555, w544, IN23[2], w556, w557);
  FullAdder U131 (w557, w546, IN24[1], w558, w559);
  FullAdder U132 (w559, w547, IN25[0], w560, w561);
  HalfAdder U133 (w550, IN20[6], Out1[20], w563);
  FullAdder U134 (w563, w552, IN21[5], w564, w565);
  FullAdder U135 (w565, w554, IN22[4], w566, w567);
  FullAdder U136 (w567, w556, IN23[3], w568, w569);
  FullAdder U137 (w569, w558, IN24[2], w570, w571);
  FullAdder U138 (w571, w560, IN25[1], w572, w573);
  FullAdder U139 (w573, w561, IN26[0], w574, w575);
  HalfAdder U140 (w564, IN21[6], Out1[21], w577);
  FullAdder U141 (w577, w566, IN22[5], w578, w579);
  FullAdder U142 (w579, w568, IN23[4], w580, w581);
  FullAdder U143 (w581, w570, IN24[3], w582, w583);
  FullAdder U144 (w583, w572, IN25[2], w584, w585);
  FullAdder U145 (w585, w574, IN26[1], w586, w587);
  FullAdder U146 (w587, w575, IN27[0], w588, w589);
  HalfAdder U147 (w578, IN22[6], Out1[22], w591);
  FullAdder U148 (w591, w580, IN23[5], w592, w593);
  FullAdder U149 (w593, w582, IN24[4], w594, w595);
  FullAdder U150 (w595, w584, IN25[3], w596, w597);
  FullAdder U151 (w597, w586, IN26[2], w598, w599);
  FullAdder U152 (w599, w588, IN27[1], w600, w601);
  FullAdder U153 (w601, w589, IN28[0], w602, w603);
  HalfAdder U154 (w592, IN23[6], Out1[23], w605);
  FullAdder U155 (w605, w594, IN24[5], w606, w607);
  FullAdder U156 (w607, w596, IN25[4], w608, w609);
  FullAdder U157 (w609, w598, IN26[3], w610, w611);
  FullAdder U158 (w611, w600, IN27[2], w612, w613);
  FullAdder U159 (w613, w602, IN28[1], w614, w615);
  FullAdder U160 (w615, w603, IN29[0], w616, w617);
  HalfAdder U161 (w606, IN24[6], Out1[24], w619);
  FullAdder U162 (w619, w608, IN25[5], w620, w621);
  FullAdder U163 (w621, w610, IN26[4], w622, w623);
  FullAdder U164 (w623, w612, IN27[3], w624, w625);
  FullAdder U165 (w625, w614, IN28[2], w626, w627);
  FullAdder U166 (w627, w616, IN29[1], w628, w629);
  FullAdder U167 (w629, w617, IN30[0], w630, w631);
  HalfAdder U168 (w620, IN25[6], Out1[25], w633);
  FullAdder U169 (w633, w622, IN26[5], w634, w635);
  FullAdder U170 (w635, w624, IN27[4], w636, w637);
  FullAdder U171 (w637, w626, IN28[3], w638, w639);
  FullAdder U172 (w639, w628, IN29[2], w640, w641);
  FullAdder U173 (w641, w630, IN30[1], w642, w643);
  FullAdder U174 (w643, w631, IN31[0], w644, w645);
  HalfAdder U175 (w634, IN26[6], Out1[26], w647);
  FullAdder U176 (w647, w636, IN27[5], w648, w649);
  FullAdder U177 (w649, w638, IN28[4], w650, w651);
  FullAdder U178 (w651, w640, IN29[3], w652, w653);
  FullAdder U179 (w653, w642, IN30[2], w654, w655);
  FullAdder U180 (w655, w644, IN31[1], w656, w657);
  FullAdder U181 (w657, w645, IN32[0], w658, w659);
  HalfAdder U182 (w648, IN27[6], Out1[27], w661);
  FullAdder U183 (w661, w650, IN28[5], w662, w663);
  FullAdder U184 (w663, w652, IN29[4], w664, w665);
  FullAdder U185 (w665, w654, IN30[3], w666, w667);
  FullAdder U186 (w667, w656, IN31[2], w668, w669);
  FullAdder U187 (w669, w658, IN32[1], w670, w671);
  FullAdder U188 (w671, w659, IN33[0], w672, w673);
  HalfAdder U189 (w662, IN28[6], Out1[28], w675);
  FullAdder U190 (w675, w664, IN29[5], w676, w677);
  FullAdder U191 (w677, w666, IN30[4], w678, w679);
  FullAdder U192 (w679, w668, IN31[3], w680, w681);
  FullAdder U193 (w681, w670, IN32[2], w682, w683);
  FullAdder U194 (w683, w672, IN33[1], w684, w685);
  FullAdder U195 (w685, w673, IN34[0], w686, w687);
  HalfAdder U196 (w676, IN29[6], Out1[29], w689);
  FullAdder U197 (w689, w678, IN30[5], w690, w691);
  FullAdder U198 (w691, w680, IN31[4], w692, w693);
  FullAdder U199 (w693, w682, IN32[3], w694, w695);
  FullAdder U200 (w695, w684, IN33[2], w696, w697);
  FullAdder U201 (w697, w686, IN34[1], w698, w699);
  FullAdder U202 (w699, w687, IN35[0], w700, w701);
  HalfAdder U203 (w690, IN30[6], Out1[30], w703);
  FullAdder U204 (w703, w692, IN31[5], w704, w705);
  FullAdder U205 (w705, w694, IN32[4], w706, w707);
  FullAdder U206 (w707, w696, IN33[3], w708, w709);
  FullAdder U207 (w709, w698, IN34[2], w710, w711);
  FullAdder U208 (w711, w700, IN35[1], w712, w713);
  FullAdder U209 (w713, w701, IN36[0], w714, w715);
  HalfAdder U210 (w704, IN31[6], Out1[31], w717);
  FullAdder U211 (w717, w706, IN32[5], w718, w719);
  FullAdder U212 (w719, w708, IN33[4], w720, w721);
  FullAdder U213 (w721, w710, IN34[3], w722, w723);
  FullAdder U214 (w723, w712, IN35[2], w724, w725);
  FullAdder U215 (w725, w714, IN36[1], w726, w727);
  FullAdder U216 (w727, w715, IN37[0], w728, w729);
  HalfAdder U217 (w718, IN32[6], Out1[32], w731);
  FullAdder U218 (w731, w720, IN33[5], w732, w733);
  FullAdder U219 (w733, w722, IN34[4], w734, w735);
  FullAdder U220 (w735, w724, IN35[3], w736, w737);
  FullAdder U221 (w737, w726, IN36[2], w738, w739);
  FullAdder U222 (w739, w728, IN37[1], w740, w741);
  FullAdder U223 (w741, w729, IN38[0], w742, w743);
  HalfAdder U224 (w732, IN33[6], Out1[33], w745);
  FullAdder U225 (w745, w734, IN34[5], w746, w747);
  FullAdder U226 (w747, w736, IN35[4], w748, w749);
  FullAdder U227 (w749, w738, IN36[3], w750, w751);
  FullAdder U228 (w751, w740, IN37[2], w752, w753);
  FullAdder U229 (w753, w742, IN38[1], w754, w755);
  FullAdder U230 (w755, w743, IN39[0], w756, w757);
  HalfAdder U231 (w746, IN34[6], Out1[34], w759);
  FullAdder U232 (w759, w748, IN35[5], w760, w761);
  FullAdder U233 (w761, w750, IN36[4], w762, w763);
  FullAdder U234 (w763, w752, IN37[3], w764, w765);
  FullAdder U235 (w765, w754, IN38[2], w766, w767);
  FullAdder U236 (w767, w756, IN39[1], w768, w769);
  FullAdder U237 (w769, w757, IN40[0], w770, w771);
  HalfAdder U238 (w760, IN35[6], Out1[35], w773);
  FullAdder U239 (w773, w762, IN36[5], w774, w775);
  FullAdder U240 (w775, w764, IN37[4], w776, w777);
  FullAdder U241 (w777, w766, IN38[3], w778, w779);
  FullAdder U242 (w779, w768, IN39[2], w780, w781);
  FullAdder U243 (w781, w770, IN40[1], w782, w783);
  FullAdder U244 (w783, w771, IN41[0], w784, w785);
  HalfAdder U245 (w774, IN36[6], Out1[36], w787);
  FullAdder U246 (w787, w776, IN37[5], Out1[37], w789);
  FullAdder U247 (w789, w778, IN38[4], Out1[38], w791);
  FullAdder U248 (w791, w780, IN39[3], Out1[39], w793);
  FullAdder U249 (w793, w782, IN40[2], Out1[40], w795);
  FullAdder U250 (w795, w784, IN41[1], Out1[41], w797);
  FullAdder U251 (w797, w785, IN42[0], Out1[42], Out1[43]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN8[7];
  assign Out2[1] = IN9[7];
  assign Out2[2] = IN10[7];
  assign Out2[3] = IN11[7];
  assign Out2[4] = IN12[7];
  assign Out2[5] = IN13[7];
  assign Out2[6] = IN14[7];
  assign Out2[7] = IN15[7];
  assign Out2[8] = IN16[7];
  assign Out2[9] = IN17[7];
  assign Out2[10] = IN18[7];
  assign Out2[11] = IN19[7];
  assign Out2[12] = IN20[7];
  assign Out2[13] = IN21[7];
  assign Out2[14] = IN22[7];
  assign Out2[15] = IN23[7];
  assign Out2[16] = IN24[7];
  assign Out2[17] = IN25[7];
  assign Out2[18] = IN26[7];
  assign Out2[19] = IN27[7];
  assign Out2[20] = IN28[7];
  assign Out2[21] = IN29[7];
  assign Out2[22] = IN30[7];
  assign Out2[23] = IN31[7];
  assign Out2[24] = IN32[7];
  assign Out2[25] = IN33[7];
  assign Out2[26] = IN34[7];
  assign Out2[27] = IN35[7];
  assign Out2[28] = IN36[7];
  assign Out2[29] = IN37[6];
  assign Out2[30] = IN38[5];
  assign Out2[31] = IN39[4];
  assign Out2[32] = IN40[3];
  assign Out2[33] = IN41[2];
  assign Out2[34] = IN42[1];
  assign Out2[35] = IN43[0];

endmodule
module RC_36_36(IN1, IN2, Out);
  input [35:0] IN1;
  input [35:0] IN2;
  output [36:0] Out;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w73);
  FullAdder U1 (IN1[1], IN2[1], w73, Out[1], w75);
  FullAdder U2 (IN1[2], IN2[2], w75, Out[2], w77);
  FullAdder U3 (IN1[3], IN2[3], w77, Out[3], w79);
  FullAdder U4 (IN1[4], IN2[4], w79, Out[4], w81);
  FullAdder U5 (IN1[5], IN2[5], w81, Out[5], w83);
  FullAdder U6 (IN1[6], IN2[6], w83, Out[6], w85);
  FullAdder U7 (IN1[7], IN2[7], w85, Out[7], w87);
  FullAdder U8 (IN1[8], IN2[8], w87, Out[8], w89);
  FullAdder U9 (IN1[9], IN2[9], w89, Out[9], w91);
  FullAdder U10 (IN1[10], IN2[10], w91, Out[10], w93);
  FullAdder U11 (IN1[11], IN2[11], w93, Out[11], w95);
  FullAdder U12 (IN1[12], IN2[12], w95, Out[12], w97);
  FullAdder U13 (IN1[13], IN2[13], w97, Out[13], w99);
  FullAdder U14 (IN1[14], IN2[14], w99, Out[14], w101);
  FullAdder U15 (IN1[15], IN2[15], w101, Out[15], w103);
  FullAdder U16 (IN1[16], IN2[16], w103, Out[16], w105);
  FullAdder U17 (IN1[17], IN2[17], w105, Out[17], w107);
  FullAdder U18 (IN1[18], IN2[18], w107, Out[18], w109);
  FullAdder U19 (IN1[19], IN2[19], w109, Out[19], w111);
  FullAdder U20 (IN1[20], IN2[20], w111, Out[20], w113);
  FullAdder U21 (IN1[21], IN2[21], w113, Out[21], w115);
  FullAdder U22 (IN1[22], IN2[22], w115, Out[22], w117);
  FullAdder U23 (IN1[23], IN2[23], w117, Out[23], w119);
  FullAdder U24 (IN1[24], IN2[24], w119, Out[24], w121);
  FullAdder U25 (IN1[25], IN2[25], w121, Out[25], w123);
  FullAdder U26 (IN1[26], IN2[26], w123, Out[26], w125);
  FullAdder U27 (IN1[27], IN2[27], w125, Out[27], w127);
  FullAdder U28 (IN1[28], IN2[28], w127, Out[28], w129);
  FullAdder U29 (IN1[29], IN2[29], w129, Out[29], w131);
  FullAdder U30 (IN1[30], IN2[30], w131, Out[30], w133);
  FullAdder U31 (IN1[31], IN2[31], w133, Out[31], w135);
  FullAdder U32 (IN1[32], IN2[32], w135, Out[32], w137);
  FullAdder U33 (IN1[33], IN2[33], w137, Out[33], w139);
  FullAdder U34 (IN1[34], IN2[34], w139, Out[34], w141);
  FullAdder U35 (IN1[35], IN2[35], w141, Out[35], Out[36]);

endmodule
module NR_8_37(IN1, IN2, Out);
  input [7:0] IN1;
  input [36:0] IN2;
  output [44:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [7:0] P8;
  wire [7:0] P9;
  wire [7:0] P10;
  wire [7:0] P11;
  wire [7:0] P12;
  wire [7:0] P13;
  wire [7:0] P14;
  wire [7:0] P15;
  wire [7:0] P16;
  wire [7:0] P17;
  wire [7:0] P18;
  wire [7:0] P19;
  wire [7:0] P20;
  wire [7:0] P21;
  wire [7:0] P22;
  wire [7:0] P23;
  wire [7:0] P24;
  wire [7:0] P25;
  wire [7:0] P26;
  wire [7:0] P27;
  wire [7:0] P28;
  wire [7:0] P29;
  wire [7:0] P30;
  wire [7:0] P31;
  wire [7:0] P32;
  wire [7:0] P33;
  wire [7:0] P34;
  wire [7:0] P35;
  wire [7:0] P36;
  wire [6:0] P37;
  wire [5:0] P38;
  wire [4:0] P39;
  wire [3:0] P40;
  wire [2:0] P41;
  wire [1:0] P42;
  wire [0:0] P43;
  wire [43:0] R1;
  wire [35:0] R2;
  wire [44:0] aOut;
  U_SP_8_37 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, R1, R2);
  RC_36_36 S2 (R1[43:8], R2, aOut[44:8]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign Out = aOut[44:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
