
module NR_57_1(
    input [56:0]IN1,
    input [0:0]IN2,
    output [56:0]Out
);
    assign Out = IN2;
endmodule
