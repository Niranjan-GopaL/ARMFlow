
module customAdder64_0(
    input [63 : 0] A,
    input [63 : 0] B,
    output [64 : 0] Sum
);

    assign Sum = A+B;

endmodule
