
module customAdder35_0(
    input [34 : 0] A,
    input [34 : 0] B,
    output [35 : 0] Sum
);

    assign Sum = A+B;

endmodule
