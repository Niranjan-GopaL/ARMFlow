
module customAdder50_0(
    input [49 : 0] A,
    input [49 : 0] B,
    output [50 : 0] Sum
);

    assign Sum = A+B;

endmodule
