//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 7
  second input length: 34
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_7_34(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39);
  input [6:0] IN1;
  input [33:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [5:0] P34;
  output [4:0] P35;
  output [3:0] P36;
  output [2:0] P37;
  output [1:0] P38;
  output [0:0] P39;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[0] = IN1[1]&IN2[33];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[1] = IN1[2]&IN2[32];
  assign P35[0] = IN1[2]&IN2[33];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[2] = IN1[3]&IN2[31];
  assign P35[1] = IN1[3]&IN2[32];
  assign P36[0] = IN1[3]&IN2[33];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[3] = IN1[4]&IN2[30];
  assign P35[2] = IN1[4]&IN2[31];
  assign P36[1] = IN1[4]&IN2[32];
  assign P37[0] = IN1[4]&IN2[33];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[4] = IN1[5]&IN2[29];
  assign P35[3] = IN1[5]&IN2[30];
  assign P36[2] = IN1[5]&IN2[31];
  assign P37[1] = IN1[5]&IN2[32];
  assign P38[0] = IN1[5]&IN2[33];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[5] = IN1[6]&IN2[28];
  assign P35[4] = IN1[6]&IN2[29];
  assign P36[3] = IN1[6]&IN2[30];
  assign P37[2] = IN1[6]&IN2[31];
  assign P38[1] = IN1[6]&IN2[32];
  assign P39[0] = IN1[6]&IN2[33];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [5:0] IN34;
  input [4:0] IN35;
  input [3:0] IN36;
  input [2:0] IN37;
  input [1:0] IN38;
  input [0:0] IN39;
  output [39:0] Out1;
  output [32:0] Out2;
  wire w239;
  wire w240;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w246;
  wire w247;
  wire w248;
  wire w249;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w623;
  wire w625;
  wire w627;
  wire w629;
  wire w631;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w239);
  FullAdder U1 (w239, IN2[0], IN2[1], w240, w241);
  FullAdder U2 (w241, IN3[0], IN3[1], w242, w243);
  FullAdder U3 (w243, IN4[0], IN4[1], w244, w245);
  FullAdder U4 (w245, IN5[0], IN5[1], w246, w247);
  FullAdder U5 (w247, IN6[0], IN6[1], w248, w249);
  HalfAdder U6 (w240, IN2[2], Out1[2], w251);
  FullAdder U7 (w251, w242, IN3[2], w252, w253);
  FullAdder U8 (w253, w244, IN4[2], w254, w255);
  FullAdder U9 (w255, w246, IN5[2], w256, w257);
  FullAdder U10 (w257, w248, IN6[2], w258, w259);
  FullAdder U11 (w259, w249, IN7[0], w260, w261);
  HalfAdder U12 (w252, IN3[3], Out1[3], w263);
  FullAdder U13 (w263, w254, IN4[3], w264, w265);
  FullAdder U14 (w265, w256, IN5[3], w266, w267);
  FullAdder U15 (w267, w258, IN6[3], w268, w269);
  FullAdder U16 (w269, w260, IN7[1], w270, w271);
  FullAdder U17 (w271, w261, IN8[0], w272, w273);
  HalfAdder U18 (w264, IN4[4], Out1[4], w275);
  FullAdder U19 (w275, w266, IN5[4], w276, w277);
  FullAdder U20 (w277, w268, IN6[4], w278, w279);
  FullAdder U21 (w279, w270, IN7[2], w280, w281);
  FullAdder U22 (w281, w272, IN8[1], w282, w283);
  FullAdder U23 (w283, w273, IN9[0], w284, w285);
  HalfAdder U24 (w276, IN5[5], Out1[5], w287);
  FullAdder U25 (w287, w278, IN6[5], w288, w289);
  FullAdder U26 (w289, w280, IN7[3], w290, w291);
  FullAdder U27 (w291, w282, IN8[2], w292, w293);
  FullAdder U28 (w293, w284, IN9[1], w294, w295);
  FullAdder U29 (w295, w285, IN10[0], w296, w297);
  HalfAdder U30 (w288, IN6[6], Out1[6], w299);
  FullAdder U31 (w299, w290, IN7[4], w300, w301);
  FullAdder U32 (w301, w292, IN8[3], w302, w303);
  FullAdder U33 (w303, w294, IN9[2], w304, w305);
  FullAdder U34 (w305, w296, IN10[1], w306, w307);
  FullAdder U35 (w307, w297, IN11[0], w308, w309);
  HalfAdder U36 (w300, IN7[5], Out1[7], w311);
  FullAdder U37 (w311, w302, IN8[4], w312, w313);
  FullAdder U38 (w313, w304, IN9[3], w314, w315);
  FullAdder U39 (w315, w306, IN10[2], w316, w317);
  FullAdder U40 (w317, w308, IN11[1], w318, w319);
  FullAdder U41 (w319, w309, IN12[0], w320, w321);
  HalfAdder U42 (w312, IN8[5], Out1[8], w323);
  FullAdder U43 (w323, w314, IN9[4], w324, w325);
  FullAdder U44 (w325, w316, IN10[3], w326, w327);
  FullAdder U45 (w327, w318, IN11[2], w328, w329);
  FullAdder U46 (w329, w320, IN12[1], w330, w331);
  FullAdder U47 (w331, w321, IN13[0], w332, w333);
  HalfAdder U48 (w324, IN9[5], Out1[9], w335);
  FullAdder U49 (w335, w326, IN10[4], w336, w337);
  FullAdder U50 (w337, w328, IN11[3], w338, w339);
  FullAdder U51 (w339, w330, IN12[2], w340, w341);
  FullAdder U52 (w341, w332, IN13[1], w342, w343);
  FullAdder U53 (w343, w333, IN14[0], w344, w345);
  HalfAdder U54 (w336, IN10[5], Out1[10], w347);
  FullAdder U55 (w347, w338, IN11[4], w348, w349);
  FullAdder U56 (w349, w340, IN12[3], w350, w351);
  FullAdder U57 (w351, w342, IN13[2], w352, w353);
  FullAdder U58 (w353, w344, IN14[1], w354, w355);
  FullAdder U59 (w355, w345, IN15[0], w356, w357);
  HalfAdder U60 (w348, IN11[5], Out1[11], w359);
  FullAdder U61 (w359, w350, IN12[4], w360, w361);
  FullAdder U62 (w361, w352, IN13[3], w362, w363);
  FullAdder U63 (w363, w354, IN14[2], w364, w365);
  FullAdder U64 (w365, w356, IN15[1], w366, w367);
  FullAdder U65 (w367, w357, IN16[0], w368, w369);
  HalfAdder U66 (w360, IN12[5], Out1[12], w371);
  FullAdder U67 (w371, w362, IN13[4], w372, w373);
  FullAdder U68 (w373, w364, IN14[3], w374, w375);
  FullAdder U69 (w375, w366, IN15[2], w376, w377);
  FullAdder U70 (w377, w368, IN16[1], w378, w379);
  FullAdder U71 (w379, w369, IN17[0], w380, w381);
  HalfAdder U72 (w372, IN13[5], Out1[13], w383);
  FullAdder U73 (w383, w374, IN14[4], w384, w385);
  FullAdder U74 (w385, w376, IN15[3], w386, w387);
  FullAdder U75 (w387, w378, IN16[2], w388, w389);
  FullAdder U76 (w389, w380, IN17[1], w390, w391);
  FullAdder U77 (w391, w381, IN18[0], w392, w393);
  HalfAdder U78 (w384, IN14[5], Out1[14], w395);
  FullAdder U79 (w395, w386, IN15[4], w396, w397);
  FullAdder U80 (w397, w388, IN16[3], w398, w399);
  FullAdder U81 (w399, w390, IN17[2], w400, w401);
  FullAdder U82 (w401, w392, IN18[1], w402, w403);
  FullAdder U83 (w403, w393, IN19[0], w404, w405);
  HalfAdder U84 (w396, IN15[5], Out1[15], w407);
  FullAdder U85 (w407, w398, IN16[4], w408, w409);
  FullAdder U86 (w409, w400, IN17[3], w410, w411);
  FullAdder U87 (w411, w402, IN18[2], w412, w413);
  FullAdder U88 (w413, w404, IN19[1], w414, w415);
  FullAdder U89 (w415, w405, IN20[0], w416, w417);
  HalfAdder U90 (w408, IN16[5], Out1[16], w419);
  FullAdder U91 (w419, w410, IN17[4], w420, w421);
  FullAdder U92 (w421, w412, IN18[3], w422, w423);
  FullAdder U93 (w423, w414, IN19[2], w424, w425);
  FullAdder U94 (w425, w416, IN20[1], w426, w427);
  FullAdder U95 (w427, w417, IN21[0], w428, w429);
  HalfAdder U96 (w420, IN17[5], Out1[17], w431);
  FullAdder U97 (w431, w422, IN18[4], w432, w433);
  FullAdder U98 (w433, w424, IN19[3], w434, w435);
  FullAdder U99 (w435, w426, IN20[2], w436, w437);
  FullAdder U100 (w437, w428, IN21[1], w438, w439);
  FullAdder U101 (w439, w429, IN22[0], w440, w441);
  HalfAdder U102 (w432, IN18[5], Out1[18], w443);
  FullAdder U103 (w443, w434, IN19[4], w444, w445);
  FullAdder U104 (w445, w436, IN20[3], w446, w447);
  FullAdder U105 (w447, w438, IN21[2], w448, w449);
  FullAdder U106 (w449, w440, IN22[1], w450, w451);
  FullAdder U107 (w451, w441, IN23[0], w452, w453);
  HalfAdder U108 (w444, IN19[5], Out1[19], w455);
  FullAdder U109 (w455, w446, IN20[4], w456, w457);
  FullAdder U110 (w457, w448, IN21[3], w458, w459);
  FullAdder U111 (w459, w450, IN22[2], w460, w461);
  FullAdder U112 (w461, w452, IN23[1], w462, w463);
  FullAdder U113 (w463, w453, IN24[0], w464, w465);
  HalfAdder U114 (w456, IN20[5], Out1[20], w467);
  FullAdder U115 (w467, w458, IN21[4], w468, w469);
  FullAdder U116 (w469, w460, IN22[3], w470, w471);
  FullAdder U117 (w471, w462, IN23[2], w472, w473);
  FullAdder U118 (w473, w464, IN24[1], w474, w475);
  FullAdder U119 (w475, w465, IN25[0], w476, w477);
  HalfAdder U120 (w468, IN21[5], Out1[21], w479);
  FullAdder U121 (w479, w470, IN22[4], w480, w481);
  FullAdder U122 (w481, w472, IN23[3], w482, w483);
  FullAdder U123 (w483, w474, IN24[2], w484, w485);
  FullAdder U124 (w485, w476, IN25[1], w486, w487);
  FullAdder U125 (w487, w477, IN26[0], w488, w489);
  HalfAdder U126 (w480, IN22[5], Out1[22], w491);
  FullAdder U127 (w491, w482, IN23[4], w492, w493);
  FullAdder U128 (w493, w484, IN24[3], w494, w495);
  FullAdder U129 (w495, w486, IN25[2], w496, w497);
  FullAdder U130 (w497, w488, IN26[1], w498, w499);
  FullAdder U131 (w499, w489, IN27[0], w500, w501);
  HalfAdder U132 (w492, IN23[5], Out1[23], w503);
  FullAdder U133 (w503, w494, IN24[4], w504, w505);
  FullAdder U134 (w505, w496, IN25[3], w506, w507);
  FullAdder U135 (w507, w498, IN26[2], w508, w509);
  FullAdder U136 (w509, w500, IN27[1], w510, w511);
  FullAdder U137 (w511, w501, IN28[0], w512, w513);
  HalfAdder U138 (w504, IN24[5], Out1[24], w515);
  FullAdder U139 (w515, w506, IN25[4], w516, w517);
  FullAdder U140 (w517, w508, IN26[3], w518, w519);
  FullAdder U141 (w519, w510, IN27[2], w520, w521);
  FullAdder U142 (w521, w512, IN28[1], w522, w523);
  FullAdder U143 (w523, w513, IN29[0], w524, w525);
  HalfAdder U144 (w516, IN25[5], Out1[25], w527);
  FullAdder U145 (w527, w518, IN26[4], w528, w529);
  FullAdder U146 (w529, w520, IN27[3], w530, w531);
  FullAdder U147 (w531, w522, IN28[2], w532, w533);
  FullAdder U148 (w533, w524, IN29[1], w534, w535);
  FullAdder U149 (w535, w525, IN30[0], w536, w537);
  HalfAdder U150 (w528, IN26[5], Out1[26], w539);
  FullAdder U151 (w539, w530, IN27[4], w540, w541);
  FullAdder U152 (w541, w532, IN28[3], w542, w543);
  FullAdder U153 (w543, w534, IN29[2], w544, w545);
  FullAdder U154 (w545, w536, IN30[1], w546, w547);
  FullAdder U155 (w547, w537, IN31[0], w548, w549);
  HalfAdder U156 (w540, IN27[5], Out1[27], w551);
  FullAdder U157 (w551, w542, IN28[4], w552, w553);
  FullAdder U158 (w553, w544, IN29[3], w554, w555);
  FullAdder U159 (w555, w546, IN30[2], w556, w557);
  FullAdder U160 (w557, w548, IN31[1], w558, w559);
  FullAdder U161 (w559, w549, IN32[0], w560, w561);
  HalfAdder U162 (w552, IN28[5], Out1[28], w563);
  FullAdder U163 (w563, w554, IN29[4], w564, w565);
  FullAdder U164 (w565, w556, IN30[3], w566, w567);
  FullAdder U165 (w567, w558, IN31[2], w568, w569);
  FullAdder U166 (w569, w560, IN32[1], w570, w571);
  FullAdder U167 (w571, w561, IN33[0], w572, w573);
  HalfAdder U168 (w564, IN29[5], Out1[29], w575);
  FullAdder U169 (w575, w566, IN30[4], w576, w577);
  FullAdder U170 (w577, w568, IN31[3], w578, w579);
  FullAdder U171 (w579, w570, IN32[2], w580, w581);
  FullAdder U172 (w581, w572, IN33[1], w582, w583);
  FullAdder U173 (w583, w573, IN34[0], w584, w585);
  HalfAdder U174 (w576, IN30[5], Out1[30], w587);
  FullAdder U175 (w587, w578, IN31[4], w588, w589);
  FullAdder U176 (w589, w580, IN32[3], w590, w591);
  FullAdder U177 (w591, w582, IN33[2], w592, w593);
  FullAdder U178 (w593, w584, IN34[1], w594, w595);
  FullAdder U179 (w595, w585, IN35[0], w596, w597);
  HalfAdder U180 (w588, IN31[5], Out1[31], w599);
  FullAdder U181 (w599, w590, IN32[4], w600, w601);
  FullAdder U182 (w601, w592, IN33[3], w602, w603);
  FullAdder U183 (w603, w594, IN34[2], w604, w605);
  FullAdder U184 (w605, w596, IN35[1], w606, w607);
  FullAdder U185 (w607, w597, IN36[0], w608, w609);
  HalfAdder U186 (w600, IN32[5], Out1[32], w611);
  FullAdder U187 (w611, w602, IN33[4], w612, w613);
  FullAdder U188 (w613, w604, IN34[3], w614, w615);
  FullAdder U189 (w615, w606, IN35[2], w616, w617);
  FullAdder U190 (w617, w608, IN36[1], w618, w619);
  FullAdder U191 (w619, w609, IN37[0], w620, w621);
  HalfAdder U192 (w612, IN33[5], Out1[33], w623);
  FullAdder U193 (w623, w614, IN34[4], Out1[34], w625);
  FullAdder U194 (w625, w616, IN35[3], Out1[35], w627);
  FullAdder U195 (w627, w618, IN36[2], Out1[36], w629);
  FullAdder U196 (w629, w620, IN37[1], Out1[37], w631);
  FullAdder U197 (w631, w621, IN38[0], Out1[38], Out1[39]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN7[6];
  assign Out2[1] = IN8[6];
  assign Out2[2] = IN9[6];
  assign Out2[3] = IN10[6];
  assign Out2[4] = IN11[6];
  assign Out2[5] = IN12[6];
  assign Out2[6] = IN13[6];
  assign Out2[7] = IN14[6];
  assign Out2[8] = IN15[6];
  assign Out2[9] = IN16[6];
  assign Out2[10] = IN17[6];
  assign Out2[11] = IN18[6];
  assign Out2[12] = IN19[6];
  assign Out2[13] = IN20[6];
  assign Out2[14] = IN21[6];
  assign Out2[15] = IN22[6];
  assign Out2[16] = IN23[6];
  assign Out2[17] = IN24[6];
  assign Out2[18] = IN25[6];
  assign Out2[19] = IN26[6];
  assign Out2[20] = IN27[6];
  assign Out2[21] = IN28[6];
  assign Out2[22] = IN29[6];
  assign Out2[23] = IN30[6];
  assign Out2[24] = IN31[6];
  assign Out2[25] = IN32[6];
  assign Out2[26] = IN33[6];
  assign Out2[27] = IN34[5];
  assign Out2[28] = IN35[4];
  assign Out2[29] = IN36[3];
  assign Out2[30] = IN37[2];
  assign Out2[31] = IN38[1];
  assign Out2[32] = IN39[0];

endmodule
module RC_33_33(IN1, IN2, Out);
  input [32:0] IN1;
  input [32:0] IN2;
  output [33:0] Out;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w67);
  FullAdder U1 (IN1[1], IN2[1], w67, Out[1], w69);
  FullAdder U2 (IN1[2], IN2[2], w69, Out[2], w71);
  FullAdder U3 (IN1[3], IN2[3], w71, Out[3], w73);
  FullAdder U4 (IN1[4], IN2[4], w73, Out[4], w75);
  FullAdder U5 (IN1[5], IN2[5], w75, Out[5], w77);
  FullAdder U6 (IN1[6], IN2[6], w77, Out[6], w79);
  FullAdder U7 (IN1[7], IN2[7], w79, Out[7], w81);
  FullAdder U8 (IN1[8], IN2[8], w81, Out[8], w83);
  FullAdder U9 (IN1[9], IN2[9], w83, Out[9], w85);
  FullAdder U10 (IN1[10], IN2[10], w85, Out[10], w87);
  FullAdder U11 (IN1[11], IN2[11], w87, Out[11], w89);
  FullAdder U12 (IN1[12], IN2[12], w89, Out[12], w91);
  FullAdder U13 (IN1[13], IN2[13], w91, Out[13], w93);
  FullAdder U14 (IN1[14], IN2[14], w93, Out[14], w95);
  FullAdder U15 (IN1[15], IN2[15], w95, Out[15], w97);
  FullAdder U16 (IN1[16], IN2[16], w97, Out[16], w99);
  FullAdder U17 (IN1[17], IN2[17], w99, Out[17], w101);
  FullAdder U18 (IN1[18], IN2[18], w101, Out[18], w103);
  FullAdder U19 (IN1[19], IN2[19], w103, Out[19], w105);
  FullAdder U20 (IN1[20], IN2[20], w105, Out[20], w107);
  FullAdder U21 (IN1[21], IN2[21], w107, Out[21], w109);
  FullAdder U22 (IN1[22], IN2[22], w109, Out[22], w111);
  FullAdder U23 (IN1[23], IN2[23], w111, Out[23], w113);
  FullAdder U24 (IN1[24], IN2[24], w113, Out[24], w115);
  FullAdder U25 (IN1[25], IN2[25], w115, Out[25], w117);
  FullAdder U26 (IN1[26], IN2[26], w117, Out[26], w119);
  FullAdder U27 (IN1[27], IN2[27], w119, Out[27], w121);
  FullAdder U28 (IN1[28], IN2[28], w121, Out[28], w123);
  FullAdder U29 (IN1[29], IN2[29], w123, Out[29], w125);
  FullAdder U30 (IN1[30], IN2[30], w125, Out[30], w127);
  FullAdder U31 (IN1[31], IN2[31], w127, Out[31], w129);
  FullAdder U32 (IN1[32], IN2[32], w129, Out[32], Out[33]);

endmodule
module NR_7_34(IN1, IN2, Out);
  input [6:0] IN1;
  input [33:0] IN2;
  output [40:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [5:0] P34;
  wire [4:0] P35;
  wire [3:0] P36;
  wire [2:0] P37;
  wire [1:0] P38;
  wire [0:0] P39;
  wire [39:0] R1;
  wire [32:0] R2;
  wire [40:0] aOut;
  U_SP_7_34 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, R1, R2);
  RC_33_33 S2 (R1[39:7], R2, aOut[40:7]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign Out = aOut[40:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
