
module customAdder47_0(
    input [46 : 0] A,
    input [46 : 0] B,
    output [47 : 0] Sum
);

    assign Sum = A+B;

endmodule
