
module NR_48_1(
    input [47:0]IN1,
    input [0:0]IN2,
    output [47:0]Out
);
    assign Out = IN2;
endmodule
