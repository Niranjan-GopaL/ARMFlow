
module customAdder51_0(
    input [50 : 0] A,
    input [50 : 0] B,
    output [51 : 0] Sum
);

    assign Sum = A+B;

endmodule
