
module customAdder39_0(
    input [38 : 0] A,
    input [38 : 0] B,
    output [39 : 0] Sum
);

    assign Sum = A+B;

endmodule
