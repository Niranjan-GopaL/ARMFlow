
module NR_56_1(
    input [55:0]IN1,
    input [0:0]IN2,
    output [55:0]Out
);
    assign Out = IN2;
endmodule
