
module customAdder54_0(
    input [53 : 0] A,
    input [53 : 0] B,
    output [54 : 0] Sum
);

    assign Sum = A+B;

endmodule
