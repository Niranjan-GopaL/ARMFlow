
module NR_1_35(
    input [0:0]IN1,
    input [34:0]IN2,
    output [34:0]Out
);
    assign Out = IN2;
endmodule
