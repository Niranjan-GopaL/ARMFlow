
module NR_41_1(
    input [40:0]IN1,
    input [0:0]IN2,
    output [40:0]Out
);
    assign Out = IN2;
endmodule
