
module customAdder59_0(
    input [58 : 0] A,
    input [58 : 0] B,
    output [59 : 0] Sum
);

    assign Sum = A+B;

endmodule
