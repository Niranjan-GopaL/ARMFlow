
module NR_1_45(
    input [0:0]IN1,
    input [44:0]IN2,
    output [44:0]Out
);
    assign Out = IN2;
endmodule
