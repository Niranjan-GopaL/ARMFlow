//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 58
  second input length: 63
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_58_63(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, P112, P113, P114, P115, P116, P117, P118, P119);
  input [57:0] IN1;
  input [62:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [29:0] P29;
  output [30:0] P30;
  output [31:0] P31;
  output [32:0] P32;
  output [33:0] P33;
  output [34:0] P34;
  output [35:0] P35;
  output [36:0] P36;
  output [37:0] P37;
  output [38:0] P38;
  output [39:0] P39;
  output [40:0] P40;
  output [41:0] P41;
  output [42:0] P42;
  output [43:0] P43;
  output [44:0] P44;
  output [45:0] P45;
  output [46:0] P46;
  output [47:0] P47;
  output [48:0] P48;
  output [49:0] P49;
  output [50:0] P50;
  output [51:0] P51;
  output [52:0] P52;
  output [53:0] P53;
  output [54:0] P54;
  output [55:0] P55;
  output [56:0] P56;
  output [57:0] P57;
  output [57:0] P58;
  output [57:0] P59;
  output [57:0] P60;
  output [57:0] P61;
  output [57:0] P62;
  output [56:0] P63;
  output [55:0] P64;
  output [54:0] P65;
  output [53:0] P66;
  output [52:0] P67;
  output [51:0] P68;
  output [50:0] P69;
  output [49:0] P70;
  output [48:0] P71;
  output [47:0] P72;
  output [46:0] P73;
  output [45:0] P74;
  output [44:0] P75;
  output [43:0] P76;
  output [42:0] P77;
  output [41:0] P78;
  output [40:0] P79;
  output [39:0] P80;
  output [38:0] P81;
  output [37:0] P82;
  output [36:0] P83;
  output [35:0] P84;
  output [34:0] P85;
  output [33:0] P86;
  output [32:0] P87;
  output [31:0] P88;
  output [30:0] P89;
  output [29:0] P90;
  output [28:0] P91;
  output [27:0] P92;
  output [26:0] P93;
  output [25:0] P94;
  output [24:0] P95;
  output [23:0] P96;
  output [22:0] P97;
  output [21:0] P98;
  output [20:0] P99;
  output [19:0] P100;
  output [18:0] P101;
  output [17:0] P102;
  output [16:0] P103;
  output [15:0] P104;
  output [14:0] P105;
  output [13:0] P106;
  output [12:0] P107;
  output [11:0] P108;
  output [10:0] P109;
  output [9:0] P110;
  output [8:0] P111;
  output [7:0] P112;
  output [6:0] P113;
  output [5:0] P114;
  output [4:0] P115;
  output [3:0] P116;
  output [2:0] P117;
  output [1:0] P118;
  output [0:0] P119;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P54[0] = IN1[0]&IN2[54];
  assign P55[0] = IN1[0]&IN2[55];
  assign P56[0] = IN1[0]&IN2[56];
  assign P57[0] = IN1[0]&IN2[57];
  assign P58[0] = IN1[0]&IN2[58];
  assign P59[0] = IN1[0]&IN2[59];
  assign P60[0] = IN1[0]&IN2[60];
  assign P61[0] = IN1[0]&IN2[61];
  assign P62[0] = IN1[0]&IN2[62];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[1] = IN1[1]&IN2[53];
  assign P55[1] = IN1[1]&IN2[54];
  assign P56[1] = IN1[1]&IN2[55];
  assign P57[1] = IN1[1]&IN2[56];
  assign P58[1] = IN1[1]&IN2[57];
  assign P59[1] = IN1[1]&IN2[58];
  assign P60[1] = IN1[1]&IN2[59];
  assign P61[1] = IN1[1]&IN2[60];
  assign P62[1] = IN1[1]&IN2[61];
  assign P63[0] = IN1[1]&IN2[62];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[2] = IN1[2]&IN2[52];
  assign P55[2] = IN1[2]&IN2[53];
  assign P56[2] = IN1[2]&IN2[54];
  assign P57[2] = IN1[2]&IN2[55];
  assign P58[2] = IN1[2]&IN2[56];
  assign P59[2] = IN1[2]&IN2[57];
  assign P60[2] = IN1[2]&IN2[58];
  assign P61[2] = IN1[2]&IN2[59];
  assign P62[2] = IN1[2]&IN2[60];
  assign P63[1] = IN1[2]&IN2[61];
  assign P64[0] = IN1[2]&IN2[62];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[3] = IN1[3]&IN2[51];
  assign P55[3] = IN1[3]&IN2[52];
  assign P56[3] = IN1[3]&IN2[53];
  assign P57[3] = IN1[3]&IN2[54];
  assign P58[3] = IN1[3]&IN2[55];
  assign P59[3] = IN1[3]&IN2[56];
  assign P60[3] = IN1[3]&IN2[57];
  assign P61[3] = IN1[3]&IN2[58];
  assign P62[3] = IN1[3]&IN2[59];
  assign P63[2] = IN1[3]&IN2[60];
  assign P64[1] = IN1[3]&IN2[61];
  assign P65[0] = IN1[3]&IN2[62];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[4] = IN1[4]&IN2[50];
  assign P55[4] = IN1[4]&IN2[51];
  assign P56[4] = IN1[4]&IN2[52];
  assign P57[4] = IN1[4]&IN2[53];
  assign P58[4] = IN1[4]&IN2[54];
  assign P59[4] = IN1[4]&IN2[55];
  assign P60[4] = IN1[4]&IN2[56];
  assign P61[4] = IN1[4]&IN2[57];
  assign P62[4] = IN1[4]&IN2[58];
  assign P63[3] = IN1[4]&IN2[59];
  assign P64[2] = IN1[4]&IN2[60];
  assign P65[1] = IN1[4]&IN2[61];
  assign P66[0] = IN1[4]&IN2[62];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[5] = IN1[5]&IN2[49];
  assign P55[5] = IN1[5]&IN2[50];
  assign P56[5] = IN1[5]&IN2[51];
  assign P57[5] = IN1[5]&IN2[52];
  assign P58[5] = IN1[5]&IN2[53];
  assign P59[5] = IN1[5]&IN2[54];
  assign P60[5] = IN1[5]&IN2[55];
  assign P61[5] = IN1[5]&IN2[56];
  assign P62[5] = IN1[5]&IN2[57];
  assign P63[4] = IN1[5]&IN2[58];
  assign P64[3] = IN1[5]&IN2[59];
  assign P65[2] = IN1[5]&IN2[60];
  assign P66[1] = IN1[5]&IN2[61];
  assign P67[0] = IN1[5]&IN2[62];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[6] = IN1[6]&IN2[48];
  assign P55[6] = IN1[6]&IN2[49];
  assign P56[6] = IN1[6]&IN2[50];
  assign P57[6] = IN1[6]&IN2[51];
  assign P58[6] = IN1[6]&IN2[52];
  assign P59[6] = IN1[6]&IN2[53];
  assign P60[6] = IN1[6]&IN2[54];
  assign P61[6] = IN1[6]&IN2[55];
  assign P62[6] = IN1[6]&IN2[56];
  assign P63[5] = IN1[6]&IN2[57];
  assign P64[4] = IN1[6]&IN2[58];
  assign P65[3] = IN1[6]&IN2[59];
  assign P66[2] = IN1[6]&IN2[60];
  assign P67[1] = IN1[6]&IN2[61];
  assign P68[0] = IN1[6]&IN2[62];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[7] = IN1[7]&IN2[47];
  assign P55[7] = IN1[7]&IN2[48];
  assign P56[7] = IN1[7]&IN2[49];
  assign P57[7] = IN1[7]&IN2[50];
  assign P58[7] = IN1[7]&IN2[51];
  assign P59[7] = IN1[7]&IN2[52];
  assign P60[7] = IN1[7]&IN2[53];
  assign P61[7] = IN1[7]&IN2[54];
  assign P62[7] = IN1[7]&IN2[55];
  assign P63[6] = IN1[7]&IN2[56];
  assign P64[5] = IN1[7]&IN2[57];
  assign P65[4] = IN1[7]&IN2[58];
  assign P66[3] = IN1[7]&IN2[59];
  assign P67[2] = IN1[7]&IN2[60];
  assign P68[1] = IN1[7]&IN2[61];
  assign P69[0] = IN1[7]&IN2[62];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[8] = IN1[8]&IN2[45];
  assign P54[8] = IN1[8]&IN2[46];
  assign P55[8] = IN1[8]&IN2[47];
  assign P56[8] = IN1[8]&IN2[48];
  assign P57[8] = IN1[8]&IN2[49];
  assign P58[8] = IN1[8]&IN2[50];
  assign P59[8] = IN1[8]&IN2[51];
  assign P60[8] = IN1[8]&IN2[52];
  assign P61[8] = IN1[8]&IN2[53];
  assign P62[8] = IN1[8]&IN2[54];
  assign P63[7] = IN1[8]&IN2[55];
  assign P64[6] = IN1[8]&IN2[56];
  assign P65[5] = IN1[8]&IN2[57];
  assign P66[4] = IN1[8]&IN2[58];
  assign P67[3] = IN1[8]&IN2[59];
  assign P68[2] = IN1[8]&IN2[60];
  assign P69[1] = IN1[8]&IN2[61];
  assign P70[0] = IN1[8]&IN2[62];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[9] = IN1[9]&IN2[44];
  assign P54[9] = IN1[9]&IN2[45];
  assign P55[9] = IN1[9]&IN2[46];
  assign P56[9] = IN1[9]&IN2[47];
  assign P57[9] = IN1[9]&IN2[48];
  assign P58[9] = IN1[9]&IN2[49];
  assign P59[9] = IN1[9]&IN2[50];
  assign P60[9] = IN1[9]&IN2[51];
  assign P61[9] = IN1[9]&IN2[52];
  assign P62[9] = IN1[9]&IN2[53];
  assign P63[8] = IN1[9]&IN2[54];
  assign P64[7] = IN1[9]&IN2[55];
  assign P65[6] = IN1[9]&IN2[56];
  assign P66[5] = IN1[9]&IN2[57];
  assign P67[4] = IN1[9]&IN2[58];
  assign P68[3] = IN1[9]&IN2[59];
  assign P69[2] = IN1[9]&IN2[60];
  assign P70[1] = IN1[9]&IN2[61];
  assign P71[0] = IN1[9]&IN2[62];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[10] = IN1[10]&IN2[39];
  assign P50[10] = IN1[10]&IN2[40];
  assign P51[10] = IN1[10]&IN2[41];
  assign P52[10] = IN1[10]&IN2[42];
  assign P53[10] = IN1[10]&IN2[43];
  assign P54[10] = IN1[10]&IN2[44];
  assign P55[10] = IN1[10]&IN2[45];
  assign P56[10] = IN1[10]&IN2[46];
  assign P57[10] = IN1[10]&IN2[47];
  assign P58[10] = IN1[10]&IN2[48];
  assign P59[10] = IN1[10]&IN2[49];
  assign P60[10] = IN1[10]&IN2[50];
  assign P61[10] = IN1[10]&IN2[51];
  assign P62[10] = IN1[10]&IN2[52];
  assign P63[9] = IN1[10]&IN2[53];
  assign P64[8] = IN1[10]&IN2[54];
  assign P65[7] = IN1[10]&IN2[55];
  assign P66[6] = IN1[10]&IN2[56];
  assign P67[5] = IN1[10]&IN2[57];
  assign P68[4] = IN1[10]&IN2[58];
  assign P69[3] = IN1[10]&IN2[59];
  assign P70[2] = IN1[10]&IN2[60];
  assign P71[1] = IN1[10]&IN2[61];
  assign P72[0] = IN1[10]&IN2[62];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[11] = IN1[11]&IN2[38];
  assign P50[11] = IN1[11]&IN2[39];
  assign P51[11] = IN1[11]&IN2[40];
  assign P52[11] = IN1[11]&IN2[41];
  assign P53[11] = IN1[11]&IN2[42];
  assign P54[11] = IN1[11]&IN2[43];
  assign P55[11] = IN1[11]&IN2[44];
  assign P56[11] = IN1[11]&IN2[45];
  assign P57[11] = IN1[11]&IN2[46];
  assign P58[11] = IN1[11]&IN2[47];
  assign P59[11] = IN1[11]&IN2[48];
  assign P60[11] = IN1[11]&IN2[49];
  assign P61[11] = IN1[11]&IN2[50];
  assign P62[11] = IN1[11]&IN2[51];
  assign P63[10] = IN1[11]&IN2[52];
  assign P64[9] = IN1[11]&IN2[53];
  assign P65[8] = IN1[11]&IN2[54];
  assign P66[7] = IN1[11]&IN2[55];
  assign P67[6] = IN1[11]&IN2[56];
  assign P68[5] = IN1[11]&IN2[57];
  assign P69[4] = IN1[11]&IN2[58];
  assign P70[3] = IN1[11]&IN2[59];
  assign P71[2] = IN1[11]&IN2[60];
  assign P72[1] = IN1[11]&IN2[61];
  assign P73[0] = IN1[11]&IN2[62];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[12] = IN1[12]&IN2[37];
  assign P50[12] = IN1[12]&IN2[38];
  assign P51[12] = IN1[12]&IN2[39];
  assign P52[12] = IN1[12]&IN2[40];
  assign P53[12] = IN1[12]&IN2[41];
  assign P54[12] = IN1[12]&IN2[42];
  assign P55[12] = IN1[12]&IN2[43];
  assign P56[12] = IN1[12]&IN2[44];
  assign P57[12] = IN1[12]&IN2[45];
  assign P58[12] = IN1[12]&IN2[46];
  assign P59[12] = IN1[12]&IN2[47];
  assign P60[12] = IN1[12]&IN2[48];
  assign P61[12] = IN1[12]&IN2[49];
  assign P62[12] = IN1[12]&IN2[50];
  assign P63[11] = IN1[12]&IN2[51];
  assign P64[10] = IN1[12]&IN2[52];
  assign P65[9] = IN1[12]&IN2[53];
  assign P66[8] = IN1[12]&IN2[54];
  assign P67[7] = IN1[12]&IN2[55];
  assign P68[6] = IN1[12]&IN2[56];
  assign P69[5] = IN1[12]&IN2[57];
  assign P70[4] = IN1[12]&IN2[58];
  assign P71[3] = IN1[12]&IN2[59];
  assign P72[2] = IN1[12]&IN2[60];
  assign P73[1] = IN1[12]&IN2[61];
  assign P74[0] = IN1[12]&IN2[62];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[13] = IN1[13]&IN2[36];
  assign P50[13] = IN1[13]&IN2[37];
  assign P51[13] = IN1[13]&IN2[38];
  assign P52[13] = IN1[13]&IN2[39];
  assign P53[13] = IN1[13]&IN2[40];
  assign P54[13] = IN1[13]&IN2[41];
  assign P55[13] = IN1[13]&IN2[42];
  assign P56[13] = IN1[13]&IN2[43];
  assign P57[13] = IN1[13]&IN2[44];
  assign P58[13] = IN1[13]&IN2[45];
  assign P59[13] = IN1[13]&IN2[46];
  assign P60[13] = IN1[13]&IN2[47];
  assign P61[13] = IN1[13]&IN2[48];
  assign P62[13] = IN1[13]&IN2[49];
  assign P63[12] = IN1[13]&IN2[50];
  assign P64[11] = IN1[13]&IN2[51];
  assign P65[10] = IN1[13]&IN2[52];
  assign P66[9] = IN1[13]&IN2[53];
  assign P67[8] = IN1[13]&IN2[54];
  assign P68[7] = IN1[13]&IN2[55];
  assign P69[6] = IN1[13]&IN2[56];
  assign P70[5] = IN1[13]&IN2[57];
  assign P71[4] = IN1[13]&IN2[58];
  assign P72[3] = IN1[13]&IN2[59];
  assign P73[2] = IN1[13]&IN2[60];
  assign P74[1] = IN1[13]&IN2[61];
  assign P75[0] = IN1[13]&IN2[62];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[14] = IN1[14]&IN2[24];
  assign P39[14] = IN1[14]&IN2[25];
  assign P40[14] = IN1[14]&IN2[26];
  assign P41[14] = IN1[14]&IN2[27];
  assign P42[14] = IN1[14]&IN2[28];
  assign P43[14] = IN1[14]&IN2[29];
  assign P44[14] = IN1[14]&IN2[30];
  assign P45[14] = IN1[14]&IN2[31];
  assign P46[14] = IN1[14]&IN2[32];
  assign P47[14] = IN1[14]&IN2[33];
  assign P48[14] = IN1[14]&IN2[34];
  assign P49[14] = IN1[14]&IN2[35];
  assign P50[14] = IN1[14]&IN2[36];
  assign P51[14] = IN1[14]&IN2[37];
  assign P52[14] = IN1[14]&IN2[38];
  assign P53[14] = IN1[14]&IN2[39];
  assign P54[14] = IN1[14]&IN2[40];
  assign P55[14] = IN1[14]&IN2[41];
  assign P56[14] = IN1[14]&IN2[42];
  assign P57[14] = IN1[14]&IN2[43];
  assign P58[14] = IN1[14]&IN2[44];
  assign P59[14] = IN1[14]&IN2[45];
  assign P60[14] = IN1[14]&IN2[46];
  assign P61[14] = IN1[14]&IN2[47];
  assign P62[14] = IN1[14]&IN2[48];
  assign P63[13] = IN1[14]&IN2[49];
  assign P64[12] = IN1[14]&IN2[50];
  assign P65[11] = IN1[14]&IN2[51];
  assign P66[10] = IN1[14]&IN2[52];
  assign P67[9] = IN1[14]&IN2[53];
  assign P68[8] = IN1[14]&IN2[54];
  assign P69[7] = IN1[14]&IN2[55];
  assign P70[6] = IN1[14]&IN2[56];
  assign P71[5] = IN1[14]&IN2[57];
  assign P72[4] = IN1[14]&IN2[58];
  assign P73[3] = IN1[14]&IN2[59];
  assign P74[2] = IN1[14]&IN2[60];
  assign P75[1] = IN1[14]&IN2[61];
  assign P76[0] = IN1[14]&IN2[62];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[15] = IN1[15]&IN2[23];
  assign P39[15] = IN1[15]&IN2[24];
  assign P40[15] = IN1[15]&IN2[25];
  assign P41[15] = IN1[15]&IN2[26];
  assign P42[15] = IN1[15]&IN2[27];
  assign P43[15] = IN1[15]&IN2[28];
  assign P44[15] = IN1[15]&IN2[29];
  assign P45[15] = IN1[15]&IN2[30];
  assign P46[15] = IN1[15]&IN2[31];
  assign P47[15] = IN1[15]&IN2[32];
  assign P48[15] = IN1[15]&IN2[33];
  assign P49[15] = IN1[15]&IN2[34];
  assign P50[15] = IN1[15]&IN2[35];
  assign P51[15] = IN1[15]&IN2[36];
  assign P52[15] = IN1[15]&IN2[37];
  assign P53[15] = IN1[15]&IN2[38];
  assign P54[15] = IN1[15]&IN2[39];
  assign P55[15] = IN1[15]&IN2[40];
  assign P56[15] = IN1[15]&IN2[41];
  assign P57[15] = IN1[15]&IN2[42];
  assign P58[15] = IN1[15]&IN2[43];
  assign P59[15] = IN1[15]&IN2[44];
  assign P60[15] = IN1[15]&IN2[45];
  assign P61[15] = IN1[15]&IN2[46];
  assign P62[15] = IN1[15]&IN2[47];
  assign P63[14] = IN1[15]&IN2[48];
  assign P64[13] = IN1[15]&IN2[49];
  assign P65[12] = IN1[15]&IN2[50];
  assign P66[11] = IN1[15]&IN2[51];
  assign P67[10] = IN1[15]&IN2[52];
  assign P68[9] = IN1[15]&IN2[53];
  assign P69[8] = IN1[15]&IN2[54];
  assign P70[7] = IN1[15]&IN2[55];
  assign P71[6] = IN1[15]&IN2[56];
  assign P72[5] = IN1[15]&IN2[57];
  assign P73[4] = IN1[15]&IN2[58];
  assign P74[3] = IN1[15]&IN2[59];
  assign P75[2] = IN1[15]&IN2[60];
  assign P76[1] = IN1[15]&IN2[61];
  assign P77[0] = IN1[15]&IN2[62];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[16] = IN1[16]&IN2[22];
  assign P39[16] = IN1[16]&IN2[23];
  assign P40[16] = IN1[16]&IN2[24];
  assign P41[16] = IN1[16]&IN2[25];
  assign P42[16] = IN1[16]&IN2[26];
  assign P43[16] = IN1[16]&IN2[27];
  assign P44[16] = IN1[16]&IN2[28];
  assign P45[16] = IN1[16]&IN2[29];
  assign P46[16] = IN1[16]&IN2[30];
  assign P47[16] = IN1[16]&IN2[31];
  assign P48[16] = IN1[16]&IN2[32];
  assign P49[16] = IN1[16]&IN2[33];
  assign P50[16] = IN1[16]&IN2[34];
  assign P51[16] = IN1[16]&IN2[35];
  assign P52[16] = IN1[16]&IN2[36];
  assign P53[16] = IN1[16]&IN2[37];
  assign P54[16] = IN1[16]&IN2[38];
  assign P55[16] = IN1[16]&IN2[39];
  assign P56[16] = IN1[16]&IN2[40];
  assign P57[16] = IN1[16]&IN2[41];
  assign P58[16] = IN1[16]&IN2[42];
  assign P59[16] = IN1[16]&IN2[43];
  assign P60[16] = IN1[16]&IN2[44];
  assign P61[16] = IN1[16]&IN2[45];
  assign P62[16] = IN1[16]&IN2[46];
  assign P63[15] = IN1[16]&IN2[47];
  assign P64[14] = IN1[16]&IN2[48];
  assign P65[13] = IN1[16]&IN2[49];
  assign P66[12] = IN1[16]&IN2[50];
  assign P67[11] = IN1[16]&IN2[51];
  assign P68[10] = IN1[16]&IN2[52];
  assign P69[9] = IN1[16]&IN2[53];
  assign P70[8] = IN1[16]&IN2[54];
  assign P71[7] = IN1[16]&IN2[55];
  assign P72[6] = IN1[16]&IN2[56];
  assign P73[5] = IN1[16]&IN2[57];
  assign P74[4] = IN1[16]&IN2[58];
  assign P75[3] = IN1[16]&IN2[59];
  assign P76[2] = IN1[16]&IN2[60];
  assign P77[1] = IN1[16]&IN2[61];
  assign P78[0] = IN1[16]&IN2[62];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[17] = IN1[17]&IN2[21];
  assign P39[17] = IN1[17]&IN2[22];
  assign P40[17] = IN1[17]&IN2[23];
  assign P41[17] = IN1[17]&IN2[24];
  assign P42[17] = IN1[17]&IN2[25];
  assign P43[17] = IN1[17]&IN2[26];
  assign P44[17] = IN1[17]&IN2[27];
  assign P45[17] = IN1[17]&IN2[28];
  assign P46[17] = IN1[17]&IN2[29];
  assign P47[17] = IN1[17]&IN2[30];
  assign P48[17] = IN1[17]&IN2[31];
  assign P49[17] = IN1[17]&IN2[32];
  assign P50[17] = IN1[17]&IN2[33];
  assign P51[17] = IN1[17]&IN2[34];
  assign P52[17] = IN1[17]&IN2[35];
  assign P53[17] = IN1[17]&IN2[36];
  assign P54[17] = IN1[17]&IN2[37];
  assign P55[17] = IN1[17]&IN2[38];
  assign P56[17] = IN1[17]&IN2[39];
  assign P57[17] = IN1[17]&IN2[40];
  assign P58[17] = IN1[17]&IN2[41];
  assign P59[17] = IN1[17]&IN2[42];
  assign P60[17] = IN1[17]&IN2[43];
  assign P61[17] = IN1[17]&IN2[44];
  assign P62[17] = IN1[17]&IN2[45];
  assign P63[16] = IN1[17]&IN2[46];
  assign P64[15] = IN1[17]&IN2[47];
  assign P65[14] = IN1[17]&IN2[48];
  assign P66[13] = IN1[17]&IN2[49];
  assign P67[12] = IN1[17]&IN2[50];
  assign P68[11] = IN1[17]&IN2[51];
  assign P69[10] = IN1[17]&IN2[52];
  assign P70[9] = IN1[17]&IN2[53];
  assign P71[8] = IN1[17]&IN2[54];
  assign P72[7] = IN1[17]&IN2[55];
  assign P73[6] = IN1[17]&IN2[56];
  assign P74[5] = IN1[17]&IN2[57];
  assign P75[4] = IN1[17]&IN2[58];
  assign P76[3] = IN1[17]&IN2[59];
  assign P77[2] = IN1[17]&IN2[60];
  assign P78[1] = IN1[17]&IN2[61];
  assign P79[0] = IN1[17]&IN2[62];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[18] = IN1[18]&IN2[20];
  assign P39[18] = IN1[18]&IN2[21];
  assign P40[18] = IN1[18]&IN2[22];
  assign P41[18] = IN1[18]&IN2[23];
  assign P42[18] = IN1[18]&IN2[24];
  assign P43[18] = IN1[18]&IN2[25];
  assign P44[18] = IN1[18]&IN2[26];
  assign P45[18] = IN1[18]&IN2[27];
  assign P46[18] = IN1[18]&IN2[28];
  assign P47[18] = IN1[18]&IN2[29];
  assign P48[18] = IN1[18]&IN2[30];
  assign P49[18] = IN1[18]&IN2[31];
  assign P50[18] = IN1[18]&IN2[32];
  assign P51[18] = IN1[18]&IN2[33];
  assign P52[18] = IN1[18]&IN2[34];
  assign P53[18] = IN1[18]&IN2[35];
  assign P54[18] = IN1[18]&IN2[36];
  assign P55[18] = IN1[18]&IN2[37];
  assign P56[18] = IN1[18]&IN2[38];
  assign P57[18] = IN1[18]&IN2[39];
  assign P58[18] = IN1[18]&IN2[40];
  assign P59[18] = IN1[18]&IN2[41];
  assign P60[18] = IN1[18]&IN2[42];
  assign P61[18] = IN1[18]&IN2[43];
  assign P62[18] = IN1[18]&IN2[44];
  assign P63[17] = IN1[18]&IN2[45];
  assign P64[16] = IN1[18]&IN2[46];
  assign P65[15] = IN1[18]&IN2[47];
  assign P66[14] = IN1[18]&IN2[48];
  assign P67[13] = IN1[18]&IN2[49];
  assign P68[12] = IN1[18]&IN2[50];
  assign P69[11] = IN1[18]&IN2[51];
  assign P70[10] = IN1[18]&IN2[52];
  assign P71[9] = IN1[18]&IN2[53];
  assign P72[8] = IN1[18]&IN2[54];
  assign P73[7] = IN1[18]&IN2[55];
  assign P74[6] = IN1[18]&IN2[56];
  assign P75[5] = IN1[18]&IN2[57];
  assign P76[4] = IN1[18]&IN2[58];
  assign P77[3] = IN1[18]&IN2[59];
  assign P78[2] = IN1[18]&IN2[60];
  assign P79[1] = IN1[18]&IN2[61];
  assign P80[0] = IN1[18]&IN2[62];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[19] = IN1[19]&IN2[19];
  assign P39[19] = IN1[19]&IN2[20];
  assign P40[19] = IN1[19]&IN2[21];
  assign P41[19] = IN1[19]&IN2[22];
  assign P42[19] = IN1[19]&IN2[23];
  assign P43[19] = IN1[19]&IN2[24];
  assign P44[19] = IN1[19]&IN2[25];
  assign P45[19] = IN1[19]&IN2[26];
  assign P46[19] = IN1[19]&IN2[27];
  assign P47[19] = IN1[19]&IN2[28];
  assign P48[19] = IN1[19]&IN2[29];
  assign P49[19] = IN1[19]&IN2[30];
  assign P50[19] = IN1[19]&IN2[31];
  assign P51[19] = IN1[19]&IN2[32];
  assign P52[19] = IN1[19]&IN2[33];
  assign P53[19] = IN1[19]&IN2[34];
  assign P54[19] = IN1[19]&IN2[35];
  assign P55[19] = IN1[19]&IN2[36];
  assign P56[19] = IN1[19]&IN2[37];
  assign P57[19] = IN1[19]&IN2[38];
  assign P58[19] = IN1[19]&IN2[39];
  assign P59[19] = IN1[19]&IN2[40];
  assign P60[19] = IN1[19]&IN2[41];
  assign P61[19] = IN1[19]&IN2[42];
  assign P62[19] = IN1[19]&IN2[43];
  assign P63[18] = IN1[19]&IN2[44];
  assign P64[17] = IN1[19]&IN2[45];
  assign P65[16] = IN1[19]&IN2[46];
  assign P66[15] = IN1[19]&IN2[47];
  assign P67[14] = IN1[19]&IN2[48];
  assign P68[13] = IN1[19]&IN2[49];
  assign P69[12] = IN1[19]&IN2[50];
  assign P70[11] = IN1[19]&IN2[51];
  assign P71[10] = IN1[19]&IN2[52];
  assign P72[9] = IN1[19]&IN2[53];
  assign P73[8] = IN1[19]&IN2[54];
  assign P74[7] = IN1[19]&IN2[55];
  assign P75[6] = IN1[19]&IN2[56];
  assign P76[5] = IN1[19]&IN2[57];
  assign P77[4] = IN1[19]&IN2[58];
  assign P78[3] = IN1[19]&IN2[59];
  assign P79[2] = IN1[19]&IN2[60];
  assign P80[1] = IN1[19]&IN2[61];
  assign P81[0] = IN1[19]&IN2[62];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[20] = IN1[20]&IN2[18];
  assign P39[20] = IN1[20]&IN2[19];
  assign P40[20] = IN1[20]&IN2[20];
  assign P41[20] = IN1[20]&IN2[21];
  assign P42[20] = IN1[20]&IN2[22];
  assign P43[20] = IN1[20]&IN2[23];
  assign P44[20] = IN1[20]&IN2[24];
  assign P45[20] = IN1[20]&IN2[25];
  assign P46[20] = IN1[20]&IN2[26];
  assign P47[20] = IN1[20]&IN2[27];
  assign P48[20] = IN1[20]&IN2[28];
  assign P49[20] = IN1[20]&IN2[29];
  assign P50[20] = IN1[20]&IN2[30];
  assign P51[20] = IN1[20]&IN2[31];
  assign P52[20] = IN1[20]&IN2[32];
  assign P53[20] = IN1[20]&IN2[33];
  assign P54[20] = IN1[20]&IN2[34];
  assign P55[20] = IN1[20]&IN2[35];
  assign P56[20] = IN1[20]&IN2[36];
  assign P57[20] = IN1[20]&IN2[37];
  assign P58[20] = IN1[20]&IN2[38];
  assign P59[20] = IN1[20]&IN2[39];
  assign P60[20] = IN1[20]&IN2[40];
  assign P61[20] = IN1[20]&IN2[41];
  assign P62[20] = IN1[20]&IN2[42];
  assign P63[19] = IN1[20]&IN2[43];
  assign P64[18] = IN1[20]&IN2[44];
  assign P65[17] = IN1[20]&IN2[45];
  assign P66[16] = IN1[20]&IN2[46];
  assign P67[15] = IN1[20]&IN2[47];
  assign P68[14] = IN1[20]&IN2[48];
  assign P69[13] = IN1[20]&IN2[49];
  assign P70[12] = IN1[20]&IN2[50];
  assign P71[11] = IN1[20]&IN2[51];
  assign P72[10] = IN1[20]&IN2[52];
  assign P73[9] = IN1[20]&IN2[53];
  assign P74[8] = IN1[20]&IN2[54];
  assign P75[7] = IN1[20]&IN2[55];
  assign P76[6] = IN1[20]&IN2[56];
  assign P77[5] = IN1[20]&IN2[57];
  assign P78[4] = IN1[20]&IN2[58];
  assign P79[3] = IN1[20]&IN2[59];
  assign P80[2] = IN1[20]&IN2[60];
  assign P81[1] = IN1[20]&IN2[61];
  assign P82[0] = IN1[20]&IN2[62];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[21] = IN1[21]&IN2[14];
  assign P36[21] = IN1[21]&IN2[15];
  assign P37[21] = IN1[21]&IN2[16];
  assign P38[21] = IN1[21]&IN2[17];
  assign P39[21] = IN1[21]&IN2[18];
  assign P40[21] = IN1[21]&IN2[19];
  assign P41[21] = IN1[21]&IN2[20];
  assign P42[21] = IN1[21]&IN2[21];
  assign P43[21] = IN1[21]&IN2[22];
  assign P44[21] = IN1[21]&IN2[23];
  assign P45[21] = IN1[21]&IN2[24];
  assign P46[21] = IN1[21]&IN2[25];
  assign P47[21] = IN1[21]&IN2[26];
  assign P48[21] = IN1[21]&IN2[27];
  assign P49[21] = IN1[21]&IN2[28];
  assign P50[21] = IN1[21]&IN2[29];
  assign P51[21] = IN1[21]&IN2[30];
  assign P52[21] = IN1[21]&IN2[31];
  assign P53[21] = IN1[21]&IN2[32];
  assign P54[21] = IN1[21]&IN2[33];
  assign P55[21] = IN1[21]&IN2[34];
  assign P56[21] = IN1[21]&IN2[35];
  assign P57[21] = IN1[21]&IN2[36];
  assign P58[21] = IN1[21]&IN2[37];
  assign P59[21] = IN1[21]&IN2[38];
  assign P60[21] = IN1[21]&IN2[39];
  assign P61[21] = IN1[21]&IN2[40];
  assign P62[21] = IN1[21]&IN2[41];
  assign P63[20] = IN1[21]&IN2[42];
  assign P64[19] = IN1[21]&IN2[43];
  assign P65[18] = IN1[21]&IN2[44];
  assign P66[17] = IN1[21]&IN2[45];
  assign P67[16] = IN1[21]&IN2[46];
  assign P68[15] = IN1[21]&IN2[47];
  assign P69[14] = IN1[21]&IN2[48];
  assign P70[13] = IN1[21]&IN2[49];
  assign P71[12] = IN1[21]&IN2[50];
  assign P72[11] = IN1[21]&IN2[51];
  assign P73[10] = IN1[21]&IN2[52];
  assign P74[9] = IN1[21]&IN2[53];
  assign P75[8] = IN1[21]&IN2[54];
  assign P76[7] = IN1[21]&IN2[55];
  assign P77[6] = IN1[21]&IN2[56];
  assign P78[5] = IN1[21]&IN2[57];
  assign P79[4] = IN1[21]&IN2[58];
  assign P80[3] = IN1[21]&IN2[59];
  assign P81[2] = IN1[21]&IN2[60];
  assign P82[1] = IN1[21]&IN2[61];
  assign P83[0] = IN1[21]&IN2[62];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[22] = IN1[22]&IN2[13];
  assign P36[22] = IN1[22]&IN2[14];
  assign P37[22] = IN1[22]&IN2[15];
  assign P38[22] = IN1[22]&IN2[16];
  assign P39[22] = IN1[22]&IN2[17];
  assign P40[22] = IN1[22]&IN2[18];
  assign P41[22] = IN1[22]&IN2[19];
  assign P42[22] = IN1[22]&IN2[20];
  assign P43[22] = IN1[22]&IN2[21];
  assign P44[22] = IN1[22]&IN2[22];
  assign P45[22] = IN1[22]&IN2[23];
  assign P46[22] = IN1[22]&IN2[24];
  assign P47[22] = IN1[22]&IN2[25];
  assign P48[22] = IN1[22]&IN2[26];
  assign P49[22] = IN1[22]&IN2[27];
  assign P50[22] = IN1[22]&IN2[28];
  assign P51[22] = IN1[22]&IN2[29];
  assign P52[22] = IN1[22]&IN2[30];
  assign P53[22] = IN1[22]&IN2[31];
  assign P54[22] = IN1[22]&IN2[32];
  assign P55[22] = IN1[22]&IN2[33];
  assign P56[22] = IN1[22]&IN2[34];
  assign P57[22] = IN1[22]&IN2[35];
  assign P58[22] = IN1[22]&IN2[36];
  assign P59[22] = IN1[22]&IN2[37];
  assign P60[22] = IN1[22]&IN2[38];
  assign P61[22] = IN1[22]&IN2[39];
  assign P62[22] = IN1[22]&IN2[40];
  assign P63[21] = IN1[22]&IN2[41];
  assign P64[20] = IN1[22]&IN2[42];
  assign P65[19] = IN1[22]&IN2[43];
  assign P66[18] = IN1[22]&IN2[44];
  assign P67[17] = IN1[22]&IN2[45];
  assign P68[16] = IN1[22]&IN2[46];
  assign P69[15] = IN1[22]&IN2[47];
  assign P70[14] = IN1[22]&IN2[48];
  assign P71[13] = IN1[22]&IN2[49];
  assign P72[12] = IN1[22]&IN2[50];
  assign P73[11] = IN1[22]&IN2[51];
  assign P74[10] = IN1[22]&IN2[52];
  assign P75[9] = IN1[22]&IN2[53];
  assign P76[8] = IN1[22]&IN2[54];
  assign P77[7] = IN1[22]&IN2[55];
  assign P78[6] = IN1[22]&IN2[56];
  assign P79[5] = IN1[22]&IN2[57];
  assign P80[4] = IN1[22]&IN2[58];
  assign P81[3] = IN1[22]&IN2[59];
  assign P82[2] = IN1[22]&IN2[60];
  assign P83[1] = IN1[22]&IN2[61];
  assign P84[0] = IN1[22]&IN2[62];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[23] = IN1[23]&IN2[12];
  assign P36[23] = IN1[23]&IN2[13];
  assign P37[23] = IN1[23]&IN2[14];
  assign P38[23] = IN1[23]&IN2[15];
  assign P39[23] = IN1[23]&IN2[16];
  assign P40[23] = IN1[23]&IN2[17];
  assign P41[23] = IN1[23]&IN2[18];
  assign P42[23] = IN1[23]&IN2[19];
  assign P43[23] = IN1[23]&IN2[20];
  assign P44[23] = IN1[23]&IN2[21];
  assign P45[23] = IN1[23]&IN2[22];
  assign P46[23] = IN1[23]&IN2[23];
  assign P47[23] = IN1[23]&IN2[24];
  assign P48[23] = IN1[23]&IN2[25];
  assign P49[23] = IN1[23]&IN2[26];
  assign P50[23] = IN1[23]&IN2[27];
  assign P51[23] = IN1[23]&IN2[28];
  assign P52[23] = IN1[23]&IN2[29];
  assign P53[23] = IN1[23]&IN2[30];
  assign P54[23] = IN1[23]&IN2[31];
  assign P55[23] = IN1[23]&IN2[32];
  assign P56[23] = IN1[23]&IN2[33];
  assign P57[23] = IN1[23]&IN2[34];
  assign P58[23] = IN1[23]&IN2[35];
  assign P59[23] = IN1[23]&IN2[36];
  assign P60[23] = IN1[23]&IN2[37];
  assign P61[23] = IN1[23]&IN2[38];
  assign P62[23] = IN1[23]&IN2[39];
  assign P63[22] = IN1[23]&IN2[40];
  assign P64[21] = IN1[23]&IN2[41];
  assign P65[20] = IN1[23]&IN2[42];
  assign P66[19] = IN1[23]&IN2[43];
  assign P67[18] = IN1[23]&IN2[44];
  assign P68[17] = IN1[23]&IN2[45];
  assign P69[16] = IN1[23]&IN2[46];
  assign P70[15] = IN1[23]&IN2[47];
  assign P71[14] = IN1[23]&IN2[48];
  assign P72[13] = IN1[23]&IN2[49];
  assign P73[12] = IN1[23]&IN2[50];
  assign P74[11] = IN1[23]&IN2[51];
  assign P75[10] = IN1[23]&IN2[52];
  assign P76[9] = IN1[23]&IN2[53];
  assign P77[8] = IN1[23]&IN2[54];
  assign P78[7] = IN1[23]&IN2[55];
  assign P79[6] = IN1[23]&IN2[56];
  assign P80[5] = IN1[23]&IN2[57];
  assign P81[4] = IN1[23]&IN2[58];
  assign P82[3] = IN1[23]&IN2[59];
  assign P83[2] = IN1[23]&IN2[60];
  assign P84[1] = IN1[23]&IN2[61];
  assign P85[0] = IN1[23]&IN2[62];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[24] = IN1[24]&IN2[11];
  assign P36[24] = IN1[24]&IN2[12];
  assign P37[24] = IN1[24]&IN2[13];
  assign P38[24] = IN1[24]&IN2[14];
  assign P39[24] = IN1[24]&IN2[15];
  assign P40[24] = IN1[24]&IN2[16];
  assign P41[24] = IN1[24]&IN2[17];
  assign P42[24] = IN1[24]&IN2[18];
  assign P43[24] = IN1[24]&IN2[19];
  assign P44[24] = IN1[24]&IN2[20];
  assign P45[24] = IN1[24]&IN2[21];
  assign P46[24] = IN1[24]&IN2[22];
  assign P47[24] = IN1[24]&IN2[23];
  assign P48[24] = IN1[24]&IN2[24];
  assign P49[24] = IN1[24]&IN2[25];
  assign P50[24] = IN1[24]&IN2[26];
  assign P51[24] = IN1[24]&IN2[27];
  assign P52[24] = IN1[24]&IN2[28];
  assign P53[24] = IN1[24]&IN2[29];
  assign P54[24] = IN1[24]&IN2[30];
  assign P55[24] = IN1[24]&IN2[31];
  assign P56[24] = IN1[24]&IN2[32];
  assign P57[24] = IN1[24]&IN2[33];
  assign P58[24] = IN1[24]&IN2[34];
  assign P59[24] = IN1[24]&IN2[35];
  assign P60[24] = IN1[24]&IN2[36];
  assign P61[24] = IN1[24]&IN2[37];
  assign P62[24] = IN1[24]&IN2[38];
  assign P63[23] = IN1[24]&IN2[39];
  assign P64[22] = IN1[24]&IN2[40];
  assign P65[21] = IN1[24]&IN2[41];
  assign P66[20] = IN1[24]&IN2[42];
  assign P67[19] = IN1[24]&IN2[43];
  assign P68[18] = IN1[24]&IN2[44];
  assign P69[17] = IN1[24]&IN2[45];
  assign P70[16] = IN1[24]&IN2[46];
  assign P71[15] = IN1[24]&IN2[47];
  assign P72[14] = IN1[24]&IN2[48];
  assign P73[13] = IN1[24]&IN2[49];
  assign P74[12] = IN1[24]&IN2[50];
  assign P75[11] = IN1[24]&IN2[51];
  assign P76[10] = IN1[24]&IN2[52];
  assign P77[9] = IN1[24]&IN2[53];
  assign P78[8] = IN1[24]&IN2[54];
  assign P79[7] = IN1[24]&IN2[55];
  assign P80[6] = IN1[24]&IN2[56];
  assign P81[5] = IN1[24]&IN2[57];
  assign P82[4] = IN1[24]&IN2[58];
  assign P83[3] = IN1[24]&IN2[59];
  assign P84[2] = IN1[24]&IN2[60];
  assign P85[1] = IN1[24]&IN2[61];
  assign P86[0] = IN1[24]&IN2[62];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[25] = IN1[25]&IN2[10];
  assign P36[25] = IN1[25]&IN2[11];
  assign P37[25] = IN1[25]&IN2[12];
  assign P38[25] = IN1[25]&IN2[13];
  assign P39[25] = IN1[25]&IN2[14];
  assign P40[25] = IN1[25]&IN2[15];
  assign P41[25] = IN1[25]&IN2[16];
  assign P42[25] = IN1[25]&IN2[17];
  assign P43[25] = IN1[25]&IN2[18];
  assign P44[25] = IN1[25]&IN2[19];
  assign P45[25] = IN1[25]&IN2[20];
  assign P46[25] = IN1[25]&IN2[21];
  assign P47[25] = IN1[25]&IN2[22];
  assign P48[25] = IN1[25]&IN2[23];
  assign P49[25] = IN1[25]&IN2[24];
  assign P50[25] = IN1[25]&IN2[25];
  assign P51[25] = IN1[25]&IN2[26];
  assign P52[25] = IN1[25]&IN2[27];
  assign P53[25] = IN1[25]&IN2[28];
  assign P54[25] = IN1[25]&IN2[29];
  assign P55[25] = IN1[25]&IN2[30];
  assign P56[25] = IN1[25]&IN2[31];
  assign P57[25] = IN1[25]&IN2[32];
  assign P58[25] = IN1[25]&IN2[33];
  assign P59[25] = IN1[25]&IN2[34];
  assign P60[25] = IN1[25]&IN2[35];
  assign P61[25] = IN1[25]&IN2[36];
  assign P62[25] = IN1[25]&IN2[37];
  assign P63[24] = IN1[25]&IN2[38];
  assign P64[23] = IN1[25]&IN2[39];
  assign P65[22] = IN1[25]&IN2[40];
  assign P66[21] = IN1[25]&IN2[41];
  assign P67[20] = IN1[25]&IN2[42];
  assign P68[19] = IN1[25]&IN2[43];
  assign P69[18] = IN1[25]&IN2[44];
  assign P70[17] = IN1[25]&IN2[45];
  assign P71[16] = IN1[25]&IN2[46];
  assign P72[15] = IN1[25]&IN2[47];
  assign P73[14] = IN1[25]&IN2[48];
  assign P74[13] = IN1[25]&IN2[49];
  assign P75[12] = IN1[25]&IN2[50];
  assign P76[11] = IN1[25]&IN2[51];
  assign P77[10] = IN1[25]&IN2[52];
  assign P78[9] = IN1[25]&IN2[53];
  assign P79[8] = IN1[25]&IN2[54];
  assign P80[7] = IN1[25]&IN2[55];
  assign P81[6] = IN1[25]&IN2[56];
  assign P82[5] = IN1[25]&IN2[57];
  assign P83[4] = IN1[25]&IN2[58];
  assign P84[3] = IN1[25]&IN2[59];
  assign P85[2] = IN1[25]&IN2[60];
  assign P86[1] = IN1[25]&IN2[61];
  assign P87[0] = IN1[25]&IN2[62];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[26] = IN1[26]&IN2[3];
  assign P30[26] = IN1[26]&IN2[4];
  assign P31[26] = IN1[26]&IN2[5];
  assign P32[26] = IN1[26]&IN2[6];
  assign P33[26] = IN1[26]&IN2[7];
  assign P34[26] = IN1[26]&IN2[8];
  assign P35[26] = IN1[26]&IN2[9];
  assign P36[26] = IN1[26]&IN2[10];
  assign P37[26] = IN1[26]&IN2[11];
  assign P38[26] = IN1[26]&IN2[12];
  assign P39[26] = IN1[26]&IN2[13];
  assign P40[26] = IN1[26]&IN2[14];
  assign P41[26] = IN1[26]&IN2[15];
  assign P42[26] = IN1[26]&IN2[16];
  assign P43[26] = IN1[26]&IN2[17];
  assign P44[26] = IN1[26]&IN2[18];
  assign P45[26] = IN1[26]&IN2[19];
  assign P46[26] = IN1[26]&IN2[20];
  assign P47[26] = IN1[26]&IN2[21];
  assign P48[26] = IN1[26]&IN2[22];
  assign P49[26] = IN1[26]&IN2[23];
  assign P50[26] = IN1[26]&IN2[24];
  assign P51[26] = IN1[26]&IN2[25];
  assign P52[26] = IN1[26]&IN2[26];
  assign P53[26] = IN1[26]&IN2[27];
  assign P54[26] = IN1[26]&IN2[28];
  assign P55[26] = IN1[26]&IN2[29];
  assign P56[26] = IN1[26]&IN2[30];
  assign P57[26] = IN1[26]&IN2[31];
  assign P58[26] = IN1[26]&IN2[32];
  assign P59[26] = IN1[26]&IN2[33];
  assign P60[26] = IN1[26]&IN2[34];
  assign P61[26] = IN1[26]&IN2[35];
  assign P62[26] = IN1[26]&IN2[36];
  assign P63[25] = IN1[26]&IN2[37];
  assign P64[24] = IN1[26]&IN2[38];
  assign P65[23] = IN1[26]&IN2[39];
  assign P66[22] = IN1[26]&IN2[40];
  assign P67[21] = IN1[26]&IN2[41];
  assign P68[20] = IN1[26]&IN2[42];
  assign P69[19] = IN1[26]&IN2[43];
  assign P70[18] = IN1[26]&IN2[44];
  assign P71[17] = IN1[26]&IN2[45];
  assign P72[16] = IN1[26]&IN2[46];
  assign P73[15] = IN1[26]&IN2[47];
  assign P74[14] = IN1[26]&IN2[48];
  assign P75[13] = IN1[26]&IN2[49];
  assign P76[12] = IN1[26]&IN2[50];
  assign P77[11] = IN1[26]&IN2[51];
  assign P78[10] = IN1[26]&IN2[52];
  assign P79[9] = IN1[26]&IN2[53];
  assign P80[8] = IN1[26]&IN2[54];
  assign P81[7] = IN1[26]&IN2[55];
  assign P82[6] = IN1[26]&IN2[56];
  assign P83[5] = IN1[26]&IN2[57];
  assign P84[4] = IN1[26]&IN2[58];
  assign P85[3] = IN1[26]&IN2[59];
  assign P86[2] = IN1[26]&IN2[60];
  assign P87[1] = IN1[26]&IN2[61];
  assign P88[0] = IN1[26]&IN2[62];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[27] = IN1[27]&IN2[2];
  assign P30[27] = IN1[27]&IN2[3];
  assign P31[27] = IN1[27]&IN2[4];
  assign P32[27] = IN1[27]&IN2[5];
  assign P33[27] = IN1[27]&IN2[6];
  assign P34[27] = IN1[27]&IN2[7];
  assign P35[27] = IN1[27]&IN2[8];
  assign P36[27] = IN1[27]&IN2[9];
  assign P37[27] = IN1[27]&IN2[10];
  assign P38[27] = IN1[27]&IN2[11];
  assign P39[27] = IN1[27]&IN2[12];
  assign P40[27] = IN1[27]&IN2[13];
  assign P41[27] = IN1[27]&IN2[14];
  assign P42[27] = IN1[27]&IN2[15];
  assign P43[27] = IN1[27]&IN2[16];
  assign P44[27] = IN1[27]&IN2[17];
  assign P45[27] = IN1[27]&IN2[18];
  assign P46[27] = IN1[27]&IN2[19];
  assign P47[27] = IN1[27]&IN2[20];
  assign P48[27] = IN1[27]&IN2[21];
  assign P49[27] = IN1[27]&IN2[22];
  assign P50[27] = IN1[27]&IN2[23];
  assign P51[27] = IN1[27]&IN2[24];
  assign P52[27] = IN1[27]&IN2[25];
  assign P53[27] = IN1[27]&IN2[26];
  assign P54[27] = IN1[27]&IN2[27];
  assign P55[27] = IN1[27]&IN2[28];
  assign P56[27] = IN1[27]&IN2[29];
  assign P57[27] = IN1[27]&IN2[30];
  assign P58[27] = IN1[27]&IN2[31];
  assign P59[27] = IN1[27]&IN2[32];
  assign P60[27] = IN1[27]&IN2[33];
  assign P61[27] = IN1[27]&IN2[34];
  assign P62[27] = IN1[27]&IN2[35];
  assign P63[26] = IN1[27]&IN2[36];
  assign P64[25] = IN1[27]&IN2[37];
  assign P65[24] = IN1[27]&IN2[38];
  assign P66[23] = IN1[27]&IN2[39];
  assign P67[22] = IN1[27]&IN2[40];
  assign P68[21] = IN1[27]&IN2[41];
  assign P69[20] = IN1[27]&IN2[42];
  assign P70[19] = IN1[27]&IN2[43];
  assign P71[18] = IN1[27]&IN2[44];
  assign P72[17] = IN1[27]&IN2[45];
  assign P73[16] = IN1[27]&IN2[46];
  assign P74[15] = IN1[27]&IN2[47];
  assign P75[14] = IN1[27]&IN2[48];
  assign P76[13] = IN1[27]&IN2[49];
  assign P77[12] = IN1[27]&IN2[50];
  assign P78[11] = IN1[27]&IN2[51];
  assign P79[10] = IN1[27]&IN2[52];
  assign P80[9] = IN1[27]&IN2[53];
  assign P81[8] = IN1[27]&IN2[54];
  assign P82[7] = IN1[27]&IN2[55];
  assign P83[6] = IN1[27]&IN2[56];
  assign P84[5] = IN1[27]&IN2[57];
  assign P85[4] = IN1[27]&IN2[58];
  assign P86[3] = IN1[27]&IN2[59];
  assign P87[2] = IN1[27]&IN2[60];
  assign P88[1] = IN1[27]&IN2[61];
  assign P89[0] = IN1[27]&IN2[62];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[28] = IN1[28]&IN2[1];
  assign P30[28] = IN1[28]&IN2[2];
  assign P31[28] = IN1[28]&IN2[3];
  assign P32[28] = IN1[28]&IN2[4];
  assign P33[28] = IN1[28]&IN2[5];
  assign P34[28] = IN1[28]&IN2[6];
  assign P35[28] = IN1[28]&IN2[7];
  assign P36[28] = IN1[28]&IN2[8];
  assign P37[28] = IN1[28]&IN2[9];
  assign P38[28] = IN1[28]&IN2[10];
  assign P39[28] = IN1[28]&IN2[11];
  assign P40[28] = IN1[28]&IN2[12];
  assign P41[28] = IN1[28]&IN2[13];
  assign P42[28] = IN1[28]&IN2[14];
  assign P43[28] = IN1[28]&IN2[15];
  assign P44[28] = IN1[28]&IN2[16];
  assign P45[28] = IN1[28]&IN2[17];
  assign P46[28] = IN1[28]&IN2[18];
  assign P47[28] = IN1[28]&IN2[19];
  assign P48[28] = IN1[28]&IN2[20];
  assign P49[28] = IN1[28]&IN2[21];
  assign P50[28] = IN1[28]&IN2[22];
  assign P51[28] = IN1[28]&IN2[23];
  assign P52[28] = IN1[28]&IN2[24];
  assign P53[28] = IN1[28]&IN2[25];
  assign P54[28] = IN1[28]&IN2[26];
  assign P55[28] = IN1[28]&IN2[27];
  assign P56[28] = IN1[28]&IN2[28];
  assign P57[28] = IN1[28]&IN2[29];
  assign P58[28] = IN1[28]&IN2[30];
  assign P59[28] = IN1[28]&IN2[31];
  assign P60[28] = IN1[28]&IN2[32];
  assign P61[28] = IN1[28]&IN2[33];
  assign P62[28] = IN1[28]&IN2[34];
  assign P63[27] = IN1[28]&IN2[35];
  assign P64[26] = IN1[28]&IN2[36];
  assign P65[25] = IN1[28]&IN2[37];
  assign P66[24] = IN1[28]&IN2[38];
  assign P67[23] = IN1[28]&IN2[39];
  assign P68[22] = IN1[28]&IN2[40];
  assign P69[21] = IN1[28]&IN2[41];
  assign P70[20] = IN1[28]&IN2[42];
  assign P71[19] = IN1[28]&IN2[43];
  assign P72[18] = IN1[28]&IN2[44];
  assign P73[17] = IN1[28]&IN2[45];
  assign P74[16] = IN1[28]&IN2[46];
  assign P75[15] = IN1[28]&IN2[47];
  assign P76[14] = IN1[28]&IN2[48];
  assign P77[13] = IN1[28]&IN2[49];
  assign P78[12] = IN1[28]&IN2[50];
  assign P79[11] = IN1[28]&IN2[51];
  assign P80[10] = IN1[28]&IN2[52];
  assign P81[9] = IN1[28]&IN2[53];
  assign P82[8] = IN1[28]&IN2[54];
  assign P83[7] = IN1[28]&IN2[55];
  assign P84[6] = IN1[28]&IN2[56];
  assign P85[5] = IN1[28]&IN2[57];
  assign P86[4] = IN1[28]&IN2[58];
  assign P87[3] = IN1[28]&IN2[59];
  assign P88[2] = IN1[28]&IN2[60];
  assign P89[1] = IN1[28]&IN2[61];
  assign P90[0] = IN1[28]&IN2[62];
  assign P29[29] = IN1[29]&IN2[0];
  assign P30[29] = IN1[29]&IN2[1];
  assign P31[29] = IN1[29]&IN2[2];
  assign P32[29] = IN1[29]&IN2[3];
  assign P33[29] = IN1[29]&IN2[4];
  assign P34[29] = IN1[29]&IN2[5];
  assign P35[29] = IN1[29]&IN2[6];
  assign P36[29] = IN1[29]&IN2[7];
  assign P37[29] = IN1[29]&IN2[8];
  assign P38[29] = IN1[29]&IN2[9];
  assign P39[29] = IN1[29]&IN2[10];
  assign P40[29] = IN1[29]&IN2[11];
  assign P41[29] = IN1[29]&IN2[12];
  assign P42[29] = IN1[29]&IN2[13];
  assign P43[29] = IN1[29]&IN2[14];
  assign P44[29] = IN1[29]&IN2[15];
  assign P45[29] = IN1[29]&IN2[16];
  assign P46[29] = IN1[29]&IN2[17];
  assign P47[29] = IN1[29]&IN2[18];
  assign P48[29] = IN1[29]&IN2[19];
  assign P49[29] = IN1[29]&IN2[20];
  assign P50[29] = IN1[29]&IN2[21];
  assign P51[29] = IN1[29]&IN2[22];
  assign P52[29] = IN1[29]&IN2[23];
  assign P53[29] = IN1[29]&IN2[24];
  assign P54[29] = IN1[29]&IN2[25];
  assign P55[29] = IN1[29]&IN2[26];
  assign P56[29] = IN1[29]&IN2[27];
  assign P57[29] = IN1[29]&IN2[28];
  assign P58[29] = IN1[29]&IN2[29];
  assign P59[29] = IN1[29]&IN2[30];
  assign P60[29] = IN1[29]&IN2[31];
  assign P61[29] = IN1[29]&IN2[32];
  assign P62[29] = IN1[29]&IN2[33];
  assign P63[28] = IN1[29]&IN2[34];
  assign P64[27] = IN1[29]&IN2[35];
  assign P65[26] = IN1[29]&IN2[36];
  assign P66[25] = IN1[29]&IN2[37];
  assign P67[24] = IN1[29]&IN2[38];
  assign P68[23] = IN1[29]&IN2[39];
  assign P69[22] = IN1[29]&IN2[40];
  assign P70[21] = IN1[29]&IN2[41];
  assign P71[20] = IN1[29]&IN2[42];
  assign P72[19] = IN1[29]&IN2[43];
  assign P73[18] = IN1[29]&IN2[44];
  assign P74[17] = IN1[29]&IN2[45];
  assign P75[16] = IN1[29]&IN2[46];
  assign P76[15] = IN1[29]&IN2[47];
  assign P77[14] = IN1[29]&IN2[48];
  assign P78[13] = IN1[29]&IN2[49];
  assign P79[12] = IN1[29]&IN2[50];
  assign P80[11] = IN1[29]&IN2[51];
  assign P81[10] = IN1[29]&IN2[52];
  assign P82[9] = IN1[29]&IN2[53];
  assign P83[8] = IN1[29]&IN2[54];
  assign P84[7] = IN1[29]&IN2[55];
  assign P85[6] = IN1[29]&IN2[56];
  assign P86[5] = IN1[29]&IN2[57];
  assign P87[4] = IN1[29]&IN2[58];
  assign P88[3] = IN1[29]&IN2[59];
  assign P89[2] = IN1[29]&IN2[60];
  assign P90[1] = IN1[29]&IN2[61];
  assign P91[0] = IN1[29]&IN2[62];
  assign P30[30] = IN1[30]&IN2[0];
  assign P31[30] = IN1[30]&IN2[1];
  assign P32[30] = IN1[30]&IN2[2];
  assign P33[30] = IN1[30]&IN2[3];
  assign P34[30] = IN1[30]&IN2[4];
  assign P35[30] = IN1[30]&IN2[5];
  assign P36[30] = IN1[30]&IN2[6];
  assign P37[30] = IN1[30]&IN2[7];
  assign P38[30] = IN1[30]&IN2[8];
  assign P39[30] = IN1[30]&IN2[9];
  assign P40[30] = IN1[30]&IN2[10];
  assign P41[30] = IN1[30]&IN2[11];
  assign P42[30] = IN1[30]&IN2[12];
  assign P43[30] = IN1[30]&IN2[13];
  assign P44[30] = IN1[30]&IN2[14];
  assign P45[30] = IN1[30]&IN2[15];
  assign P46[30] = IN1[30]&IN2[16];
  assign P47[30] = IN1[30]&IN2[17];
  assign P48[30] = IN1[30]&IN2[18];
  assign P49[30] = IN1[30]&IN2[19];
  assign P50[30] = IN1[30]&IN2[20];
  assign P51[30] = IN1[30]&IN2[21];
  assign P52[30] = IN1[30]&IN2[22];
  assign P53[30] = IN1[30]&IN2[23];
  assign P54[30] = IN1[30]&IN2[24];
  assign P55[30] = IN1[30]&IN2[25];
  assign P56[30] = IN1[30]&IN2[26];
  assign P57[30] = IN1[30]&IN2[27];
  assign P58[30] = IN1[30]&IN2[28];
  assign P59[30] = IN1[30]&IN2[29];
  assign P60[30] = IN1[30]&IN2[30];
  assign P61[30] = IN1[30]&IN2[31];
  assign P62[30] = IN1[30]&IN2[32];
  assign P63[29] = IN1[30]&IN2[33];
  assign P64[28] = IN1[30]&IN2[34];
  assign P65[27] = IN1[30]&IN2[35];
  assign P66[26] = IN1[30]&IN2[36];
  assign P67[25] = IN1[30]&IN2[37];
  assign P68[24] = IN1[30]&IN2[38];
  assign P69[23] = IN1[30]&IN2[39];
  assign P70[22] = IN1[30]&IN2[40];
  assign P71[21] = IN1[30]&IN2[41];
  assign P72[20] = IN1[30]&IN2[42];
  assign P73[19] = IN1[30]&IN2[43];
  assign P74[18] = IN1[30]&IN2[44];
  assign P75[17] = IN1[30]&IN2[45];
  assign P76[16] = IN1[30]&IN2[46];
  assign P77[15] = IN1[30]&IN2[47];
  assign P78[14] = IN1[30]&IN2[48];
  assign P79[13] = IN1[30]&IN2[49];
  assign P80[12] = IN1[30]&IN2[50];
  assign P81[11] = IN1[30]&IN2[51];
  assign P82[10] = IN1[30]&IN2[52];
  assign P83[9] = IN1[30]&IN2[53];
  assign P84[8] = IN1[30]&IN2[54];
  assign P85[7] = IN1[30]&IN2[55];
  assign P86[6] = IN1[30]&IN2[56];
  assign P87[5] = IN1[30]&IN2[57];
  assign P88[4] = IN1[30]&IN2[58];
  assign P89[3] = IN1[30]&IN2[59];
  assign P90[2] = IN1[30]&IN2[60];
  assign P91[1] = IN1[30]&IN2[61];
  assign P92[0] = IN1[30]&IN2[62];
  assign P31[31] = IN1[31]&IN2[0];
  assign P32[31] = IN1[31]&IN2[1];
  assign P33[31] = IN1[31]&IN2[2];
  assign P34[31] = IN1[31]&IN2[3];
  assign P35[31] = IN1[31]&IN2[4];
  assign P36[31] = IN1[31]&IN2[5];
  assign P37[31] = IN1[31]&IN2[6];
  assign P38[31] = IN1[31]&IN2[7];
  assign P39[31] = IN1[31]&IN2[8];
  assign P40[31] = IN1[31]&IN2[9];
  assign P41[31] = IN1[31]&IN2[10];
  assign P42[31] = IN1[31]&IN2[11];
  assign P43[31] = IN1[31]&IN2[12];
  assign P44[31] = IN1[31]&IN2[13];
  assign P45[31] = IN1[31]&IN2[14];
  assign P46[31] = IN1[31]&IN2[15];
  assign P47[31] = IN1[31]&IN2[16];
  assign P48[31] = IN1[31]&IN2[17];
  assign P49[31] = IN1[31]&IN2[18];
  assign P50[31] = IN1[31]&IN2[19];
  assign P51[31] = IN1[31]&IN2[20];
  assign P52[31] = IN1[31]&IN2[21];
  assign P53[31] = IN1[31]&IN2[22];
  assign P54[31] = IN1[31]&IN2[23];
  assign P55[31] = IN1[31]&IN2[24];
  assign P56[31] = IN1[31]&IN2[25];
  assign P57[31] = IN1[31]&IN2[26];
  assign P58[31] = IN1[31]&IN2[27];
  assign P59[31] = IN1[31]&IN2[28];
  assign P60[31] = IN1[31]&IN2[29];
  assign P61[31] = IN1[31]&IN2[30];
  assign P62[31] = IN1[31]&IN2[31];
  assign P63[30] = IN1[31]&IN2[32];
  assign P64[29] = IN1[31]&IN2[33];
  assign P65[28] = IN1[31]&IN2[34];
  assign P66[27] = IN1[31]&IN2[35];
  assign P67[26] = IN1[31]&IN2[36];
  assign P68[25] = IN1[31]&IN2[37];
  assign P69[24] = IN1[31]&IN2[38];
  assign P70[23] = IN1[31]&IN2[39];
  assign P71[22] = IN1[31]&IN2[40];
  assign P72[21] = IN1[31]&IN2[41];
  assign P73[20] = IN1[31]&IN2[42];
  assign P74[19] = IN1[31]&IN2[43];
  assign P75[18] = IN1[31]&IN2[44];
  assign P76[17] = IN1[31]&IN2[45];
  assign P77[16] = IN1[31]&IN2[46];
  assign P78[15] = IN1[31]&IN2[47];
  assign P79[14] = IN1[31]&IN2[48];
  assign P80[13] = IN1[31]&IN2[49];
  assign P81[12] = IN1[31]&IN2[50];
  assign P82[11] = IN1[31]&IN2[51];
  assign P83[10] = IN1[31]&IN2[52];
  assign P84[9] = IN1[31]&IN2[53];
  assign P85[8] = IN1[31]&IN2[54];
  assign P86[7] = IN1[31]&IN2[55];
  assign P87[6] = IN1[31]&IN2[56];
  assign P88[5] = IN1[31]&IN2[57];
  assign P89[4] = IN1[31]&IN2[58];
  assign P90[3] = IN1[31]&IN2[59];
  assign P91[2] = IN1[31]&IN2[60];
  assign P92[1] = IN1[31]&IN2[61];
  assign P93[0] = IN1[31]&IN2[62];
  assign P32[32] = IN1[32]&IN2[0];
  assign P33[32] = IN1[32]&IN2[1];
  assign P34[32] = IN1[32]&IN2[2];
  assign P35[32] = IN1[32]&IN2[3];
  assign P36[32] = IN1[32]&IN2[4];
  assign P37[32] = IN1[32]&IN2[5];
  assign P38[32] = IN1[32]&IN2[6];
  assign P39[32] = IN1[32]&IN2[7];
  assign P40[32] = IN1[32]&IN2[8];
  assign P41[32] = IN1[32]&IN2[9];
  assign P42[32] = IN1[32]&IN2[10];
  assign P43[32] = IN1[32]&IN2[11];
  assign P44[32] = IN1[32]&IN2[12];
  assign P45[32] = IN1[32]&IN2[13];
  assign P46[32] = IN1[32]&IN2[14];
  assign P47[32] = IN1[32]&IN2[15];
  assign P48[32] = IN1[32]&IN2[16];
  assign P49[32] = IN1[32]&IN2[17];
  assign P50[32] = IN1[32]&IN2[18];
  assign P51[32] = IN1[32]&IN2[19];
  assign P52[32] = IN1[32]&IN2[20];
  assign P53[32] = IN1[32]&IN2[21];
  assign P54[32] = IN1[32]&IN2[22];
  assign P55[32] = IN1[32]&IN2[23];
  assign P56[32] = IN1[32]&IN2[24];
  assign P57[32] = IN1[32]&IN2[25];
  assign P58[32] = IN1[32]&IN2[26];
  assign P59[32] = IN1[32]&IN2[27];
  assign P60[32] = IN1[32]&IN2[28];
  assign P61[32] = IN1[32]&IN2[29];
  assign P62[32] = IN1[32]&IN2[30];
  assign P63[31] = IN1[32]&IN2[31];
  assign P64[30] = IN1[32]&IN2[32];
  assign P65[29] = IN1[32]&IN2[33];
  assign P66[28] = IN1[32]&IN2[34];
  assign P67[27] = IN1[32]&IN2[35];
  assign P68[26] = IN1[32]&IN2[36];
  assign P69[25] = IN1[32]&IN2[37];
  assign P70[24] = IN1[32]&IN2[38];
  assign P71[23] = IN1[32]&IN2[39];
  assign P72[22] = IN1[32]&IN2[40];
  assign P73[21] = IN1[32]&IN2[41];
  assign P74[20] = IN1[32]&IN2[42];
  assign P75[19] = IN1[32]&IN2[43];
  assign P76[18] = IN1[32]&IN2[44];
  assign P77[17] = IN1[32]&IN2[45];
  assign P78[16] = IN1[32]&IN2[46];
  assign P79[15] = IN1[32]&IN2[47];
  assign P80[14] = IN1[32]&IN2[48];
  assign P81[13] = IN1[32]&IN2[49];
  assign P82[12] = IN1[32]&IN2[50];
  assign P83[11] = IN1[32]&IN2[51];
  assign P84[10] = IN1[32]&IN2[52];
  assign P85[9] = IN1[32]&IN2[53];
  assign P86[8] = IN1[32]&IN2[54];
  assign P87[7] = IN1[32]&IN2[55];
  assign P88[6] = IN1[32]&IN2[56];
  assign P89[5] = IN1[32]&IN2[57];
  assign P90[4] = IN1[32]&IN2[58];
  assign P91[3] = IN1[32]&IN2[59];
  assign P92[2] = IN1[32]&IN2[60];
  assign P93[1] = IN1[32]&IN2[61];
  assign P94[0] = IN1[32]&IN2[62];
  assign P33[33] = IN1[33]&IN2[0];
  assign P34[33] = IN1[33]&IN2[1];
  assign P35[33] = IN1[33]&IN2[2];
  assign P36[33] = IN1[33]&IN2[3];
  assign P37[33] = IN1[33]&IN2[4];
  assign P38[33] = IN1[33]&IN2[5];
  assign P39[33] = IN1[33]&IN2[6];
  assign P40[33] = IN1[33]&IN2[7];
  assign P41[33] = IN1[33]&IN2[8];
  assign P42[33] = IN1[33]&IN2[9];
  assign P43[33] = IN1[33]&IN2[10];
  assign P44[33] = IN1[33]&IN2[11];
  assign P45[33] = IN1[33]&IN2[12];
  assign P46[33] = IN1[33]&IN2[13];
  assign P47[33] = IN1[33]&IN2[14];
  assign P48[33] = IN1[33]&IN2[15];
  assign P49[33] = IN1[33]&IN2[16];
  assign P50[33] = IN1[33]&IN2[17];
  assign P51[33] = IN1[33]&IN2[18];
  assign P52[33] = IN1[33]&IN2[19];
  assign P53[33] = IN1[33]&IN2[20];
  assign P54[33] = IN1[33]&IN2[21];
  assign P55[33] = IN1[33]&IN2[22];
  assign P56[33] = IN1[33]&IN2[23];
  assign P57[33] = IN1[33]&IN2[24];
  assign P58[33] = IN1[33]&IN2[25];
  assign P59[33] = IN1[33]&IN2[26];
  assign P60[33] = IN1[33]&IN2[27];
  assign P61[33] = IN1[33]&IN2[28];
  assign P62[33] = IN1[33]&IN2[29];
  assign P63[32] = IN1[33]&IN2[30];
  assign P64[31] = IN1[33]&IN2[31];
  assign P65[30] = IN1[33]&IN2[32];
  assign P66[29] = IN1[33]&IN2[33];
  assign P67[28] = IN1[33]&IN2[34];
  assign P68[27] = IN1[33]&IN2[35];
  assign P69[26] = IN1[33]&IN2[36];
  assign P70[25] = IN1[33]&IN2[37];
  assign P71[24] = IN1[33]&IN2[38];
  assign P72[23] = IN1[33]&IN2[39];
  assign P73[22] = IN1[33]&IN2[40];
  assign P74[21] = IN1[33]&IN2[41];
  assign P75[20] = IN1[33]&IN2[42];
  assign P76[19] = IN1[33]&IN2[43];
  assign P77[18] = IN1[33]&IN2[44];
  assign P78[17] = IN1[33]&IN2[45];
  assign P79[16] = IN1[33]&IN2[46];
  assign P80[15] = IN1[33]&IN2[47];
  assign P81[14] = IN1[33]&IN2[48];
  assign P82[13] = IN1[33]&IN2[49];
  assign P83[12] = IN1[33]&IN2[50];
  assign P84[11] = IN1[33]&IN2[51];
  assign P85[10] = IN1[33]&IN2[52];
  assign P86[9] = IN1[33]&IN2[53];
  assign P87[8] = IN1[33]&IN2[54];
  assign P88[7] = IN1[33]&IN2[55];
  assign P89[6] = IN1[33]&IN2[56];
  assign P90[5] = IN1[33]&IN2[57];
  assign P91[4] = IN1[33]&IN2[58];
  assign P92[3] = IN1[33]&IN2[59];
  assign P93[2] = IN1[33]&IN2[60];
  assign P94[1] = IN1[33]&IN2[61];
  assign P95[0] = IN1[33]&IN2[62];
  assign P34[34] = IN1[34]&IN2[0];
  assign P35[34] = IN1[34]&IN2[1];
  assign P36[34] = IN1[34]&IN2[2];
  assign P37[34] = IN1[34]&IN2[3];
  assign P38[34] = IN1[34]&IN2[4];
  assign P39[34] = IN1[34]&IN2[5];
  assign P40[34] = IN1[34]&IN2[6];
  assign P41[34] = IN1[34]&IN2[7];
  assign P42[34] = IN1[34]&IN2[8];
  assign P43[34] = IN1[34]&IN2[9];
  assign P44[34] = IN1[34]&IN2[10];
  assign P45[34] = IN1[34]&IN2[11];
  assign P46[34] = IN1[34]&IN2[12];
  assign P47[34] = IN1[34]&IN2[13];
  assign P48[34] = IN1[34]&IN2[14];
  assign P49[34] = IN1[34]&IN2[15];
  assign P50[34] = IN1[34]&IN2[16];
  assign P51[34] = IN1[34]&IN2[17];
  assign P52[34] = IN1[34]&IN2[18];
  assign P53[34] = IN1[34]&IN2[19];
  assign P54[34] = IN1[34]&IN2[20];
  assign P55[34] = IN1[34]&IN2[21];
  assign P56[34] = IN1[34]&IN2[22];
  assign P57[34] = IN1[34]&IN2[23];
  assign P58[34] = IN1[34]&IN2[24];
  assign P59[34] = IN1[34]&IN2[25];
  assign P60[34] = IN1[34]&IN2[26];
  assign P61[34] = IN1[34]&IN2[27];
  assign P62[34] = IN1[34]&IN2[28];
  assign P63[33] = IN1[34]&IN2[29];
  assign P64[32] = IN1[34]&IN2[30];
  assign P65[31] = IN1[34]&IN2[31];
  assign P66[30] = IN1[34]&IN2[32];
  assign P67[29] = IN1[34]&IN2[33];
  assign P68[28] = IN1[34]&IN2[34];
  assign P69[27] = IN1[34]&IN2[35];
  assign P70[26] = IN1[34]&IN2[36];
  assign P71[25] = IN1[34]&IN2[37];
  assign P72[24] = IN1[34]&IN2[38];
  assign P73[23] = IN1[34]&IN2[39];
  assign P74[22] = IN1[34]&IN2[40];
  assign P75[21] = IN1[34]&IN2[41];
  assign P76[20] = IN1[34]&IN2[42];
  assign P77[19] = IN1[34]&IN2[43];
  assign P78[18] = IN1[34]&IN2[44];
  assign P79[17] = IN1[34]&IN2[45];
  assign P80[16] = IN1[34]&IN2[46];
  assign P81[15] = IN1[34]&IN2[47];
  assign P82[14] = IN1[34]&IN2[48];
  assign P83[13] = IN1[34]&IN2[49];
  assign P84[12] = IN1[34]&IN2[50];
  assign P85[11] = IN1[34]&IN2[51];
  assign P86[10] = IN1[34]&IN2[52];
  assign P87[9] = IN1[34]&IN2[53];
  assign P88[8] = IN1[34]&IN2[54];
  assign P89[7] = IN1[34]&IN2[55];
  assign P90[6] = IN1[34]&IN2[56];
  assign P91[5] = IN1[34]&IN2[57];
  assign P92[4] = IN1[34]&IN2[58];
  assign P93[3] = IN1[34]&IN2[59];
  assign P94[2] = IN1[34]&IN2[60];
  assign P95[1] = IN1[34]&IN2[61];
  assign P96[0] = IN1[34]&IN2[62];
  assign P35[35] = IN1[35]&IN2[0];
  assign P36[35] = IN1[35]&IN2[1];
  assign P37[35] = IN1[35]&IN2[2];
  assign P38[35] = IN1[35]&IN2[3];
  assign P39[35] = IN1[35]&IN2[4];
  assign P40[35] = IN1[35]&IN2[5];
  assign P41[35] = IN1[35]&IN2[6];
  assign P42[35] = IN1[35]&IN2[7];
  assign P43[35] = IN1[35]&IN2[8];
  assign P44[35] = IN1[35]&IN2[9];
  assign P45[35] = IN1[35]&IN2[10];
  assign P46[35] = IN1[35]&IN2[11];
  assign P47[35] = IN1[35]&IN2[12];
  assign P48[35] = IN1[35]&IN2[13];
  assign P49[35] = IN1[35]&IN2[14];
  assign P50[35] = IN1[35]&IN2[15];
  assign P51[35] = IN1[35]&IN2[16];
  assign P52[35] = IN1[35]&IN2[17];
  assign P53[35] = IN1[35]&IN2[18];
  assign P54[35] = IN1[35]&IN2[19];
  assign P55[35] = IN1[35]&IN2[20];
  assign P56[35] = IN1[35]&IN2[21];
  assign P57[35] = IN1[35]&IN2[22];
  assign P58[35] = IN1[35]&IN2[23];
  assign P59[35] = IN1[35]&IN2[24];
  assign P60[35] = IN1[35]&IN2[25];
  assign P61[35] = IN1[35]&IN2[26];
  assign P62[35] = IN1[35]&IN2[27];
  assign P63[34] = IN1[35]&IN2[28];
  assign P64[33] = IN1[35]&IN2[29];
  assign P65[32] = IN1[35]&IN2[30];
  assign P66[31] = IN1[35]&IN2[31];
  assign P67[30] = IN1[35]&IN2[32];
  assign P68[29] = IN1[35]&IN2[33];
  assign P69[28] = IN1[35]&IN2[34];
  assign P70[27] = IN1[35]&IN2[35];
  assign P71[26] = IN1[35]&IN2[36];
  assign P72[25] = IN1[35]&IN2[37];
  assign P73[24] = IN1[35]&IN2[38];
  assign P74[23] = IN1[35]&IN2[39];
  assign P75[22] = IN1[35]&IN2[40];
  assign P76[21] = IN1[35]&IN2[41];
  assign P77[20] = IN1[35]&IN2[42];
  assign P78[19] = IN1[35]&IN2[43];
  assign P79[18] = IN1[35]&IN2[44];
  assign P80[17] = IN1[35]&IN2[45];
  assign P81[16] = IN1[35]&IN2[46];
  assign P82[15] = IN1[35]&IN2[47];
  assign P83[14] = IN1[35]&IN2[48];
  assign P84[13] = IN1[35]&IN2[49];
  assign P85[12] = IN1[35]&IN2[50];
  assign P86[11] = IN1[35]&IN2[51];
  assign P87[10] = IN1[35]&IN2[52];
  assign P88[9] = IN1[35]&IN2[53];
  assign P89[8] = IN1[35]&IN2[54];
  assign P90[7] = IN1[35]&IN2[55];
  assign P91[6] = IN1[35]&IN2[56];
  assign P92[5] = IN1[35]&IN2[57];
  assign P93[4] = IN1[35]&IN2[58];
  assign P94[3] = IN1[35]&IN2[59];
  assign P95[2] = IN1[35]&IN2[60];
  assign P96[1] = IN1[35]&IN2[61];
  assign P97[0] = IN1[35]&IN2[62];
  assign P36[36] = IN1[36]&IN2[0];
  assign P37[36] = IN1[36]&IN2[1];
  assign P38[36] = IN1[36]&IN2[2];
  assign P39[36] = IN1[36]&IN2[3];
  assign P40[36] = IN1[36]&IN2[4];
  assign P41[36] = IN1[36]&IN2[5];
  assign P42[36] = IN1[36]&IN2[6];
  assign P43[36] = IN1[36]&IN2[7];
  assign P44[36] = IN1[36]&IN2[8];
  assign P45[36] = IN1[36]&IN2[9];
  assign P46[36] = IN1[36]&IN2[10];
  assign P47[36] = IN1[36]&IN2[11];
  assign P48[36] = IN1[36]&IN2[12];
  assign P49[36] = IN1[36]&IN2[13];
  assign P50[36] = IN1[36]&IN2[14];
  assign P51[36] = IN1[36]&IN2[15];
  assign P52[36] = IN1[36]&IN2[16];
  assign P53[36] = IN1[36]&IN2[17];
  assign P54[36] = IN1[36]&IN2[18];
  assign P55[36] = IN1[36]&IN2[19];
  assign P56[36] = IN1[36]&IN2[20];
  assign P57[36] = IN1[36]&IN2[21];
  assign P58[36] = IN1[36]&IN2[22];
  assign P59[36] = IN1[36]&IN2[23];
  assign P60[36] = IN1[36]&IN2[24];
  assign P61[36] = IN1[36]&IN2[25];
  assign P62[36] = IN1[36]&IN2[26];
  assign P63[35] = IN1[36]&IN2[27];
  assign P64[34] = IN1[36]&IN2[28];
  assign P65[33] = IN1[36]&IN2[29];
  assign P66[32] = IN1[36]&IN2[30];
  assign P67[31] = IN1[36]&IN2[31];
  assign P68[30] = IN1[36]&IN2[32];
  assign P69[29] = IN1[36]&IN2[33];
  assign P70[28] = IN1[36]&IN2[34];
  assign P71[27] = IN1[36]&IN2[35];
  assign P72[26] = IN1[36]&IN2[36];
  assign P73[25] = IN1[36]&IN2[37];
  assign P74[24] = IN1[36]&IN2[38];
  assign P75[23] = IN1[36]&IN2[39];
  assign P76[22] = IN1[36]&IN2[40];
  assign P77[21] = IN1[36]&IN2[41];
  assign P78[20] = IN1[36]&IN2[42];
  assign P79[19] = IN1[36]&IN2[43];
  assign P80[18] = IN1[36]&IN2[44];
  assign P81[17] = IN1[36]&IN2[45];
  assign P82[16] = IN1[36]&IN2[46];
  assign P83[15] = IN1[36]&IN2[47];
  assign P84[14] = IN1[36]&IN2[48];
  assign P85[13] = IN1[36]&IN2[49];
  assign P86[12] = IN1[36]&IN2[50];
  assign P87[11] = IN1[36]&IN2[51];
  assign P88[10] = IN1[36]&IN2[52];
  assign P89[9] = IN1[36]&IN2[53];
  assign P90[8] = IN1[36]&IN2[54];
  assign P91[7] = IN1[36]&IN2[55];
  assign P92[6] = IN1[36]&IN2[56];
  assign P93[5] = IN1[36]&IN2[57];
  assign P94[4] = IN1[36]&IN2[58];
  assign P95[3] = IN1[36]&IN2[59];
  assign P96[2] = IN1[36]&IN2[60];
  assign P97[1] = IN1[36]&IN2[61];
  assign P98[0] = IN1[36]&IN2[62];
  assign P37[37] = IN1[37]&IN2[0];
  assign P38[37] = IN1[37]&IN2[1];
  assign P39[37] = IN1[37]&IN2[2];
  assign P40[37] = IN1[37]&IN2[3];
  assign P41[37] = IN1[37]&IN2[4];
  assign P42[37] = IN1[37]&IN2[5];
  assign P43[37] = IN1[37]&IN2[6];
  assign P44[37] = IN1[37]&IN2[7];
  assign P45[37] = IN1[37]&IN2[8];
  assign P46[37] = IN1[37]&IN2[9];
  assign P47[37] = IN1[37]&IN2[10];
  assign P48[37] = IN1[37]&IN2[11];
  assign P49[37] = IN1[37]&IN2[12];
  assign P50[37] = IN1[37]&IN2[13];
  assign P51[37] = IN1[37]&IN2[14];
  assign P52[37] = IN1[37]&IN2[15];
  assign P53[37] = IN1[37]&IN2[16];
  assign P54[37] = IN1[37]&IN2[17];
  assign P55[37] = IN1[37]&IN2[18];
  assign P56[37] = IN1[37]&IN2[19];
  assign P57[37] = IN1[37]&IN2[20];
  assign P58[37] = IN1[37]&IN2[21];
  assign P59[37] = IN1[37]&IN2[22];
  assign P60[37] = IN1[37]&IN2[23];
  assign P61[37] = IN1[37]&IN2[24];
  assign P62[37] = IN1[37]&IN2[25];
  assign P63[36] = IN1[37]&IN2[26];
  assign P64[35] = IN1[37]&IN2[27];
  assign P65[34] = IN1[37]&IN2[28];
  assign P66[33] = IN1[37]&IN2[29];
  assign P67[32] = IN1[37]&IN2[30];
  assign P68[31] = IN1[37]&IN2[31];
  assign P69[30] = IN1[37]&IN2[32];
  assign P70[29] = IN1[37]&IN2[33];
  assign P71[28] = IN1[37]&IN2[34];
  assign P72[27] = IN1[37]&IN2[35];
  assign P73[26] = IN1[37]&IN2[36];
  assign P74[25] = IN1[37]&IN2[37];
  assign P75[24] = IN1[37]&IN2[38];
  assign P76[23] = IN1[37]&IN2[39];
  assign P77[22] = IN1[37]&IN2[40];
  assign P78[21] = IN1[37]&IN2[41];
  assign P79[20] = IN1[37]&IN2[42];
  assign P80[19] = IN1[37]&IN2[43];
  assign P81[18] = IN1[37]&IN2[44];
  assign P82[17] = IN1[37]&IN2[45];
  assign P83[16] = IN1[37]&IN2[46];
  assign P84[15] = IN1[37]&IN2[47];
  assign P85[14] = IN1[37]&IN2[48];
  assign P86[13] = IN1[37]&IN2[49];
  assign P87[12] = IN1[37]&IN2[50];
  assign P88[11] = IN1[37]&IN2[51];
  assign P89[10] = IN1[37]&IN2[52];
  assign P90[9] = IN1[37]&IN2[53];
  assign P91[8] = IN1[37]&IN2[54];
  assign P92[7] = IN1[37]&IN2[55];
  assign P93[6] = IN1[37]&IN2[56];
  assign P94[5] = IN1[37]&IN2[57];
  assign P95[4] = IN1[37]&IN2[58];
  assign P96[3] = IN1[37]&IN2[59];
  assign P97[2] = IN1[37]&IN2[60];
  assign P98[1] = IN1[37]&IN2[61];
  assign P99[0] = IN1[37]&IN2[62];
  assign P38[38] = IN1[38]&IN2[0];
  assign P39[38] = IN1[38]&IN2[1];
  assign P40[38] = IN1[38]&IN2[2];
  assign P41[38] = IN1[38]&IN2[3];
  assign P42[38] = IN1[38]&IN2[4];
  assign P43[38] = IN1[38]&IN2[5];
  assign P44[38] = IN1[38]&IN2[6];
  assign P45[38] = IN1[38]&IN2[7];
  assign P46[38] = IN1[38]&IN2[8];
  assign P47[38] = IN1[38]&IN2[9];
  assign P48[38] = IN1[38]&IN2[10];
  assign P49[38] = IN1[38]&IN2[11];
  assign P50[38] = IN1[38]&IN2[12];
  assign P51[38] = IN1[38]&IN2[13];
  assign P52[38] = IN1[38]&IN2[14];
  assign P53[38] = IN1[38]&IN2[15];
  assign P54[38] = IN1[38]&IN2[16];
  assign P55[38] = IN1[38]&IN2[17];
  assign P56[38] = IN1[38]&IN2[18];
  assign P57[38] = IN1[38]&IN2[19];
  assign P58[38] = IN1[38]&IN2[20];
  assign P59[38] = IN1[38]&IN2[21];
  assign P60[38] = IN1[38]&IN2[22];
  assign P61[38] = IN1[38]&IN2[23];
  assign P62[38] = IN1[38]&IN2[24];
  assign P63[37] = IN1[38]&IN2[25];
  assign P64[36] = IN1[38]&IN2[26];
  assign P65[35] = IN1[38]&IN2[27];
  assign P66[34] = IN1[38]&IN2[28];
  assign P67[33] = IN1[38]&IN2[29];
  assign P68[32] = IN1[38]&IN2[30];
  assign P69[31] = IN1[38]&IN2[31];
  assign P70[30] = IN1[38]&IN2[32];
  assign P71[29] = IN1[38]&IN2[33];
  assign P72[28] = IN1[38]&IN2[34];
  assign P73[27] = IN1[38]&IN2[35];
  assign P74[26] = IN1[38]&IN2[36];
  assign P75[25] = IN1[38]&IN2[37];
  assign P76[24] = IN1[38]&IN2[38];
  assign P77[23] = IN1[38]&IN2[39];
  assign P78[22] = IN1[38]&IN2[40];
  assign P79[21] = IN1[38]&IN2[41];
  assign P80[20] = IN1[38]&IN2[42];
  assign P81[19] = IN1[38]&IN2[43];
  assign P82[18] = IN1[38]&IN2[44];
  assign P83[17] = IN1[38]&IN2[45];
  assign P84[16] = IN1[38]&IN2[46];
  assign P85[15] = IN1[38]&IN2[47];
  assign P86[14] = IN1[38]&IN2[48];
  assign P87[13] = IN1[38]&IN2[49];
  assign P88[12] = IN1[38]&IN2[50];
  assign P89[11] = IN1[38]&IN2[51];
  assign P90[10] = IN1[38]&IN2[52];
  assign P91[9] = IN1[38]&IN2[53];
  assign P92[8] = IN1[38]&IN2[54];
  assign P93[7] = IN1[38]&IN2[55];
  assign P94[6] = IN1[38]&IN2[56];
  assign P95[5] = IN1[38]&IN2[57];
  assign P96[4] = IN1[38]&IN2[58];
  assign P97[3] = IN1[38]&IN2[59];
  assign P98[2] = IN1[38]&IN2[60];
  assign P99[1] = IN1[38]&IN2[61];
  assign P100[0] = IN1[38]&IN2[62];
  assign P39[39] = IN1[39]&IN2[0];
  assign P40[39] = IN1[39]&IN2[1];
  assign P41[39] = IN1[39]&IN2[2];
  assign P42[39] = IN1[39]&IN2[3];
  assign P43[39] = IN1[39]&IN2[4];
  assign P44[39] = IN1[39]&IN2[5];
  assign P45[39] = IN1[39]&IN2[6];
  assign P46[39] = IN1[39]&IN2[7];
  assign P47[39] = IN1[39]&IN2[8];
  assign P48[39] = IN1[39]&IN2[9];
  assign P49[39] = IN1[39]&IN2[10];
  assign P50[39] = IN1[39]&IN2[11];
  assign P51[39] = IN1[39]&IN2[12];
  assign P52[39] = IN1[39]&IN2[13];
  assign P53[39] = IN1[39]&IN2[14];
  assign P54[39] = IN1[39]&IN2[15];
  assign P55[39] = IN1[39]&IN2[16];
  assign P56[39] = IN1[39]&IN2[17];
  assign P57[39] = IN1[39]&IN2[18];
  assign P58[39] = IN1[39]&IN2[19];
  assign P59[39] = IN1[39]&IN2[20];
  assign P60[39] = IN1[39]&IN2[21];
  assign P61[39] = IN1[39]&IN2[22];
  assign P62[39] = IN1[39]&IN2[23];
  assign P63[38] = IN1[39]&IN2[24];
  assign P64[37] = IN1[39]&IN2[25];
  assign P65[36] = IN1[39]&IN2[26];
  assign P66[35] = IN1[39]&IN2[27];
  assign P67[34] = IN1[39]&IN2[28];
  assign P68[33] = IN1[39]&IN2[29];
  assign P69[32] = IN1[39]&IN2[30];
  assign P70[31] = IN1[39]&IN2[31];
  assign P71[30] = IN1[39]&IN2[32];
  assign P72[29] = IN1[39]&IN2[33];
  assign P73[28] = IN1[39]&IN2[34];
  assign P74[27] = IN1[39]&IN2[35];
  assign P75[26] = IN1[39]&IN2[36];
  assign P76[25] = IN1[39]&IN2[37];
  assign P77[24] = IN1[39]&IN2[38];
  assign P78[23] = IN1[39]&IN2[39];
  assign P79[22] = IN1[39]&IN2[40];
  assign P80[21] = IN1[39]&IN2[41];
  assign P81[20] = IN1[39]&IN2[42];
  assign P82[19] = IN1[39]&IN2[43];
  assign P83[18] = IN1[39]&IN2[44];
  assign P84[17] = IN1[39]&IN2[45];
  assign P85[16] = IN1[39]&IN2[46];
  assign P86[15] = IN1[39]&IN2[47];
  assign P87[14] = IN1[39]&IN2[48];
  assign P88[13] = IN1[39]&IN2[49];
  assign P89[12] = IN1[39]&IN2[50];
  assign P90[11] = IN1[39]&IN2[51];
  assign P91[10] = IN1[39]&IN2[52];
  assign P92[9] = IN1[39]&IN2[53];
  assign P93[8] = IN1[39]&IN2[54];
  assign P94[7] = IN1[39]&IN2[55];
  assign P95[6] = IN1[39]&IN2[56];
  assign P96[5] = IN1[39]&IN2[57];
  assign P97[4] = IN1[39]&IN2[58];
  assign P98[3] = IN1[39]&IN2[59];
  assign P99[2] = IN1[39]&IN2[60];
  assign P100[1] = IN1[39]&IN2[61];
  assign P101[0] = IN1[39]&IN2[62];
  assign P40[40] = IN1[40]&IN2[0];
  assign P41[40] = IN1[40]&IN2[1];
  assign P42[40] = IN1[40]&IN2[2];
  assign P43[40] = IN1[40]&IN2[3];
  assign P44[40] = IN1[40]&IN2[4];
  assign P45[40] = IN1[40]&IN2[5];
  assign P46[40] = IN1[40]&IN2[6];
  assign P47[40] = IN1[40]&IN2[7];
  assign P48[40] = IN1[40]&IN2[8];
  assign P49[40] = IN1[40]&IN2[9];
  assign P50[40] = IN1[40]&IN2[10];
  assign P51[40] = IN1[40]&IN2[11];
  assign P52[40] = IN1[40]&IN2[12];
  assign P53[40] = IN1[40]&IN2[13];
  assign P54[40] = IN1[40]&IN2[14];
  assign P55[40] = IN1[40]&IN2[15];
  assign P56[40] = IN1[40]&IN2[16];
  assign P57[40] = IN1[40]&IN2[17];
  assign P58[40] = IN1[40]&IN2[18];
  assign P59[40] = IN1[40]&IN2[19];
  assign P60[40] = IN1[40]&IN2[20];
  assign P61[40] = IN1[40]&IN2[21];
  assign P62[40] = IN1[40]&IN2[22];
  assign P63[39] = IN1[40]&IN2[23];
  assign P64[38] = IN1[40]&IN2[24];
  assign P65[37] = IN1[40]&IN2[25];
  assign P66[36] = IN1[40]&IN2[26];
  assign P67[35] = IN1[40]&IN2[27];
  assign P68[34] = IN1[40]&IN2[28];
  assign P69[33] = IN1[40]&IN2[29];
  assign P70[32] = IN1[40]&IN2[30];
  assign P71[31] = IN1[40]&IN2[31];
  assign P72[30] = IN1[40]&IN2[32];
  assign P73[29] = IN1[40]&IN2[33];
  assign P74[28] = IN1[40]&IN2[34];
  assign P75[27] = IN1[40]&IN2[35];
  assign P76[26] = IN1[40]&IN2[36];
  assign P77[25] = IN1[40]&IN2[37];
  assign P78[24] = IN1[40]&IN2[38];
  assign P79[23] = IN1[40]&IN2[39];
  assign P80[22] = IN1[40]&IN2[40];
  assign P81[21] = IN1[40]&IN2[41];
  assign P82[20] = IN1[40]&IN2[42];
  assign P83[19] = IN1[40]&IN2[43];
  assign P84[18] = IN1[40]&IN2[44];
  assign P85[17] = IN1[40]&IN2[45];
  assign P86[16] = IN1[40]&IN2[46];
  assign P87[15] = IN1[40]&IN2[47];
  assign P88[14] = IN1[40]&IN2[48];
  assign P89[13] = IN1[40]&IN2[49];
  assign P90[12] = IN1[40]&IN2[50];
  assign P91[11] = IN1[40]&IN2[51];
  assign P92[10] = IN1[40]&IN2[52];
  assign P93[9] = IN1[40]&IN2[53];
  assign P94[8] = IN1[40]&IN2[54];
  assign P95[7] = IN1[40]&IN2[55];
  assign P96[6] = IN1[40]&IN2[56];
  assign P97[5] = IN1[40]&IN2[57];
  assign P98[4] = IN1[40]&IN2[58];
  assign P99[3] = IN1[40]&IN2[59];
  assign P100[2] = IN1[40]&IN2[60];
  assign P101[1] = IN1[40]&IN2[61];
  assign P102[0] = IN1[40]&IN2[62];
  assign P41[41] = IN1[41]&IN2[0];
  assign P42[41] = IN1[41]&IN2[1];
  assign P43[41] = IN1[41]&IN2[2];
  assign P44[41] = IN1[41]&IN2[3];
  assign P45[41] = IN1[41]&IN2[4];
  assign P46[41] = IN1[41]&IN2[5];
  assign P47[41] = IN1[41]&IN2[6];
  assign P48[41] = IN1[41]&IN2[7];
  assign P49[41] = IN1[41]&IN2[8];
  assign P50[41] = IN1[41]&IN2[9];
  assign P51[41] = IN1[41]&IN2[10];
  assign P52[41] = IN1[41]&IN2[11];
  assign P53[41] = IN1[41]&IN2[12];
  assign P54[41] = IN1[41]&IN2[13];
  assign P55[41] = IN1[41]&IN2[14];
  assign P56[41] = IN1[41]&IN2[15];
  assign P57[41] = IN1[41]&IN2[16];
  assign P58[41] = IN1[41]&IN2[17];
  assign P59[41] = IN1[41]&IN2[18];
  assign P60[41] = IN1[41]&IN2[19];
  assign P61[41] = IN1[41]&IN2[20];
  assign P62[41] = IN1[41]&IN2[21];
  assign P63[40] = IN1[41]&IN2[22];
  assign P64[39] = IN1[41]&IN2[23];
  assign P65[38] = IN1[41]&IN2[24];
  assign P66[37] = IN1[41]&IN2[25];
  assign P67[36] = IN1[41]&IN2[26];
  assign P68[35] = IN1[41]&IN2[27];
  assign P69[34] = IN1[41]&IN2[28];
  assign P70[33] = IN1[41]&IN2[29];
  assign P71[32] = IN1[41]&IN2[30];
  assign P72[31] = IN1[41]&IN2[31];
  assign P73[30] = IN1[41]&IN2[32];
  assign P74[29] = IN1[41]&IN2[33];
  assign P75[28] = IN1[41]&IN2[34];
  assign P76[27] = IN1[41]&IN2[35];
  assign P77[26] = IN1[41]&IN2[36];
  assign P78[25] = IN1[41]&IN2[37];
  assign P79[24] = IN1[41]&IN2[38];
  assign P80[23] = IN1[41]&IN2[39];
  assign P81[22] = IN1[41]&IN2[40];
  assign P82[21] = IN1[41]&IN2[41];
  assign P83[20] = IN1[41]&IN2[42];
  assign P84[19] = IN1[41]&IN2[43];
  assign P85[18] = IN1[41]&IN2[44];
  assign P86[17] = IN1[41]&IN2[45];
  assign P87[16] = IN1[41]&IN2[46];
  assign P88[15] = IN1[41]&IN2[47];
  assign P89[14] = IN1[41]&IN2[48];
  assign P90[13] = IN1[41]&IN2[49];
  assign P91[12] = IN1[41]&IN2[50];
  assign P92[11] = IN1[41]&IN2[51];
  assign P93[10] = IN1[41]&IN2[52];
  assign P94[9] = IN1[41]&IN2[53];
  assign P95[8] = IN1[41]&IN2[54];
  assign P96[7] = IN1[41]&IN2[55];
  assign P97[6] = IN1[41]&IN2[56];
  assign P98[5] = IN1[41]&IN2[57];
  assign P99[4] = IN1[41]&IN2[58];
  assign P100[3] = IN1[41]&IN2[59];
  assign P101[2] = IN1[41]&IN2[60];
  assign P102[1] = IN1[41]&IN2[61];
  assign P103[0] = IN1[41]&IN2[62];
  assign P42[42] = IN1[42]&IN2[0];
  assign P43[42] = IN1[42]&IN2[1];
  assign P44[42] = IN1[42]&IN2[2];
  assign P45[42] = IN1[42]&IN2[3];
  assign P46[42] = IN1[42]&IN2[4];
  assign P47[42] = IN1[42]&IN2[5];
  assign P48[42] = IN1[42]&IN2[6];
  assign P49[42] = IN1[42]&IN2[7];
  assign P50[42] = IN1[42]&IN2[8];
  assign P51[42] = IN1[42]&IN2[9];
  assign P52[42] = IN1[42]&IN2[10];
  assign P53[42] = IN1[42]&IN2[11];
  assign P54[42] = IN1[42]&IN2[12];
  assign P55[42] = IN1[42]&IN2[13];
  assign P56[42] = IN1[42]&IN2[14];
  assign P57[42] = IN1[42]&IN2[15];
  assign P58[42] = IN1[42]&IN2[16];
  assign P59[42] = IN1[42]&IN2[17];
  assign P60[42] = IN1[42]&IN2[18];
  assign P61[42] = IN1[42]&IN2[19];
  assign P62[42] = IN1[42]&IN2[20];
  assign P63[41] = IN1[42]&IN2[21];
  assign P64[40] = IN1[42]&IN2[22];
  assign P65[39] = IN1[42]&IN2[23];
  assign P66[38] = IN1[42]&IN2[24];
  assign P67[37] = IN1[42]&IN2[25];
  assign P68[36] = IN1[42]&IN2[26];
  assign P69[35] = IN1[42]&IN2[27];
  assign P70[34] = IN1[42]&IN2[28];
  assign P71[33] = IN1[42]&IN2[29];
  assign P72[32] = IN1[42]&IN2[30];
  assign P73[31] = IN1[42]&IN2[31];
  assign P74[30] = IN1[42]&IN2[32];
  assign P75[29] = IN1[42]&IN2[33];
  assign P76[28] = IN1[42]&IN2[34];
  assign P77[27] = IN1[42]&IN2[35];
  assign P78[26] = IN1[42]&IN2[36];
  assign P79[25] = IN1[42]&IN2[37];
  assign P80[24] = IN1[42]&IN2[38];
  assign P81[23] = IN1[42]&IN2[39];
  assign P82[22] = IN1[42]&IN2[40];
  assign P83[21] = IN1[42]&IN2[41];
  assign P84[20] = IN1[42]&IN2[42];
  assign P85[19] = IN1[42]&IN2[43];
  assign P86[18] = IN1[42]&IN2[44];
  assign P87[17] = IN1[42]&IN2[45];
  assign P88[16] = IN1[42]&IN2[46];
  assign P89[15] = IN1[42]&IN2[47];
  assign P90[14] = IN1[42]&IN2[48];
  assign P91[13] = IN1[42]&IN2[49];
  assign P92[12] = IN1[42]&IN2[50];
  assign P93[11] = IN1[42]&IN2[51];
  assign P94[10] = IN1[42]&IN2[52];
  assign P95[9] = IN1[42]&IN2[53];
  assign P96[8] = IN1[42]&IN2[54];
  assign P97[7] = IN1[42]&IN2[55];
  assign P98[6] = IN1[42]&IN2[56];
  assign P99[5] = IN1[42]&IN2[57];
  assign P100[4] = IN1[42]&IN2[58];
  assign P101[3] = IN1[42]&IN2[59];
  assign P102[2] = IN1[42]&IN2[60];
  assign P103[1] = IN1[42]&IN2[61];
  assign P104[0] = IN1[42]&IN2[62];
  assign P43[43] = IN1[43]&IN2[0];
  assign P44[43] = IN1[43]&IN2[1];
  assign P45[43] = IN1[43]&IN2[2];
  assign P46[43] = IN1[43]&IN2[3];
  assign P47[43] = IN1[43]&IN2[4];
  assign P48[43] = IN1[43]&IN2[5];
  assign P49[43] = IN1[43]&IN2[6];
  assign P50[43] = IN1[43]&IN2[7];
  assign P51[43] = IN1[43]&IN2[8];
  assign P52[43] = IN1[43]&IN2[9];
  assign P53[43] = IN1[43]&IN2[10];
  assign P54[43] = IN1[43]&IN2[11];
  assign P55[43] = IN1[43]&IN2[12];
  assign P56[43] = IN1[43]&IN2[13];
  assign P57[43] = IN1[43]&IN2[14];
  assign P58[43] = IN1[43]&IN2[15];
  assign P59[43] = IN1[43]&IN2[16];
  assign P60[43] = IN1[43]&IN2[17];
  assign P61[43] = IN1[43]&IN2[18];
  assign P62[43] = IN1[43]&IN2[19];
  assign P63[42] = IN1[43]&IN2[20];
  assign P64[41] = IN1[43]&IN2[21];
  assign P65[40] = IN1[43]&IN2[22];
  assign P66[39] = IN1[43]&IN2[23];
  assign P67[38] = IN1[43]&IN2[24];
  assign P68[37] = IN1[43]&IN2[25];
  assign P69[36] = IN1[43]&IN2[26];
  assign P70[35] = IN1[43]&IN2[27];
  assign P71[34] = IN1[43]&IN2[28];
  assign P72[33] = IN1[43]&IN2[29];
  assign P73[32] = IN1[43]&IN2[30];
  assign P74[31] = IN1[43]&IN2[31];
  assign P75[30] = IN1[43]&IN2[32];
  assign P76[29] = IN1[43]&IN2[33];
  assign P77[28] = IN1[43]&IN2[34];
  assign P78[27] = IN1[43]&IN2[35];
  assign P79[26] = IN1[43]&IN2[36];
  assign P80[25] = IN1[43]&IN2[37];
  assign P81[24] = IN1[43]&IN2[38];
  assign P82[23] = IN1[43]&IN2[39];
  assign P83[22] = IN1[43]&IN2[40];
  assign P84[21] = IN1[43]&IN2[41];
  assign P85[20] = IN1[43]&IN2[42];
  assign P86[19] = IN1[43]&IN2[43];
  assign P87[18] = IN1[43]&IN2[44];
  assign P88[17] = IN1[43]&IN2[45];
  assign P89[16] = IN1[43]&IN2[46];
  assign P90[15] = IN1[43]&IN2[47];
  assign P91[14] = IN1[43]&IN2[48];
  assign P92[13] = IN1[43]&IN2[49];
  assign P93[12] = IN1[43]&IN2[50];
  assign P94[11] = IN1[43]&IN2[51];
  assign P95[10] = IN1[43]&IN2[52];
  assign P96[9] = IN1[43]&IN2[53];
  assign P97[8] = IN1[43]&IN2[54];
  assign P98[7] = IN1[43]&IN2[55];
  assign P99[6] = IN1[43]&IN2[56];
  assign P100[5] = IN1[43]&IN2[57];
  assign P101[4] = IN1[43]&IN2[58];
  assign P102[3] = IN1[43]&IN2[59];
  assign P103[2] = IN1[43]&IN2[60];
  assign P104[1] = IN1[43]&IN2[61];
  assign P105[0] = IN1[43]&IN2[62];
  assign P44[44] = IN1[44]&IN2[0];
  assign P45[44] = IN1[44]&IN2[1];
  assign P46[44] = IN1[44]&IN2[2];
  assign P47[44] = IN1[44]&IN2[3];
  assign P48[44] = IN1[44]&IN2[4];
  assign P49[44] = IN1[44]&IN2[5];
  assign P50[44] = IN1[44]&IN2[6];
  assign P51[44] = IN1[44]&IN2[7];
  assign P52[44] = IN1[44]&IN2[8];
  assign P53[44] = IN1[44]&IN2[9];
  assign P54[44] = IN1[44]&IN2[10];
  assign P55[44] = IN1[44]&IN2[11];
  assign P56[44] = IN1[44]&IN2[12];
  assign P57[44] = IN1[44]&IN2[13];
  assign P58[44] = IN1[44]&IN2[14];
  assign P59[44] = IN1[44]&IN2[15];
  assign P60[44] = IN1[44]&IN2[16];
  assign P61[44] = IN1[44]&IN2[17];
  assign P62[44] = IN1[44]&IN2[18];
  assign P63[43] = IN1[44]&IN2[19];
  assign P64[42] = IN1[44]&IN2[20];
  assign P65[41] = IN1[44]&IN2[21];
  assign P66[40] = IN1[44]&IN2[22];
  assign P67[39] = IN1[44]&IN2[23];
  assign P68[38] = IN1[44]&IN2[24];
  assign P69[37] = IN1[44]&IN2[25];
  assign P70[36] = IN1[44]&IN2[26];
  assign P71[35] = IN1[44]&IN2[27];
  assign P72[34] = IN1[44]&IN2[28];
  assign P73[33] = IN1[44]&IN2[29];
  assign P74[32] = IN1[44]&IN2[30];
  assign P75[31] = IN1[44]&IN2[31];
  assign P76[30] = IN1[44]&IN2[32];
  assign P77[29] = IN1[44]&IN2[33];
  assign P78[28] = IN1[44]&IN2[34];
  assign P79[27] = IN1[44]&IN2[35];
  assign P80[26] = IN1[44]&IN2[36];
  assign P81[25] = IN1[44]&IN2[37];
  assign P82[24] = IN1[44]&IN2[38];
  assign P83[23] = IN1[44]&IN2[39];
  assign P84[22] = IN1[44]&IN2[40];
  assign P85[21] = IN1[44]&IN2[41];
  assign P86[20] = IN1[44]&IN2[42];
  assign P87[19] = IN1[44]&IN2[43];
  assign P88[18] = IN1[44]&IN2[44];
  assign P89[17] = IN1[44]&IN2[45];
  assign P90[16] = IN1[44]&IN2[46];
  assign P91[15] = IN1[44]&IN2[47];
  assign P92[14] = IN1[44]&IN2[48];
  assign P93[13] = IN1[44]&IN2[49];
  assign P94[12] = IN1[44]&IN2[50];
  assign P95[11] = IN1[44]&IN2[51];
  assign P96[10] = IN1[44]&IN2[52];
  assign P97[9] = IN1[44]&IN2[53];
  assign P98[8] = IN1[44]&IN2[54];
  assign P99[7] = IN1[44]&IN2[55];
  assign P100[6] = IN1[44]&IN2[56];
  assign P101[5] = IN1[44]&IN2[57];
  assign P102[4] = IN1[44]&IN2[58];
  assign P103[3] = IN1[44]&IN2[59];
  assign P104[2] = IN1[44]&IN2[60];
  assign P105[1] = IN1[44]&IN2[61];
  assign P106[0] = IN1[44]&IN2[62];
  assign P45[45] = IN1[45]&IN2[0];
  assign P46[45] = IN1[45]&IN2[1];
  assign P47[45] = IN1[45]&IN2[2];
  assign P48[45] = IN1[45]&IN2[3];
  assign P49[45] = IN1[45]&IN2[4];
  assign P50[45] = IN1[45]&IN2[5];
  assign P51[45] = IN1[45]&IN2[6];
  assign P52[45] = IN1[45]&IN2[7];
  assign P53[45] = IN1[45]&IN2[8];
  assign P54[45] = IN1[45]&IN2[9];
  assign P55[45] = IN1[45]&IN2[10];
  assign P56[45] = IN1[45]&IN2[11];
  assign P57[45] = IN1[45]&IN2[12];
  assign P58[45] = IN1[45]&IN2[13];
  assign P59[45] = IN1[45]&IN2[14];
  assign P60[45] = IN1[45]&IN2[15];
  assign P61[45] = IN1[45]&IN2[16];
  assign P62[45] = IN1[45]&IN2[17];
  assign P63[44] = IN1[45]&IN2[18];
  assign P64[43] = IN1[45]&IN2[19];
  assign P65[42] = IN1[45]&IN2[20];
  assign P66[41] = IN1[45]&IN2[21];
  assign P67[40] = IN1[45]&IN2[22];
  assign P68[39] = IN1[45]&IN2[23];
  assign P69[38] = IN1[45]&IN2[24];
  assign P70[37] = IN1[45]&IN2[25];
  assign P71[36] = IN1[45]&IN2[26];
  assign P72[35] = IN1[45]&IN2[27];
  assign P73[34] = IN1[45]&IN2[28];
  assign P74[33] = IN1[45]&IN2[29];
  assign P75[32] = IN1[45]&IN2[30];
  assign P76[31] = IN1[45]&IN2[31];
  assign P77[30] = IN1[45]&IN2[32];
  assign P78[29] = IN1[45]&IN2[33];
  assign P79[28] = IN1[45]&IN2[34];
  assign P80[27] = IN1[45]&IN2[35];
  assign P81[26] = IN1[45]&IN2[36];
  assign P82[25] = IN1[45]&IN2[37];
  assign P83[24] = IN1[45]&IN2[38];
  assign P84[23] = IN1[45]&IN2[39];
  assign P85[22] = IN1[45]&IN2[40];
  assign P86[21] = IN1[45]&IN2[41];
  assign P87[20] = IN1[45]&IN2[42];
  assign P88[19] = IN1[45]&IN2[43];
  assign P89[18] = IN1[45]&IN2[44];
  assign P90[17] = IN1[45]&IN2[45];
  assign P91[16] = IN1[45]&IN2[46];
  assign P92[15] = IN1[45]&IN2[47];
  assign P93[14] = IN1[45]&IN2[48];
  assign P94[13] = IN1[45]&IN2[49];
  assign P95[12] = IN1[45]&IN2[50];
  assign P96[11] = IN1[45]&IN2[51];
  assign P97[10] = IN1[45]&IN2[52];
  assign P98[9] = IN1[45]&IN2[53];
  assign P99[8] = IN1[45]&IN2[54];
  assign P100[7] = IN1[45]&IN2[55];
  assign P101[6] = IN1[45]&IN2[56];
  assign P102[5] = IN1[45]&IN2[57];
  assign P103[4] = IN1[45]&IN2[58];
  assign P104[3] = IN1[45]&IN2[59];
  assign P105[2] = IN1[45]&IN2[60];
  assign P106[1] = IN1[45]&IN2[61];
  assign P107[0] = IN1[45]&IN2[62];
  assign P46[46] = IN1[46]&IN2[0];
  assign P47[46] = IN1[46]&IN2[1];
  assign P48[46] = IN1[46]&IN2[2];
  assign P49[46] = IN1[46]&IN2[3];
  assign P50[46] = IN1[46]&IN2[4];
  assign P51[46] = IN1[46]&IN2[5];
  assign P52[46] = IN1[46]&IN2[6];
  assign P53[46] = IN1[46]&IN2[7];
  assign P54[46] = IN1[46]&IN2[8];
  assign P55[46] = IN1[46]&IN2[9];
  assign P56[46] = IN1[46]&IN2[10];
  assign P57[46] = IN1[46]&IN2[11];
  assign P58[46] = IN1[46]&IN2[12];
  assign P59[46] = IN1[46]&IN2[13];
  assign P60[46] = IN1[46]&IN2[14];
  assign P61[46] = IN1[46]&IN2[15];
  assign P62[46] = IN1[46]&IN2[16];
  assign P63[45] = IN1[46]&IN2[17];
  assign P64[44] = IN1[46]&IN2[18];
  assign P65[43] = IN1[46]&IN2[19];
  assign P66[42] = IN1[46]&IN2[20];
  assign P67[41] = IN1[46]&IN2[21];
  assign P68[40] = IN1[46]&IN2[22];
  assign P69[39] = IN1[46]&IN2[23];
  assign P70[38] = IN1[46]&IN2[24];
  assign P71[37] = IN1[46]&IN2[25];
  assign P72[36] = IN1[46]&IN2[26];
  assign P73[35] = IN1[46]&IN2[27];
  assign P74[34] = IN1[46]&IN2[28];
  assign P75[33] = IN1[46]&IN2[29];
  assign P76[32] = IN1[46]&IN2[30];
  assign P77[31] = IN1[46]&IN2[31];
  assign P78[30] = IN1[46]&IN2[32];
  assign P79[29] = IN1[46]&IN2[33];
  assign P80[28] = IN1[46]&IN2[34];
  assign P81[27] = IN1[46]&IN2[35];
  assign P82[26] = IN1[46]&IN2[36];
  assign P83[25] = IN1[46]&IN2[37];
  assign P84[24] = IN1[46]&IN2[38];
  assign P85[23] = IN1[46]&IN2[39];
  assign P86[22] = IN1[46]&IN2[40];
  assign P87[21] = IN1[46]&IN2[41];
  assign P88[20] = IN1[46]&IN2[42];
  assign P89[19] = IN1[46]&IN2[43];
  assign P90[18] = IN1[46]&IN2[44];
  assign P91[17] = IN1[46]&IN2[45];
  assign P92[16] = IN1[46]&IN2[46];
  assign P93[15] = IN1[46]&IN2[47];
  assign P94[14] = IN1[46]&IN2[48];
  assign P95[13] = IN1[46]&IN2[49];
  assign P96[12] = IN1[46]&IN2[50];
  assign P97[11] = IN1[46]&IN2[51];
  assign P98[10] = IN1[46]&IN2[52];
  assign P99[9] = IN1[46]&IN2[53];
  assign P100[8] = IN1[46]&IN2[54];
  assign P101[7] = IN1[46]&IN2[55];
  assign P102[6] = IN1[46]&IN2[56];
  assign P103[5] = IN1[46]&IN2[57];
  assign P104[4] = IN1[46]&IN2[58];
  assign P105[3] = IN1[46]&IN2[59];
  assign P106[2] = IN1[46]&IN2[60];
  assign P107[1] = IN1[46]&IN2[61];
  assign P108[0] = IN1[46]&IN2[62];
  assign P47[47] = IN1[47]&IN2[0];
  assign P48[47] = IN1[47]&IN2[1];
  assign P49[47] = IN1[47]&IN2[2];
  assign P50[47] = IN1[47]&IN2[3];
  assign P51[47] = IN1[47]&IN2[4];
  assign P52[47] = IN1[47]&IN2[5];
  assign P53[47] = IN1[47]&IN2[6];
  assign P54[47] = IN1[47]&IN2[7];
  assign P55[47] = IN1[47]&IN2[8];
  assign P56[47] = IN1[47]&IN2[9];
  assign P57[47] = IN1[47]&IN2[10];
  assign P58[47] = IN1[47]&IN2[11];
  assign P59[47] = IN1[47]&IN2[12];
  assign P60[47] = IN1[47]&IN2[13];
  assign P61[47] = IN1[47]&IN2[14];
  assign P62[47] = IN1[47]&IN2[15];
  assign P63[46] = IN1[47]&IN2[16];
  assign P64[45] = IN1[47]&IN2[17];
  assign P65[44] = IN1[47]&IN2[18];
  assign P66[43] = IN1[47]&IN2[19];
  assign P67[42] = IN1[47]&IN2[20];
  assign P68[41] = IN1[47]&IN2[21];
  assign P69[40] = IN1[47]&IN2[22];
  assign P70[39] = IN1[47]&IN2[23];
  assign P71[38] = IN1[47]&IN2[24];
  assign P72[37] = IN1[47]&IN2[25];
  assign P73[36] = IN1[47]&IN2[26];
  assign P74[35] = IN1[47]&IN2[27];
  assign P75[34] = IN1[47]&IN2[28];
  assign P76[33] = IN1[47]&IN2[29];
  assign P77[32] = IN1[47]&IN2[30];
  assign P78[31] = IN1[47]&IN2[31];
  assign P79[30] = IN1[47]&IN2[32];
  assign P80[29] = IN1[47]&IN2[33];
  assign P81[28] = IN1[47]&IN2[34];
  assign P82[27] = IN1[47]&IN2[35];
  assign P83[26] = IN1[47]&IN2[36];
  assign P84[25] = IN1[47]&IN2[37];
  assign P85[24] = IN1[47]&IN2[38];
  assign P86[23] = IN1[47]&IN2[39];
  assign P87[22] = IN1[47]&IN2[40];
  assign P88[21] = IN1[47]&IN2[41];
  assign P89[20] = IN1[47]&IN2[42];
  assign P90[19] = IN1[47]&IN2[43];
  assign P91[18] = IN1[47]&IN2[44];
  assign P92[17] = IN1[47]&IN2[45];
  assign P93[16] = IN1[47]&IN2[46];
  assign P94[15] = IN1[47]&IN2[47];
  assign P95[14] = IN1[47]&IN2[48];
  assign P96[13] = IN1[47]&IN2[49];
  assign P97[12] = IN1[47]&IN2[50];
  assign P98[11] = IN1[47]&IN2[51];
  assign P99[10] = IN1[47]&IN2[52];
  assign P100[9] = IN1[47]&IN2[53];
  assign P101[8] = IN1[47]&IN2[54];
  assign P102[7] = IN1[47]&IN2[55];
  assign P103[6] = IN1[47]&IN2[56];
  assign P104[5] = IN1[47]&IN2[57];
  assign P105[4] = IN1[47]&IN2[58];
  assign P106[3] = IN1[47]&IN2[59];
  assign P107[2] = IN1[47]&IN2[60];
  assign P108[1] = IN1[47]&IN2[61];
  assign P109[0] = IN1[47]&IN2[62];
  assign P48[48] = IN1[48]&IN2[0];
  assign P49[48] = IN1[48]&IN2[1];
  assign P50[48] = IN1[48]&IN2[2];
  assign P51[48] = IN1[48]&IN2[3];
  assign P52[48] = IN1[48]&IN2[4];
  assign P53[48] = IN1[48]&IN2[5];
  assign P54[48] = IN1[48]&IN2[6];
  assign P55[48] = IN1[48]&IN2[7];
  assign P56[48] = IN1[48]&IN2[8];
  assign P57[48] = IN1[48]&IN2[9];
  assign P58[48] = IN1[48]&IN2[10];
  assign P59[48] = IN1[48]&IN2[11];
  assign P60[48] = IN1[48]&IN2[12];
  assign P61[48] = IN1[48]&IN2[13];
  assign P62[48] = IN1[48]&IN2[14];
  assign P63[47] = IN1[48]&IN2[15];
  assign P64[46] = IN1[48]&IN2[16];
  assign P65[45] = IN1[48]&IN2[17];
  assign P66[44] = IN1[48]&IN2[18];
  assign P67[43] = IN1[48]&IN2[19];
  assign P68[42] = IN1[48]&IN2[20];
  assign P69[41] = IN1[48]&IN2[21];
  assign P70[40] = IN1[48]&IN2[22];
  assign P71[39] = IN1[48]&IN2[23];
  assign P72[38] = IN1[48]&IN2[24];
  assign P73[37] = IN1[48]&IN2[25];
  assign P74[36] = IN1[48]&IN2[26];
  assign P75[35] = IN1[48]&IN2[27];
  assign P76[34] = IN1[48]&IN2[28];
  assign P77[33] = IN1[48]&IN2[29];
  assign P78[32] = IN1[48]&IN2[30];
  assign P79[31] = IN1[48]&IN2[31];
  assign P80[30] = IN1[48]&IN2[32];
  assign P81[29] = IN1[48]&IN2[33];
  assign P82[28] = IN1[48]&IN2[34];
  assign P83[27] = IN1[48]&IN2[35];
  assign P84[26] = IN1[48]&IN2[36];
  assign P85[25] = IN1[48]&IN2[37];
  assign P86[24] = IN1[48]&IN2[38];
  assign P87[23] = IN1[48]&IN2[39];
  assign P88[22] = IN1[48]&IN2[40];
  assign P89[21] = IN1[48]&IN2[41];
  assign P90[20] = IN1[48]&IN2[42];
  assign P91[19] = IN1[48]&IN2[43];
  assign P92[18] = IN1[48]&IN2[44];
  assign P93[17] = IN1[48]&IN2[45];
  assign P94[16] = IN1[48]&IN2[46];
  assign P95[15] = IN1[48]&IN2[47];
  assign P96[14] = IN1[48]&IN2[48];
  assign P97[13] = IN1[48]&IN2[49];
  assign P98[12] = IN1[48]&IN2[50];
  assign P99[11] = IN1[48]&IN2[51];
  assign P100[10] = IN1[48]&IN2[52];
  assign P101[9] = IN1[48]&IN2[53];
  assign P102[8] = IN1[48]&IN2[54];
  assign P103[7] = IN1[48]&IN2[55];
  assign P104[6] = IN1[48]&IN2[56];
  assign P105[5] = IN1[48]&IN2[57];
  assign P106[4] = IN1[48]&IN2[58];
  assign P107[3] = IN1[48]&IN2[59];
  assign P108[2] = IN1[48]&IN2[60];
  assign P109[1] = IN1[48]&IN2[61];
  assign P110[0] = IN1[48]&IN2[62];
  assign P49[49] = IN1[49]&IN2[0];
  assign P50[49] = IN1[49]&IN2[1];
  assign P51[49] = IN1[49]&IN2[2];
  assign P52[49] = IN1[49]&IN2[3];
  assign P53[49] = IN1[49]&IN2[4];
  assign P54[49] = IN1[49]&IN2[5];
  assign P55[49] = IN1[49]&IN2[6];
  assign P56[49] = IN1[49]&IN2[7];
  assign P57[49] = IN1[49]&IN2[8];
  assign P58[49] = IN1[49]&IN2[9];
  assign P59[49] = IN1[49]&IN2[10];
  assign P60[49] = IN1[49]&IN2[11];
  assign P61[49] = IN1[49]&IN2[12];
  assign P62[49] = IN1[49]&IN2[13];
  assign P63[48] = IN1[49]&IN2[14];
  assign P64[47] = IN1[49]&IN2[15];
  assign P65[46] = IN1[49]&IN2[16];
  assign P66[45] = IN1[49]&IN2[17];
  assign P67[44] = IN1[49]&IN2[18];
  assign P68[43] = IN1[49]&IN2[19];
  assign P69[42] = IN1[49]&IN2[20];
  assign P70[41] = IN1[49]&IN2[21];
  assign P71[40] = IN1[49]&IN2[22];
  assign P72[39] = IN1[49]&IN2[23];
  assign P73[38] = IN1[49]&IN2[24];
  assign P74[37] = IN1[49]&IN2[25];
  assign P75[36] = IN1[49]&IN2[26];
  assign P76[35] = IN1[49]&IN2[27];
  assign P77[34] = IN1[49]&IN2[28];
  assign P78[33] = IN1[49]&IN2[29];
  assign P79[32] = IN1[49]&IN2[30];
  assign P80[31] = IN1[49]&IN2[31];
  assign P81[30] = IN1[49]&IN2[32];
  assign P82[29] = IN1[49]&IN2[33];
  assign P83[28] = IN1[49]&IN2[34];
  assign P84[27] = IN1[49]&IN2[35];
  assign P85[26] = IN1[49]&IN2[36];
  assign P86[25] = IN1[49]&IN2[37];
  assign P87[24] = IN1[49]&IN2[38];
  assign P88[23] = IN1[49]&IN2[39];
  assign P89[22] = IN1[49]&IN2[40];
  assign P90[21] = IN1[49]&IN2[41];
  assign P91[20] = IN1[49]&IN2[42];
  assign P92[19] = IN1[49]&IN2[43];
  assign P93[18] = IN1[49]&IN2[44];
  assign P94[17] = IN1[49]&IN2[45];
  assign P95[16] = IN1[49]&IN2[46];
  assign P96[15] = IN1[49]&IN2[47];
  assign P97[14] = IN1[49]&IN2[48];
  assign P98[13] = IN1[49]&IN2[49];
  assign P99[12] = IN1[49]&IN2[50];
  assign P100[11] = IN1[49]&IN2[51];
  assign P101[10] = IN1[49]&IN2[52];
  assign P102[9] = IN1[49]&IN2[53];
  assign P103[8] = IN1[49]&IN2[54];
  assign P104[7] = IN1[49]&IN2[55];
  assign P105[6] = IN1[49]&IN2[56];
  assign P106[5] = IN1[49]&IN2[57];
  assign P107[4] = IN1[49]&IN2[58];
  assign P108[3] = IN1[49]&IN2[59];
  assign P109[2] = IN1[49]&IN2[60];
  assign P110[1] = IN1[49]&IN2[61];
  assign P111[0] = IN1[49]&IN2[62];
  assign P50[50] = IN1[50]&IN2[0];
  assign P51[50] = IN1[50]&IN2[1];
  assign P52[50] = IN1[50]&IN2[2];
  assign P53[50] = IN1[50]&IN2[3];
  assign P54[50] = IN1[50]&IN2[4];
  assign P55[50] = IN1[50]&IN2[5];
  assign P56[50] = IN1[50]&IN2[6];
  assign P57[50] = IN1[50]&IN2[7];
  assign P58[50] = IN1[50]&IN2[8];
  assign P59[50] = IN1[50]&IN2[9];
  assign P60[50] = IN1[50]&IN2[10];
  assign P61[50] = IN1[50]&IN2[11];
  assign P62[50] = IN1[50]&IN2[12];
  assign P63[49] = IN1[50]&IN2[13];
  assign P64[48] = IN1[50]&IN2[14];
  assign P65[47] = IN1[50]&IN2[15];
  assign P66[46] = IN1[50]&IN2[16];
  assign P67[45] = IN1[50]&IN2[17];
  assign P68[44] = IN1[50]&IN2[18];
  assign P69[43] = IN1[50]&IN2[19];
  assign P70[42] = IN1[50]&IN2[20];
  assign P71[41] = IN1[50]&IN2[21];
  assign P72[40] = IN1[50]&IN2[22];
  assign P73[39] = IN1[50]&IN2[23];
  assign P74[38] = IN1[50]&IN2[24];
  assign P75[37] = IN1[50]&IN2[25];
  assign P76[36] = IN1[50]&IN2[26];
  assign P77[35] = IN1[50]&IN2[27];
  assign P78[34] = IN1[50]&IN2[28];
  assign P79[33] = IN1[50]&IN2[29];
  assign P80[32] = IN1[50]&IN2[30];
  assign P81[31] = IN1[50]&IN2[31];
  assign P82[30] = IN1[50]&IN2[32];
  assign P83[29] = IN1[50]&IN2[33];
  assign P84[28] = IN1[50]&IN2[34];
  assign P85[27] = IN1[50]&IN2[35];
  assign P86[26] = IN1[50]&IN2[36];
  assign P87[25] = IN1[50]&IN2[37];
  assign P88[24] = IN1[50]&IN2[38];
  assign P89[23] = IN1[50]&IN2[39];
  assign P90[22] = IN1[50]&IN2[40];
  assign P91[21] = IN1[50]&IN2[41];
  assign P92[20] = IN1[50]&IN2[42];
  assign P93[19] = IN1[50]&IN2[43];
  assign P94[18] = IN1[50]&IN2[44];
  assign P95[17] = IN1[50]&IN2[45];
  assign P96[16] = IN1[50]&IN2[46];
  assign P97[15] = IN1[50]&IN2[47];
  assign P98[14] = IN1[50]&IN2[48];
  assign P99[13] = IN1[50]&IN2[49];
  assign P100[12] = IN1[50]&IN2[50];
  assign P101[11] = IN1[50]&IN2[51];
  assign P102[10] = IN1[50]&IN2[52];
  assign P103[9] = IN1[50]&IN2[53];
  assign P104[8] = IN1[50]&IN2[54];
  assign P105[7] = IN1[50]&IN2[55];
  assign P106[6] = IN1[50]&IN2[56];
  assign P107[5] = IN1[50]&IN2[57];
  assign P108[4] = IN1[50]&IN2[58];
  assign P109[3] = IN1[50]&IN2[59];
  assign P110[2] = IN1[50]&IN2[60];
  assign P111[1] = IN1[50]&IN2[61];
  assign P112[0] = IN1[50]&IN2[62];
  assign P51[51] = IN1[51]&IN2[0];
  assign P52[51] = IN1[51]&IN2[1];
  assign P53[51] = IN1[51]&IN2[2];
  assign P54[51] = IN1[51]&IN2[3];
  assign P55[51] = IN1[51]&IN2[4];
  assign P56[51] = IN1[51]&IN2[5];
  assign P57[51] = IN1[51]&IN2[6];
  assign P58[51] = IN1[51]&IN2[7];
  assign P59[51] = IN1[51]&IN2[8];
  assign P60[51] = IN1[51]&IN2[9];
  assign P61[51] = IN1[51]&IN2[10];
  assign P62[51] = IN1[51]&IN2[11];
  assign P63[50] = IN1[51]&IN2[12];
  assign P64[49] = IN1[51]&IN2[13];
  assign P65[48] = IN1[51]&IN2[14];
  assign P66[47] = IN1[51]&IN2[15];
  assign P67[46] = IN1[51]&IN2[16];
  assign P68[45] = IN1[51]&IN2[17];
  assign P69[44] = IN1[51]&IN2[18];
  assign P70[43] = IN1[51]&IN2[19];
  assign P71[42] = IN1[51]&IN2[20];
  assign P72[41] = IN1[51]&IN2[21];
  assign P73[40] = IN1[51]&IN2[22];
  assign P74[39] = IN1[51]&IN2[23];
  assign P75[38] = IN1[51]&IN2[24];
  assign P76[37] = IN1[51]&IN2[25];
  assign P77[36] = IN1[51]&IN2[26];
  assign P78[35] = IN1[51]&IN2[27];
  assign P79[34] = IN1[51]&IN2[28];
  assign P80[33] = IN1[51]&IN2[29];
  assign P81[32] = IN1[51]&IN2[30];
  assign P82[31] = IN1[51]&IN2[31];
  assign P83[30] = IN1[51]&IN2[32];
  assign P84[29] = IN1[51]&IN2[33];
  assign P85[28] = IN1[51]&IN2[34];
  assign P86[27] = IN1[51]&IN2[35];
  assign P87[26] = IN1[51]&IN2[36];
  assign P88[25] = IN1[51]&IN2[37];
  assign P89[24] = IN1[51]&IN2[38];
  assign P90[23] = IN1[51]&IN2[39];
  assign P91[22] = IN1[51]&IN2[40];
  assign P92[21] = IN1[51]&IN2[41];
  assign P93[20] = IN1[51]&IN2[42];
  assign P94[19] = IN1[51]&IN2[43];
  assign P95[18] = IN1[51]&IN2[44];
  assign P96[17] = IN1[51]&IN2[45];
  assign P97[16] = IN1[51]&IN2[46];
  assign P98[15] = IN1[51]&IN2[47];
  assign P99[14] = IN1[51]&IN2[48];
  assign P100[13] = IN1[51]&IN2[49];
  assign P101[12] = IN1[51]&IN2[50];
  assign P102[11] = IN1[51]&IN2[51];
  assign P103[10] = IN1[51]&IN2[52];
  assign P104[9] = IN1[51]&IN2[53];
  assign P105[8] = IN1[51]&IN2[54];
  assign P106[7] = IN1[51]&IN2[55];
  assign P107[6] = IN1[51]&IN2[56];
  assign P108[5] = IN1[51]&IN2[57];
  assign P109[4] = IN1[51]&IN2[58];
  assign P110[3] = IN1[51]&IN2[59];
  assign P111[2] = IN1[51]&IN2[60];
  assign P112[1] = IN1[51]&IN2[61];
  assign P113[0] = IN1[51]&IN2[62];
  assign P52[52] = IN1[52]&IN2[0];
  assign P53[52] = IN1[52]&IN2[1];
  assign P54[52] = IN1[52]&IN2[2];
  assign P55[52] = IN1[52]&IN2[3];
  assign P56[52] = IN1[52]&IN2[4];
  assign P57[52] = IN1[52]&IN2[5];
  assign P58[52] = IN1[52]&IN2[6];
  assign P59[52] = IN1[52]&IN2[7];
  assign P60[52] = IN1[52]&IN2[8];
  assign P61[52] = IN1[52]&IN2[9];
  assign P62[52] = IN1[52]&IN2[10];
  assign P63[51] = IN1[52]&IN2[11];
  assign P64[50] = IN1[52]&IN2[12];
  assign P65[49] = IN1[52]&IN2[13];
  assign P66[48] = IN1[52]&IN2[14];
  assign P67[47] = IN1[52]&IN2[15];
  assign P68[46] = IN1[52]&IN2[16];
  assign P69[45] = IN1[52]&IN2[17];
  assign P70[44] = IN1[52]&IN2[18];
  assign P71[43] = IN1[52]&IN2[19];
  assign P72[42] = IN1[52]&IN2[20];
  assign P73[41] = IN1[52]&IN2[21];
  assign P74[40] = IN1[52]&IN2[22];
  assign P75[39] = IN1[52]&IN2[23];
  assign P76[38] = IN1[52]&IN2[24];
  assign P77[37] = IN1[52]&IN2[25];
  assign P78[36] = IN1[52]&IN2[26];
  assign P79[35] = IN1[52]&IN2[27];
  assign P80[34] = IN1[52]&IN2[28];
  assign P81[33] = IN1[52]&IN2[29];
  assign P82[32] = IN1[52]&IN2[30];
  assign P83[31] = IN1[52]&IN2[31];
  assign P84[30] = IN1[52]&IN2[32];
  assign P85[29] = IN1[52]&IN2[33];
  assign P86[28] = IN1[52]&IN2[34];
  assign P87[27] = IN1[52]&IN2[35];
  assign P88[26] = IN1[52]&IN2[36];
  assign P89[25] = IN1[52]&IN2[37];
  assign P90[24] = IN1[52]&IN2[38];
  assign P91[23] = IN1[52]&IN2[39];
  assign P92[22] = IN1[52]&IN2[40];
  assign P93[21] = IN1[52]&IN2[41];
  assign P94[20] = IN1[52]&IN2[42];
  assign P95[19] = IN1[52]&IN2[43];
  assign P96[18] = IN1[52]&IN2[44];
  assign P97[17] = IN1[52]&IN2[45];
  assign P98[16] = IN1[52]&IN2[46];
  assign P99[15] = IN1[52]&IN2[47];
  assign P100[14] = IN1[52]&IN2[48];
  assign P101[13] = IN1[52]&IN2[49];
  assign P102[12] = IN1[52]&IN2[50];
  assign P103[11] = IN1[52]&IN2[51];
  assign P104[10] = IN1[52]&IN2[52];
  assign P105[9] = IN1[52]&IN2[53];
  assign P106[8] = IN1[52]&IN2[54];
  assign P107[7] = IN1[52]&IN2[55];
  assign P108[6] = IN1[52]&IN2[56];
  assign P109[5] = IN1[52]&IN2[57];
  assign P110[4] = IN1[52]&IN2[58];
  assign P111[3] = IN1[52]&IN2[59];
  assign P112[2] = IN1[52]&IN2[60];
  assign P113[1] = IN1[52]&IN2[61];
  assign P114[0] = IN1[52]&IN2[62];
  assign P53[53] = IN1[53]&IN2[0];
  assign P54[53] = IN1[53]&IN2[1];
  assign P55[53] = IN1[53]&IN2[2];
  assign P56[53] = IN1[53]&IN2[3];
  assign P57[53] = IN1[53]&IN2[4];
  assign P58[53] = IN1[53]&IN2[5];
  assign P59[53] = IN1[53]&IN2[6];
  assign P60[53] = IN1[53]&IN2[7];
  assign P61[53] = IN1[53]&IN2[8];
  assign P62[53] = IN1[53]&IN2[9];
  assign P63[52] = IN1[53]&IN2[10];
  assign P64[51] = IN1[53]&IN2[11];
  assign P65[50] = IN1[53]&IN2[12];
  assign P66[49] = IN1[53]&IN2[13];
  assign P67[48] = IN1[53]&IN2[14];
  assign P68[47] = IN1[53]&IN2[15];
  assign P69[46] = IN1[53]&IN2[16];
  assign P70[45] = IN1[53]&IN2[17];
  assign P71[44] = IN1[53]&IN2[18];
  assign P72[43] = IN1[53]&IN2[19];
  assign P73[42] = IN1[53]&IN2[20];
  assign P74[41] = IN1[53]&IN2[21];
  assign P75[40] = IN1[53]&IN2[22];
  assign P76[39] = IN1[53]&IN2[23];
  assign P77[38] = IN1[53]&IN2[24];
  assign P78[37] = IN1[53]&IN2[25];
  assign P79[36] = IN1[53]&IN2[26];
  assign P80[35] = IN1[53]&IN2[27];
  assign P81[34] = IN1[53]&IN2[28];
  assign P82[33] = IN1[53]&IN2[29];
  assign P83[32] = IN1[53]&IN2[30];
  assign P84[31] = IN1[53]&IN2[31];
  assign P85[30] = IN1[53]&IN2[32];
  assign P86[29] = IN1[53]&IN2[33];
  assign P87[28] = IN1[53]&IN2[34];
  assign P88[27] = IN1[53]&IN2[35];
  assign P89[26] = IN1[53]&IN2[36];
  assign P90[25] = IN1[53]&IN2[37];
  assign P91[24] = IN1[53]&IN2[38];
  assign P92[23] = IN1[53]&IN2[39];
  assign P93[22] = IN1[53]&IN2[40];
  assign P94[21] = IN1[53]&IN2[41];
  assign P95[20] = IN1[53]&IN2[42];
  assign P96[19] = IN1[53]&IN2[43];
  assign P97[18] = IN1[53]&IN2[44];
  assign P98[17] = IN1[53]&IN2[45];
  assign P99[16] = IN1[53]&IN2[46];
  assign P100[15] = IN1[53]&IN2[47];
  assign P101[14] = IN1[53]&IN2[48];
  assign P102[13] = IN1[53]&IN2[49];
  assign P103[12] = IN1[53]&IN2[50];
  assign P104[11] = IN1[53]&IN2[51];
  assign P105[10] = IN1[53]&IN2[52];
  assign P106[9] = IN1[53]&IN2[53];
  assign P107[8] = IN1[53]&IN2[54];
  assign P108[7] = IN1[53]&IN2[55];
  assign P109[6] = IN1[53]&IN2[56];
  assign P110[5] = IN1[53]&IN2[57];
  assign P111[4] = IN1[53]&IN2[58];
  assign P112[3] = IN1[53]&IN2[59];
  assign P113[2] = IN1[53]&IN2[60];
  assign P114[1] = IN1[53]&IN2[61];
  assign P115[0] = IN1[53]&IN2[62];
  assign P54[54] = IN1[54]&IN2[0];
  assign P55[54] = IN1[54]&IN2[1];
  assign P56[54] = IN1[54]&IN2[2];
  assign P57[54] = IN1[54]&IN2[3];
  assign P58[54] = IN1[54]&IN2[4];
  assign P59[54] = IN1[54]&IN2[5];
  assign P60[54] = IN1[54]&IN2[6];
  assign P61[54] = IN1[54]&IN2[7];
  assign P62[54] = IN1[54]&IN2[8];
  assign P63[53] = IN1[54]&IN2[9];
  assign P64[52] = IN1[54]&IN2[10];
  assign P65[51] = IN1[54]&IN2[11];
  assign P66[50] = IN1[54]&IN2[12];
  assign P67[49] = IN1[54]&IN2[13];
  assign P68[48] = IN1[54]&IN2[14];
  assign P69[47] = IN1[54]&IN2[15];
  assign P70[46] = IN1[54]&IN2[16];
  assign P71[45] = IN1[54]&IN2[17];
  assign P72[44] = IN1[54]&IN2[18];
  assign P73[43] = IN1[54]&IN2[19];
  assign P74[42] = IN1[54]&IN2[20];
  assign P75[41] = IN1[54]&IN2[21];
  assign P76[40] = IN1[54]&IN2[22];
  assign P77[39] = IN1[54]&IN2[23];
  assign P78[38] = IN1[54]&IN2[24];
  assign P79[37] = IN1[54]&IN2[25];
  assign P80[36] = IN1[54]&IN2[26];
  assign P81[35] = IN1[54]&IN2[27];
  assign P82[34] = IN1[54]&IN2[28];
  assign P83[33] = IN1[54]&IN2[29];
  assign P84[32] = IN1[54]&IN2[30];
  assign P85[31] = IN1[54]&IN2[31];
  assign P86[30] = IN1[54]&IN2[32];
  assign P87[29] = IN1[54]&IN2[33];
  assign P88[28] = IN1[54]&IN2[34];
  assign P89[27] = IN1[54]&IN2[35];
  assign P90[26] = IN1[54]&IN2[36];
  assign P91[25] = IN1[54]&IN2[37];
  assign P92[24] = IN1[54]&IN2[38];
  assign P93[23] = IN1[54]&IN2[39];
  assign P94[22] = IN1[54]&IN2[40];
  assign P95[21] = IN1[54]&IN2[41];
  assign P96[20] = IN1[54]&IN2[42];
  assign P97[19] = IN1[54]&IN2[43];
  assign P98[18] = IN1[54]&IN2[44];
  assign P99[17] = IN1[54]&IN2[45];
  assign P100[16] = IN1[54]&IN2[46];
  assign P101[15] = IN1[54]&IN2[47];
  assign P102[14] = IN1[54]&IN2[48];
  assign P103[13] = IN1[54]&IN2[49];
  assign P104[12] = IN1[54]&IN2[50];
  assign P105[11] = IN1[54]&IN2[51];
  assign P106[10] = IN1[54]&IN2[52];
  assign P107[9] = IN1[54]&IN2[53];
  assign P108[8] = IN1[54]&IN2[54];
  assign P109[7] = IN1[54]&IN2[55];
  assign P110[6] = IN1[54]&IN2[56];
  assign P111[5] = IN1[54]&IN2[57];
  assign P112[4] = IN1[54]&IN2[58];
  assign P113[3] = IN1[54]&IN2[59];
  assign P114[2] = IN1[54]&IN2[60];
  assign P115[1] = IN1[54]&IN2[61];
  assign P116[0] = IN1[54]&IN2[62];
  assign P55[55] = IN1[55]&IN2[0];
  assign P56[55] = IN1[55]&IN2[1];
  assign P57[55] = IN1[55]&IN2[2];
  assign P58[55] = IN1[55]&IN2[3];
  assign P59[55] = IN1[55]&IN2[4];
  assign P60[55] = IN1[55]&IN2[5];
  assign P61[55] = IN1[55]&IN2[6];
  assign P62[55] = IN1[55]&IN2[7];
  assign P63[54] = IN1[55]&IN2[8];
  assign P64[53] = IN1[55]&IN2[9];
  assign P65[52] = IN1[55]&IN2[10];
  assign P66[51] = IN1[55]&IN2[11];
  assign P67[50] = IN1[55]&IN2[12];
  assign P68[49] = IN1[55]&IN2[13];
  assign P69[48] = IN1[55]&IN2[14];
  assign P70[47] = IN1[55]&IN2[15];
  assign P71[46] = IN1[55]&IN2[16];
  assign P72[45] = IN1[55]&IN2[17];
  assign P73[44] = IN1[55]&IN2[18];
  assign P74[43] = IN1[55]&IN2[19];
  assign P75[42] = IN1[55]&IN2[20];
  assign P76[41] = IN1[55]&IN2[21];
  assign P77[40] = IN1[55]&IN2[22];
  assign P78[39] = IN1[55]&IN2[23];
  assign P79[38] = IN1[55]&IN2[24];
  assign P80[37] = IN1[55]&IN2[25];
  assign P81[36] = IN1[55]&IN2[26];
  assign P82[35] = IN1[55]&IN2[27];
  assign P83[34] = IN1[55]&IN2[28];
  assign P84[33] = IN1[55]&IN2[29];
  assign P85[32] = IN1[55]&IN2[30];
  assign P86[31] = IN1[55]&IN2[31];
  assign P87[30] = IN1[55]&IN2[32];
  assign P88[29] = IN1[55]&IN2[33];
  assign P89[28] = IN1[55]&IN2[34];
  assign P90[27] = IN1[55]&IN2[35];
  assign P91[26] = IN1[55]&IN2[36];
  assign P92[25] = IN1[55]&IN2[37];
  assign P93[24] = IN1[55]&IN2[38];
  assign P94[23] = IN1[55]&IN2[39];
  assign P95[22] = IN1[55]&IN2[40];
  assign P96[21] = IN1[55]&IN2[41];
  assign P97[20] = IN1[55]&IN2[42];
  assign P98[19] = IN1[55]&IN2[43];
  assign P99[18] = IN1[55]&IN2[44];
  assign P100[17] = IN1[55]&IN2[45];
  assign P101[16] = IN1[55]&IN2[46];
  assign P102[15] = IN1[55]&IN2[47];
  assign P103[14] = IN1[55]&IN2[48];
  assign P104[13] = IN1[55]&IN2[49];
  assign P105[12] = IN1[55]&IN2[50];
  assign P106[11] = IN1[55]&IN2[51];
  assign P107[10] = IN1[55]&IN2[52];
  assign P108[9] = IN1[55]&IN2[53];
  assign P109[8] = IN1[55]&IN2[54];
  assign P110[7] = IN1[55]&IN2[55];
  assign P111[6] = IN1[55]&IN2[56];
  assign P112[5] = IN1[55]&IN2[57];
  assign P113[4] = IN1[55]&IN2[58];
  assign P114[3] = IN1[55]&IN2[59];
  assign P115[2] = IN1[55]&IN2[60];
  assign P116[1] = IN1[55]&IN2[61];
  assign P117[0] = IN1[55]&IN2[62];
  assign P56[56] = IN1[56]&IN2[0];
  assign P57[56] = IN1[56]&IN2[1];
  assign P58[56] = IN1[56]&IN2[2];
  assign P59[56] = IN1[56]&IN2[3];
  assign P60[56] = IN1[56]&IN2[4];
  assign P61[56] = IN1[56]&IN2[5];
  assign P62[56] = IN1[56]&IN2[6];
  assign P63[55] = IN1[56]&IN2[7];
  assign P64[54] = IN1[56]&IN2[8];
  assign P65[53] = IN1[56]&IN2[9];
  assign P66[52] = IN1[56]&IN2[10];
  assign P67[51] = IN1[56]&IN2[11];
  assign P68[50] = IN1[56]&IN2[12];
  assign P69[49] = IN1[56]&IN2[13];
  assign P70[48] = IN1[56]&IN2[14];
  assign P71[47] = IN1[56]&IN2[15];
  assign P72[46] = IN1[56]&IN2[16];
  assign P73[45] = IN1[56]&IN2[17];
  assign P74[44] = IN1[56]&IN2[18];
  assign P75[43] = IN1[56]&IN2[19];
  assign P76[42] = IN1[56]&IN2[20];
  assign P77[41] = IN1[56]&IN2[21];
  assign P78[40] = IN1[56]&IN2[22];
  assign P79[39] = IN1[56]&IN2[23];
  assign P80[38] = IN1[56]&IN2[24];
  assign P81[37] = IN1[56]&IN2[25];
  assign P82[36] = IN1[56]&IN2[26];
  assign P83[35] = IN1[56]&IN2[27];
  assign P84[34] = IN1[56]&IN2[28];
  assign P85[33] = IN1[56]&IN2[29];
  assign P86[32] = IN1[56]&IN2[30];
  assign P87[31] = IN1[56]&IN2[31];
  assign P88[30] = IN1[56]&IN2[32];
  assign P89[29] = IN1[56]&IN2[33];
  assign P90[28] = IN1[56]&IN2[34];
  assign P91[27] = IN1[56]&IN2[35];
  assign P92[26] = IN1[56]&IN2[36];
  assign P93[25] = IN1[56]&IN2[37];
  assign P94[24] = IN1[56]&IN2[38];
  assign P95[23] = IN1[56]&IN2[39];
  assign P96[22] = IN1[56]&IN2[40];
  assign P97[21] = IN1[56]&IN2[41];
  assign P98[20] = IN1[56]&IN2[42];
  assign P99[19] = IN1[56]&IN2[43];
  assign P100[18] = IN1[56]&IN2[44];
  assign P101[17] = IN1[56]&IN2[45];
  assign P102[16] = IN1[56]&IN2[46];
  assign P103[15] = IN1[56]&IN2[47];
  assign P104[14] = IN1[56]&IN2[48];
  assign P105[13] = IN1[56]&IN2[49];
  assign P106[12] = IN1[56]&IN2[50];
  assign P107[11] = IN1[56]&IN2[51];
  assign P108[10] = IN1[56]&IN2[52];
  assign P109[9] = IN1[56]&IN2[53];
  assign P110[8] = IN1[56]&IN2[54];
  assign P111[7] = IN1[56]&IN2[55];
  assign P112[6] = IN1[56]&IN2[56];
  assign P113[5] = IN1[56]&IN2[57];
  assign P114[4] = IN1[56]&IN2[58];
  assign P115[3] = IN1[56]&IN2[59];
  assign P116[2] = IN1[56]&IN2[60];
  assign P117[1] = IN1[56]&IN2[61];
  assign P118[0] = IN1[56]&IN2[62];
  assign P57[57] = IN1[57]&IN2[0];
  assign P58[57] = IN1[57]&IN2[1];
  assign P59[57] = IN1[57]&IN2[2];
  assign P60[57] = IN1[57]&IN2[3];
  assign P61[57] = IN1[57]&IN2[4];
  assign P62[57] = IN1[57]&IN2[5];
  assign P63[56] = IN1[57]&IN2[6];
  assign P64[55] = IN1[57]&IN2[7];
  assign P65[54] = IN1[57]&IN2[8];
  assign P66[53] = IN1[57]&IN2[9];
  assign P67[52] = IN1[57]&IN2[10];
  assign P68[51] = IN1[57]&IN2[11];
  assign P69[50] = IN1[57]&IN2[12];
  assign P70[49] = IN1[57]&IN2[13];
  assign P71[48] = IN1[57]&IN2[14];
  assign P72[47] = IN1[57]&IN2[15];
  assign P73[46] = IN1[57]&IN2[16];
  assign P74[45] = IN1[57]&IN2[17];
  assign P75[44] = IN1[57]&IN2[18];
  assign P76[43] = IN1[57]&IN2[19];
  assign P77[42] = IN1[57]&IN2[20];
  assign P78[41] = IN1[57]&IN2[21];
  assign P79[40] = IN1[57]&IN2[22];
  assign P80[39] = IN1[57]&IN2[23];
  assign P81[38] = IN1[57]&IN2[24];
  assign P82[37] = IN1[57]&IN2[25];
  assign P83[36] = IN1[57]&IN2[26];
  assign P84[35] = IN1[57]&IN2[27];
  assign P85[34] = IN1[57]&IN2[28];
  assign P86[33] = IN1[57]&IN2[29];
  assign P87[32] = IN1[57]&IN2[30];
  assign P88[31] = IN1[57]&IN2[31];
  assign P89[30] = IN1[57]&IN2[32];
  assign P90[29] = IN1[57]&IN2[33];
  assign P91[28] = IN1[57]&IN2[34];
  assign P92[27] = IN1[57]&IN2[35];
  assign P93[26] = IN1[57]&IN2[36];
  assign P94[25] = IN1[57]&IN2[37];
  assign P95[24] = IN1[57]&IN2[38];
  assign P96[23] = IN1[57]&IN2[39];
  assign P97[22] = IN1[57]&IN2[40];
  assign P98[21] = IN1[57]&IN2[41];
  assign P99[20] = IN1[57]&IN2[42];
  assign P100[19] = IN1[57]&IN2[43];
  assign P101[18] = IN1[57]&IN2[44];
  assign P102[17] = IN1[57]&IN2[45];
  assign P103[16] = IN1[57]&IN2[46];
  assign P104[15] = IN1[57]&IN2[47];
  assign P105[14] = IN1[57]&IN2[48];
  assign P106[13] = IN1[57]&IN2[49];
  assign P107[12] = IN1[57]&IN2[50];
  assign P108[11] = IN1[57]&IN2[51];
  assign P109[10] = IN1[57]&IN2[52];
  assign P110[9] = IN1[57]&IN2[53];
  assign P111[8] = IN1[57]&IN2[54];
  assign P112[7] = IN1[57]&IN2[55];
  assign P113[6] = IN1[57]&IN2[56];
  assign P114[5] = IN1[57]&IN2[57];
  assign P115[4] = IN1[57]&IN2[58];
  assign P116[3] = IN1[57]&IN2[59];
  assign P117[2] = IN1[57]&IN2[60];
  assign P118[1] = IN1[57]&IN2[61];
  assign P119[0] = IN1[57]&IN2[62];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, IN79, IN80, IN81, IN82, IN83, IN84, IN85, IN86, IN87, IN88, IN89, IN90, IN91, IN92, IN93, IN94, IN95, IN96, IN97, IN98, IN99, IN100, IN101, IN102, IN103, IN104, IN105, IN106, IN107, IN108, IN109, IN110, IN111, IN112, IN113, IN114, IN115, IN116, IN117, IN118, IN119, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [29:0] IN29;
  input [30:0] IN30;
  input [31:0] IN31;
  input [32:0] IN32;
  input [33:0] IN33;
  input [34:0] IN34;
  input [35:0] IN35;
  input [36:0] IN36;
  input [37:0] IN37;
  input [38:0] IN38;
  input [39:0] IN39;
  input [40:0] IN40;
  input [41:0] IN41;
  input [42:0] IN42;
  input [43:0] IN43;
  input [44:0] IN44;
  input [45:0] IN45;
  input [46:0] IN46;
  input [47:0] IN47;
  input [48:0] IN48;
  input [49:0] IN49;
  input [50:0] IN50;
  input [51:0] IN51;
  input [52:0] IN52;
  input [53:0] IN53;
  input [54:0] IN54;
  input [55:0] IN55;
  input [56:0] IN56;
  input [57:0] IN57;
  input [57:0] IN58;
  input [57:0] IN59;
  input [57:0] IN60;
  input [57:0] IN61;
  input [57:0] IN62;
  input [56:0] IN63;
  input [55:0] IN64;
  input [54:0] IN65;
  input [53:0] IN66;
  input [52:0] IN67;
  input [51:0] IN68;
  input [50:0] IN69;
  input [49:0] IN70;
  input [48:0] IN71;
  input [47:0] IN72;
  input [46:0] IN73;
  input [45:0] IN74;
  input [44:0] IN75;
  input [43:0] IN76;
  input [42:0] IN77;
  input [41:0] IN78;
  input [40:0] IN79;
  input [39:0] IN80;
  input [38:0] IN81;
  input [37:0] IN82;
  input [36:0] IN83;
  input [35:0] IN84;
  input [34:0] IN85;
  input [33:0] IN86;
  input [32:0] IN87;
  input [31:0] IN88;
  input [30:0] IN89;
  input [29:0] IN90;
  input [28:0] IN91;
  input [27:0] IN92;
  input [26:0] IN93;
  input [25:0] IN94;
  input [24:0] IN95;
  input [23:0] IN96;
  input [22:0] IN97;
  input [21:0] IN98;
  input [20:0] IN99;
  input [19:0] IN100;
  input [18:0] IN101;
  input [17:0] IN102;
  input [16:0] IN103;
  input [15:0] IN104;
  input [14:0] IN105;
  input [13:0] IN106;
  input [12:0] IN107;
  input [11:0] IN108;
  input [10:0] IN109;
  input [9:0] IN110;
  input [8:0] IN111;
  input [7:0] IN112;
  input [6:0] IN113;
  input [5:0] IN114;
  input [4:0] IN115;
  input [3:0] IN116;
  input [2:0] IN117;
  input [1:0] IN118;
  input [0:0] IN119;
  output [119:0] Out1;
  output [61:0] Out2;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3662;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3685;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3734;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3742;
  wire w3743;
  wire w3744;
  wire w3745;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3762;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3785;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3814;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3836;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3849;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3862;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3883;
  wire w3884;
  wire w3885;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3894;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3930;
  wire w3931;
  wire w3932;
  wire w3933;
  wire w3934;
  wire w3935;
  wire w3936;
  wire w3937;
  wire w3938;
  wire w3939;
  wire w3940;
  wire w3941;
  wire w3942;
  wire w3943;
  wire w3944;
  wire w3945;
  wire w3946;
  wire w3947;
  wire w3948;
  wire w3949;
  wire w3950;
  wire w3951;
  wire w3952;
  wire w3953;
  wire w3954;
  wire w3955;
  wire w3956;
  wire w3957;
  wire w3958;
  wire w3959;
  wire w3960;
  wire w3961;
  wire w3962;
  wire w3963;
  wire w3964;
  wire w3965;
  wire w3966;
  wire w3967;
  wire w3968;
  wire w3969;
  wire w3970;
  wire w3971;
  wire w3972;
  wire w3973;
  wire w3974;
  wire w3975;
  wire w3976;
  wire w3977;
  wire w3978;
  wire w3979;
  wire w3980;
  wire w3981;
  wire w3982;
  wire w3983;
  wire w3984;
  wire w3985;
  wire w3986;
  wire w3987;
  wire w3988;
  wire w3989;
  wire w3990;
  wire w3991;
  wire w3992;
  wire w3993;
  wire w3994;
  wire w3995;
  wire w3997;
  wire w3998;
  wire w3999;
  wire w4000;
  wire w4001;
  wire w4002;
  wire w4003;
  wire w4004;
  wire w4005;
  wire w4006;
  wire w4007;
  wire w4008;
  wire w4009;
  wire w4010;
  wire w4011;
  wire w4012;
  wire w4013;
  wire w4014;
  wire w4015;
  wire w4016;
  wire w4017;
  wire w4018;
  wire w4019;
  wire w4020;
  wire w4021;
  wire w4022;
  wire w4023;
  wire w4024;
  wire w4025;
  wire w4026;
  wire w4027;
  wire w4028;
  wire w4029;
  wire w4030;
  wire w4031;
  wire w4032;
  wire w4033;
  wire w4034;
  wire w4035;
  wire w4036;
  wire w4037;
  wire w4038;
  wire w4039;
  wire w4040;
  wire w4041;
  wire w4042;
  wire w4043;
  wire w4044;
  wire w4045;
  wire w4046;
  wire w4047;
  wire w4048;
  wire w4049;
  wire w4050;
  wire w4051;
  wire w4052;
  wire w4053;
  wire w4054;
  wire w4055;
  wire w4056;
  wire w4057;
  wire w4058;
  wire w4059;
  wire w4060;
  wire w4061;
  wire w4062;
  wire w4063;
  wire w4064;
  wire w4065;
  wire w4066;
  wire w4067;
  wire w4068;
  wire w4069;
  wire w4070;
  wire w4071;
  wire w4072;
  wire w4073;
  wire w4074;
  wire w4075;
  wire w4076;
  wire w4077;
  wire w4078;
  wire w4079;
  wire w4080;
  wire w4081;
  wire w4082;
  wire w4083;
  wire w4084;
  wire w4085;
  wire w4086;
  wire w4087;
  wire w4088;
  wire w4089;
  wire w4090;
  wire w4091;
  wire w4092;
  wire w4093;
  wire w4094;
  wire w4095;
  wire w4096;
  wire w4097;
  wire w4098;
  wire w4099;
  wire w4100;
  wire w4101;
  wire w4102;
  wire w4103;
  wire w4104;
  wire w4105;
  wire w4106;
  wire w4107;
  wire w4108;
  wire w4109;
  wire w4111;
  wire w4112;
  wire w4113;
  wire w4114;
  wire w4115;
  wire w4116;
  wire w4117;
  wire w4118;
  wire w4119;
  wire w4120;
  wire w4121;
  wire w4122;
  wire w4123;
  wire w4124;
  wire w4125;
  wire w4126;
  wire w4127;
  wire w4128;
  wire w4129;
  wire w4130;
  wire w4131;
  wire w4132;
  wire w4133;
  wire w4134;
  wire w4135;
  wire w4136;
  wire w4137;
  wire w4138;
  wire w4139;
  wire w4140;
  wire w4141;
  wire w4142;
  wire w4143;
  wire w4144;
  wire w4145;
  wire w4146;
  wire w4147;
  wire w4148;
  wire w4149;
  wire w4150;
  wire w4151;
  wire w4152;
  wire w4153;
  wire w4154;
  wire w4155;
  wire w4156;
  wire w4157;
  wire w4158;
  wire w4159;
  wire w4160;
  wire w4161;
  wire w4162;
  wire w4163;
  wire w4164;
  wire w4165;
  wire w4166;
  wire w4167;
  wire w4168;
  wire w4169;
  wire w4170;
  wire w4171;
  wire w4172;
  wire w4173;
  wire w4174;
  wire w4175;
  wire w4176;
  wire w4177;
  wire w4178;
  wire w4179;
  wire w4180;
  wire w4181;
  wire w4182;
  wire w4183;
  wire w4184;
  wire w4185;
  wire w4186;
  wire w4187;
  wire w4188;
  wire w4189;
  wire w4190;
  wire w4191;
  wire w4192;
  wire w4193;
  wire w4194;
  wire w4195;
  wire w4196;
  wire w4197;
  wire w4198;
  wire w4199;
  wire w4200;
  wire w4201;
  wire w4202;
  wire w4203;
  wire w4204;
  wire w4205;
  wire w4206;
  wire w4207;
  wire w4208;
  wire w4209;
  wire w4210;
  wire w4211;
  wire w4212;
  wire w4213;
  wire w4214;
  wire w4215;
  wire w4216;
  wire w4217;
  wire w4218;
  wire w4219;
  wire w4220;
  wire w4221;
  wire w4222;
  wire w4223;
  wire w4225;
  wire w4226;
  wire w4227;
  wire w4228;
  wire w4229;
  wire w4230;
  wire w4231;
  wire w4232;
  wire w4233;
  wire w4234;
  wire w4235;
  wire w4236;
  wire w4237;
  wire w4238;
  wire w4239;
  wire w4240;
  wire w4241;
  wire w4242;
  wire w4243;
  wire w4244;
  wire w4245;
  wire w4246;
  wire w4247;
  wire w4248;
  wire w4249;
  wire w4250;
  wire w4251;
  wire w4252;
  wire w4253;
  wire w4254;
  wire w4255;
  wire w4256;
  wire w4257;
  wire w4258;
  wire w4259;
  wire w4260;
  wire w4261;
  wire w4262;
  wire w4263;
  wire w4264;
  wire w4265;
  wire w4266;
  wire w4267;
  wire w4268;
  wire w4269;
  wire w4270;
  wire w4271;
  wire w4272;
  wire w4273;
  wire w4274;
  wire w4275;
  wire w4276;
  wire w4277;
  wire w4278;
  wire w4279;
  wire w4280;
  wire w4281;
  wire w4282;
  wire w4283;
  wire w4284;
  wire w4285;
  wire w4286;
  wire w4287;
  wire w4288;
  wire w4289;
  wire w4290;
  wire w4291;
  wire w4292;
  wire w4293;
  wire w4294;
  wire w4295;
  wire w4296;
  wire w4297;
  wire w4298;
  wire w4299;
  wire w4300;
  wire w4301;
  wire w4302;
  wire w4303;
  wire w4304;
  wire w4305;
  wire w4306;
  wire w4307;
  wire w4308;
  wire w4309;
  wire w4310;
  wire w4311;
  wire w4312;
  wire w4313;
  wire w4314;
  wire w4315;
  wire w4316;
  wire w4317;
  wire w4318;
  wire w4319;
  wire w4320;
  wire w4321;
  wire w4322;
  wire w4323;
  wire w4324;
  wire w4325;
  wire w4326;
  wire w4327;
  wire w4328;
  wire w4329;
  wire w4330;
  wire w4331;
  wire w4332;
  wire w4333;
  wire w4334;
  wire w4335;
  wire w4336;
  wire w4337;
  wire w4339;
  wire w4340;
  wire w4341;
  wire w4342;
  wire w4343;
  wire w4344;
  wire w4345;
  wire w4346;
  wire w4347;
  wire w4348;
  wire w4349;
  wire w4350;
  wire w4351;
  wire w4352;
  wire w4353;
  wire w4354;
  wire w4355;
  wire w4356;
  wire w4357;
  wire w4358;
  wire w4359;
  wire w4360;
  wire w4361;
  wire w4362;
  wire w4363;
  wire w4364;
  wire w4365;
  wire w4366;
  wire w4367;
  wire w4368;
  wire w4369;
  wire w4370;
  wire w4371;
  wire w4372;
  wire w4373;
  wire w4374;
  wire w4375;
  wire w4376;
  wire w4377;
  wire w4378;
  wire w4379;
  wire w4380;
  wire w4381;
  wire w4382;
  wire w4383;
  wire w4384;
  wire w4385;
  wire w4386;
  wire w4387;
  wire w4388;
  wire w4389;
  wire w4390;
  wire w4391;
  wire w4392;
  wire w4393;
  wire w4394;
  wire w4395;
  wire w4396;
  wire w4397;
  wire w4398;
  wire w4399;
  wire w4400;
  wire w4401;
  wire w4402;
  wire w4403;
  wire w4404;
  wire w4405;
  wire w4406;
  wire w4407;
  wire w4408;
  wire w4409;
  wire w4410;
  wire w4411;
  wire w4412;
  wire w4413;
  wire w4414;
  wire w4415;
  wire w4416;
  wire w4417;
  wire w4418;
  wire w4419;
  wire w4420;
  wire w4421;
  wire w4422;
  wire w4423;
  wire w4424;
  wire w4425;
  wire w4426;
  wire w4427;
  wire w4428;
  wire w4429;
  wire w4430;
  wire w4431;
  wire w4432;
  wire w4433;
  wire w4434;
  wire w4435;
  wire w4436;
  wire w4437;
  wire w4438;
  wire w4439;
  wire w4440;
  wire w4441;
  wire w4442;
  wire w4443;
  wire w4444;
  wire w4445;
  wire w4446;
  wire w4447;
  wire w4448;
  wire w4449;
  wire w4450;
  wire w4451;
  wire w4453;
  wire w4454;
  wire w4455;
  wire w4456;
  wire w4457;
  wire w4458;
  wire w4459;
  wire w4460;
  wire w4461;
  wire w4462;
  wire w4463;
  wire w4464;
  wire w4465;
  wire w4466;
  wire w4467;
  wire w4468;
  wire w4469;
  wire w4470;
  wire w4471;
  wire w4472;
  wire w4473;
  wire w4474;
  wire w4475;
  wire w4476;
  wire w4477;
  wire w4478;
  wire w4479;
  wire w4480;
  wire w4481;
  wire w4482;
  wire w4483;
  wire w4484;
  wire w4485;
  wire w4486;
  wire w4487;
  wire w4488;
  wire w4489;
  wire w4490;
  wire w4491;
  wire w4492;
  wire w4493;
  wire w4494;
  wire w4495;
  wire w4496;
  wire w4497;
  wire w4498;
  wire w4499;
  wire w4500;
  wire w4501;
  wire w4502;
  wire w4503;
  wire w4504;
  wire w4505;
  wire w4506;
  wire w4507;
  wire w4508;
  wire w4509;
  wire w4510;
  wire w4511;
  wire w4512;
  wire w4513;
  wire w4514;
  wire w4515;
  wire w4516;
  wire w4517;
  wire w4518;
  wire w4519;
  wire w4520;
  wire w4521;
  wire w4522;
  wire w4523;
  wire w4524;
  wire w4525;
  wire w4526;
  wire w4527;
  wire w4528;
  wire w4529;
  wire w4530;
  wire w4531;
  wire w4532;
  wire w4533;
  wire w4534;
  wire w4535;
  wire w4536;
  wire w4537;
  wire w4538;
  wire w4539;
  wire w4540;
  wire w4541;
  wire w4542;
  wire w4543;
  wire w4544;
  wire w4545;
  wire w4546;
  wire w4547;
  wire w4548;
  wire w4549;
  wire w4550;
  wire w4551;
  wire w4552;
  wire w4553;
  wire w4554;
  wire w4555;
  wire w4556;
  wire w4557;
  wire w4558;
  wire w4559;
  wire w4560;
  wire w4561;
  wire w4562;
  wire w4563;
  wire w4564;
  wire w4565;
  wire w4567;
  wire w4568;
  wire w4569;
  wire w4570;
  wire w4571;
  wire w4572;
  wire w4573;
  wire w4574;
  wire w4575;
  wire w4576;
  wire w4577;
  wire w4578;
  wire w4579;
  wire w4580;
  wire w4581;
  wire w4582;
  wire w4583;
  wire w4584;
  wire w4585;
  wire w4586;
  wire w4587;
  wire w4588;
  wire w4589;
  wire w4590;
  wire w4591;
  wire w4592;
  wire w4593;
  wire w4594;
  wire w4595;
  wire w4596;
  wire w4597;
  wire w4598;
  wire w4599;
  wire w4600;
  wire w4601;
  wire w4602;
  wire w4603;
  wire w4604;
  wire w4605;
  wire w4606;
  wire w4607;
  wire w4608;
  wire w4609;
  wire w4610;
  wire w4611;
  wire w4612;
  wire w4613;
  wire w4614;
  wire w4615;
  wire w4616;
  wire w4617;
  wire w4618;
  wire w4619;
  wire w4620;
  wire w4621;
  wire w4622;
  wire w4623;
  wire w4624;
  wire w4625;
  wire w4626;
  wire w4627;
  wire w4628;
  wire w4629;
  wire w4630;
  wire w4631;
  wire w4632;
  wire w4633;
  wire w4634;
  wire w4635;
  wire w4636;
  wire w4637;
  wire w4638;
  wire w4639;
  wire w4640;
  wire w4641;
  wire w4642;
  wire w4643;
  wire w4644;
  wire w4645;
  wire w4646;
  wire w4647;
  wire w4648;
  wire w4649;
  wire w4650;
  wire w4651;
  wire w4652;
  wire w4653;
  wire w4654;
  wire w4655;
  wire w4656;
  wire w4657;
  wire w4658;
  wire w4659;
  wire w4660;
  wire w4661;
  wire w4662;
  wire w4663;
  wire w4664;
  wire w4665;
  wire w4666;
  wire w4667;
  wire w4668;
  wire w4669;
  wire w4670;
  wire w4671;
  wire w4672;
  wire w4673;
  wire w4674;
  wire w4675;
  wire w4676;
  wire w4677;
  wire w4678;
  wire w4679;
  wire w4681;
  wire w4682;
  wire w4683;
  wire w4684;
  wire w4685;
  wire w4686;
  wire w4687;
  wire w4688;
  wire w4689;
  wire w4690;
  wire w4691;
  wire w4692;
  wire w4693;
  wire w4694;
  wire w4695;
  wire w4696;
  wire w4697;
  wire w4698;
  wire w4699;
  wire w4700;
  wire w4701;
  wire w4702;
  wire w4703;
  wire w4704;
  wire w4705;
  wire w4706;
  wire w4707;
  wire w4708;
  wire w4709;
  wire w4710;
  wire w4711;
  wire w4712;
  wire w4713;
  wire w4714;
  wire w4715;
  wire w4716;
  wire w4717;
  wire w4718;
  wire w4719;
  wire w4720;
  wire w4721;
  wire w4722;
  wire w4723;
  wire w4724;
  wire w4725;
  wire w4726;
  wire w4727;
  wire w4728;
  wire w4729;
  wire w4730;
  wire w4731;
  wire w4732;
  wire w4733;
  wire w4734;
  wire w4735;
  wire w4736;
  wire w4737;
  wire w4738;
  wire w4739;
  wire w4740;
  wire w4741;
  wire w4742;
  wire w4743;
  wire w4744;
  wire w4745;
  wire w4746;
  wire w4747;
  wire w4748;
  wire w4749;
  wire w4750;
  wire w4751;
  wire w4752;
  wire w4753;
  wire w4754;
  wire w4755;
  wire w4756;
  wire w4757;
  wire w4758;
  wire w4759;
  wire w4760;
  wire w4761;
  wire w4762;
  wire w4763;
  wire w4764;
  wire w4765;
  wire w4766;
  wire w4767;
  wire w4768;
  wire w4769;
  wire w4770;
  wire w4771;
  wire w4772;
  wire w4773;
  wire w4774;
  wire w4775;
  wire w4776;
  wire w4777;
  wire w4778;
  wire w4779;
  wire w4780;
  wire w4781;
  wire w4782;
  wire w4783;
  wire w4784;
  wire w4785;
  wire w4786;
  wire w4787;
  wire w4788;
  wire w4789;
  wire w4790;
  wire w4791;
  wire w4792;
  wire w4793;
  wire w4795;
  wire w4796;
  wire w4797;
  wire w4798;
  wire w4799;
  wire w4800;
  wire w4801;
  wire w4802;
  wire w4803;
  wire w4804;
  wire w4805;
  wire w4806;
  wire w4807;
  wire w4808;
  wire w4809;
  wire w4810;
  wire w4811;
  wire w4812;
  wire w4813;
  wire w4814;
  wire w4815;
  wire w4816;
  wire w4817;
  wire w4818;
  wire w4819;
  wire w4820;
  wire w4821;
  wire w4822;
  wire w4823;
  wire w4824;
  wire w4825;
  wire w4826;
  wire w4827;
  wire w4828;
  wire w4829;
  wire w4830;
  wire w4831;
  wire w4832;
  wire w4833;
  wire w4834;
  wire w4835;
  wire w4836;
  wire w4837;
  wire w4838;
  wire w4839;
  wire w4840;
  wire w4841;
  wire w4842;
  wire w4843;
  wire w4844;
  wire w4845;
  wire w4846;
  wire w4847;
  wire w4848;
  wire w4849;
  wire w4850;
  wire w4851;
  wire w4852;
  wire w4853;
  wire w4854;
  wire w4855;
  wire w4856;
  wire w4857;
  wire w4858;
  wire w4859;
  wire w4860;
  wire w4861;
  wire w4862;
  wire w4863;
  wire w4864;
  wire w4865;
  wire w4866;
  wire w4867;
  wire w4868;
  wire w4869;
  wire w4870;
  wire w4871;
  wire w4872;
  wire w4873;
  wire w4874;
  wire w4875;
  wire w4876;
  wire w4877;
  wire w4878;
  wire w4879;
  wire w4880;
  wire w4881;
  wire w4882;
  wire w4883;
  wire w4884;
  wire w4885;
  wire w4886;
  wire w4887;
  wire w4888;
  wire w4889;
  wire w4890;
  wire w4891;
  wire w4892;
  wire w4893;
  wire w4894;
  wire w4895;
  wire w4896;
  wire w4897;
  wire w4898;
  wire w4899;
  wire w4900;
  wire w4901;
  wire w4902;
  wire w4903;
  wire w4904;
  wire w4905;
  wire w4906;
  wire w4907;
  wire w4909;
  wire w4910;
  wire w4911;
  wire w4912;
  wire w4913;
  wire w4914;
  wire w4915;
  wire w4916;
  wire w4917;
  wire w4918;
  wire w4919;
  wire w4920;
  wire w4921;
  wire w4922;
  wire w4923;
  wire w4924;
  wire w4925;
  wire w4926;
  wire w4927;
  wire w4928;
  wire w4929;
  wire w4930;
  wire w4931;
  wire w4932;
  wire w4933;
  wire w4934;
  wire w4935;
  wire w4936;
  wire w4937;
  wire w4938;
  wire w4939;
  wire w4940;
  wire w4941;
  wire w4942;
  wire w4943;
  wire w4944;
  wire w4945;
  wire w4946;
  wire w4947;
  wire w4948;
  wire w4949;
  wire w4950;
  wire w4951;
  wire w4952;
  wire w4953;
  wire w4954;
  wire w4955;
  wire w4956;
  wire w4957;
  wire w4958;
  wire w4959;
  wire w4960;
  wire w4961;
  wire w4962;
  wire w4963;
  wire w4964;
  wire w4965;
  wire w4966;
  wire w4967;
  wire w4968;
  wire w4969;
  wire w4970;
  wire w4971;
  wire w4972;
  wire w4973;
  wire w4974;
  wire w4975;
  wire w4976;
  wire w4977;
  wire w4978;
  wire w4979;
  wire w4980;
  wire w4981;
  wire w4982;
  wire w4983;
  wire w4984;
  wire w4985;
  wire w4986;
  wire w4987;
  wire w4988;
  wire w4989;
  wire w4990;
  wire w4991;
  wire w4992;
  wire w4993;
  wire w4994;
  wire w4995;
  wire w4996;
  wire w4997;
  wire w4998;
  wire w4999;
  wire w5000;
  wire w5001;
  wire w5002;
  wire w5003;
  wire w5004;
  wire w5005;
  wire w5006;
  wire w5007;
  wire w5008;
  wire w5009;
  wire w5010;
  wire w5011;
  wire w5012;
  wire w5013;
  wire w5014;
  wire w5015;
  wire w5016;
  wire w5017;
  wire w5018;
  wire w5019;
  wire w5020;
  wire w5021;
  wire w5023;
  wire w5024;
  wire w5025;
  wire w5026;
  wire w5027;
  wire w5028;
  wire w5029;
  wire w5030;
  wire w5031;
  wire w5032;
  wire w5033;
  wire w5034;
  wire w5035;
  wire w5036;
  wire w5037;
  wire w5038;
  wire w5039;
  wire w5040;
  wire w5041;
  wire w5042;
  wire w5043;
  wire w5044;
  wire w5045;
  wire w5046;
  wire w5047;
  wire w5048;
  wire w5049;
  wire w5050;
  wire w5051;
  wire w5052;
  wire w5053;
  wire w5054;
  wire w5055;
  wire w5056;
  wire w5057;
  wire w5058;
  wire w5059;
  wire w5060;
  wire w5061;
  wire w5062;
  wire w5063;
  wire w5064;
  wire w5065;
  wire w5066;
  wire w5067;
  wire w5068;
  wire w5069;
  wire w5070;
  wire w5071;
  wire w5072;
  wire w5073;
  wire w5074;
  wire w5075;
  wire w5076;
  wire w5077;
  wire w5078;
  wire w5079;
  wire w5080;
  wire w5081;
  wire w5082;
  wire w5083;
  wire w5084;
  wire w5085;
  wire w5086;
  wire w5087;
  wire w5088;
  wire w5089;
  wire w5090;
  wire w5091;
  wire w5092;
  wire w5093;
  wire w5094;
  wire w5095;
  wire w5096;
  wire w5097;
  wire w5098;
  wire w5099;
  wire w5100;
  wire w5101;
  wire w5102;
  wire w5103;
  wire w5104;
  wire w5105;
  wire w5106;
  wire w5107;
  wire w5108;
  wire w5109;
  wire w5110;
  wire w5111;
  wire w5112;
  wire w5113;
  wire w5114;
  wire w5115;
  wire w5116;
  wire w5117;
  wire w5118;
  wire w5119;
  wire w5120;
  wire w5121;
  wire w5122;
  wire w5123;
  wire w5124;
  wire w5125;
  wire w5126;
  wire w5127;
  wire w5128;
  wire w5129;
  wire w5130;
  wire w5131;
  wire w5132;
  wire w5133;
  wire w5134;
  wire w5135;
  wire w5137;
  wire w5138;
  wire w5139;
  wire w5140;
  wire w5141;
  wire w5142;
  wire w5143;
  wire w5144;
  wire w5145;
  wire w5146;
  wire w5147;
  wire w5148;
  wire w5149;
  wire w5150;
  wire w5151;
  wire w5152;
  wire w5153;
  wire w5154;
  wire w5155;
  wire w5156;
  wire w5157;
  wire w5158;
  wire w5159;
  wire w5160;
  wire w5161;
  wire w5162;
  wire w5163;
  wire w5164;
  wire w5165;
  wire w5166;
  wire w5167;
  wire w5168;
  wire w5169;
  wire w5170;
  wire w5171;
  wire w5172;
  wire w5173;
  wire w5174;
  wire w5175;
  wire w5176;
  wire w5177;
  wire w5178;
  wire w5179;
  wire w5180;
  wire w5181;
  wire w5182;
  wire w5183;
  wire w5184;
  wire w5185;
  wire w5186;
  wire w5187;
  wire w5188;
  wire w5189;
  wire w5190;
  wire w5191;
  wire w5192;
  wire w5193;
  wire w5194;
  wire w5195;
  wire w5196;
  wire w5197;
  wire w5198;
  wire w5199;
  wire w5200;
  wire w5201;
  wire w5202;
  wire w5203;
  wire w5204;
  wire w5205;
  wire w5206;
  wire w5207;
  wire w5208;
  wire w5209;
  wire w5210;
  wire w5211;
  wire w5212;
  wire w5213;
  wire w5214;
  wire w5215;
  wire w5216;
  wire w5217;
  wire w5218;
  wire w5219;
  wire w5220;
  wire w5221;
  wire w5222;
  wire w5223;
  wire w5224;
  wire w5225;
  wire w5226;
  wire w5227;
  wire w5228;
  wire w5229;
  wire w5230;
  wire w5231;
  wire w5232;
  wire w5233;
  wire w5234;
  wire w5235;
  wire w5236;
  wire w5237;
  wire w5238;
  wire w5239;
  wire w5240;
  wire w5241;
  wire w5242;
  wire w5243;
  wire w5244;
  wire w5245;
  wire w5246;
  wire w5247;
  wire w5248;
  wire w5249;
  wire w5251;
  wire w5252;
  wire w5253;
  wire w5254;
  wire w5255;
  wire w5256;
  wire w5257;
  wire w5258;
  wire w5259;
  wire w5260;
  wire w5261;
  wire w5262;
  wire w5263;
  wire w5264;
  wire w5265;
  wire w5266;
  wire w5267;
  wire w5268;
  wire w5269;
  wire w5270;
  wire w5271;
  wire w5272;
  wire w5273;
  wire w5274;
  wire w5275;
  wire w5276;
  wire w5277;
  wire w5278;
  wire w5279;
  wire w5280;
  wire w5281;
  wire w5282;
  wire w5283;
  wire w5284;
  wire w5285;
  wire w5286;
  wire w5287;
  wire w5288;
  wire w5289;
  wire w5290;
  wire w5291;
  wire w5292;
  wire w5293;
  wire w5294;
  wire w5295;
  wire w5296;
  wire w5297;
  wire w5298;
  wire w5299;
  wire w5300;
  wire w5301;
  wire w5302;
  wire w5303;
  wire w5304;
  wire w5305;
  wire w5306;
  wire w5307;
  wire w5308;
  wire w5309;
  wire w5310;
  wire w5311;
  wire w5312;
  wire w5313;
  wire w5314;
  wire w5315;
  wire w5316;
  wire w5317;
  wire w5318;
  wire w5319;
  wire w5320;
  wire w5321;
  wire w5322;
  wire w5323;
  wire w5324;
  wire w5325;
  wire w5326;
  wire w5327;
  wire w5328;
  wire w5329;
  wire w5330;
  wire w5331;
  wire w5332;
  wire w5333;
  wire w5334;
  wire w5335;
  wire w5336;
  wire w5337;
  wire w5338;
  wire w5339;
  wire w5340;
  wire w5341;
  wire w5342;
  wire w5343;
  wire w5344;
  wire w5345;
  wire w5346;
  wire w5347;
  wire w5348;
  wire w5349;
  wire w5350;
  wire w5351;
  wire w5352;
  wire w5353;
  wire w5354;
  wire w5355;
  wire w5356;
  wire w5357;
  wire w5358;
  wire w5359;
  wire w5360;
  wire w5361;
  wire w5362;
  wire w5363;
  wire w5365;
  wire w5366;
  wire w5367;
  wire w5368;
  wire w5369;
  wire w5370;
  wire w5371;
  wire w5372;
  wire w5373;
  wire w5374;
  wire w5375;
  wire w5376;
  wire w5377;
  wire w5378;
  wire w5379;
  wire w5380;
  wire w5381;
  wire w5382;
  wire w5383;
  wire w5384;
  wire w5385;
  wire w5386;
  wire w5387;
  wire w5388;
  wire w5389;
  wire w5390;
  wire w5391;
  wire w5392;
  wire w5393;
  wire w5394;
  wire w5395;
  wire w5396;
  wire w5397;
  wire w5398;
  wire w5399;
  wire w5400;
  wire w5401;
  wire w5402;
  wire w5403;
  wire w5404;
  wire w5405;
  wire w5406;
  wire w5407;
  wire w5408;
  wire w5409;
  wire w5410;
  wire w5411;
  wire w5412;
  wire w5413;
  wire w5414;
  wire w5415;
  wire w5416;
  wire w5417;
  wire w5418;
  wire w5419;
  wire w5420;
  wire w5421;
  wire w5422;
  wire w5423;
  wire w5424;
  wire w5425;
  wire w5426;
  wire w5427;
  wire w5428;
  wire w5429;
  wire w5430;
  wire w5431;
  wire w5432;
  wire w5433;
  wire w5434;
  wire w5435;
  wire w5436;
  wire w5437;
  wire w5438;
  wire w5439;
  wire w5440;
  wire w5441;
  wire w5442;
  wire w5443;
  wire w5444;
  wire w5445;
  wire w5446;
  wire w5447;
  wire w5448;
  wire w5449;
  wire w5450;
  wire w5451;
  wire w5452;
  wire w5453;
  wire w5454;
  wire w5455;
  wire w5456;
  wire w5457;
  wire w5458;
  wire w5459;
  wire w5460;
  wire w5461;
  wire w5462;
  wire w5463;
  wire w5464;
  wire w5465;
  wire w5466;
  wire w5467;
  wire w5468;
  wire w5469;
  wire w5470;
  wire w5471;
  wire w5472;
  wire w5473;
  wire w5474;
  wire w5475;
  wire w5476;
  wire w5477;
  wire w5479;
  wire w5480;
  wire w5481;
  wire w5482;
  wire w5483;
  wire w5484;
  wire w5485;
  wire w5486;
  wire w5487;
  wire w5488;
  wire w5489;
  wire w5490;
  wire w5491;
  wire w5492;
  wire w5493;
  wire w5494;
  wire w5495;
  wire w5496;
  wire w5497;
  wire w5498;
  wire w5499;
  wire w5500;
  wire w5501;
  wire w5502;
  wire w5503;
  wire w5504;
  wire w5505;
  wire w5506;
  wire w5507;
  wire w5508;
  wire w5509;
  wire w5510;
  wire w5511;
  wire w5512;
  wire w5513;
  wire w5514;
  wire w5515;
  wire w5516;
  wire w5517;
  wire w5518;
  wire w5519;
  wire w5520;
  wire w5521;
  wire w5522;
  wire w5523;
  wire w5524;
  wire w5525;
  wire w5526;
  wire w5527;
  wire w5528;
  wire w5529;
  wire w5530;
  wire w5531;
  wire w5532;
  wire w5533;
  wire w5534;
  wire w5535;
  wire w5536;
  wire w5537;
  wire w5538;
  wire w5539;
  wire w5540;
  wire w5541;
  wire w5542;
  wire w5543;
  wire w5544;
  wire w5545;
  wire w5546;
  wire w5547;
  wire w5548;
  wire w5549;
  wire w5550;
  wire w5551;
  wire w5552;
  wire w5553;
  wire w5554;
  wire w5555;
  wire w5556;
  wire w5557;
  wire w5558;
  wire w5559;
  wire w5560;
  wire w5561;
  wire w5562;
  wire w5563;
  wire w5564;
  wire w5565;
  wire w5566;
  wire w5567;
  wire w5568;
  wire w5569;
  wire w5570;
  wire w5571;
  wire w5572;
  wire w5573;
  wire w5574;
  wire w5575;
  wire w5576;
  wire w5577;
  wire w5578;
  wire w5579;
  wire w5580;
  wire w5581;
  wire w5582;
  wire w5583;
  wire w5584;
  wire w5585;
  wire w5586;
  wire w5587;
  wire w5588;
  wire w5589;
  wire w5590;
  wire w5591;
  wire w5593;
  wire w5594;
  wire w5595;
  wire w5596;
  wire w5597;
  wire w5598;
  wire w5599;
  wire w5600;
  wire w5601;
  wire w5602;
  wire w5603;
  wire w5604;
  wire w5605;
  wire w5606;
  wire w5607;
  wire w5608;
  wire w5609;
  wire w5610;
  wire w5611;
  wire w5612;
  wire w5613;
  wire w5614;
  wire w5615;
  wire w5616;
  wire w5617;
  wire w5618;
  wire w5619;
  wire w5620;
  wire w5621;
  wire w5622;
  wire w5623;
  wire w5624;
  wire w5625;
  wire w5626;
  wire w5627;
  wire w5628;
  wire w5629;
  wire w5630;
  wire w5631;
  wire w5632;
  wire w5633;
  wire w5634;
  wire w5635;
  wire w5636;
  wire w5637;
  wire w5638;
  wire w5639;
  wire w5640;
  wire w5641;
  wire w5642;
  wire w5643;
  wire w5644;
  wire w5645;
  wire w5646;
  wire w5647;
  wire w5648;
  wire w5649;
  wire w5650;
  wire w5651;
  wire w5652;
  wire w5653;
  wire w5654;
  wire w5655;
  wire w5656;
  wire w5657;
  wire w5658;
  wire w5659;
  wire w5660;
  wire w5661;
  wire w5662;
  wire w5663;
  wire w5664;
  wire w5665;
  wire w5666;
  wire w5667;
  wire w5668;
  wire w5669;
  wire w5670;
  wire w5671;
  wire w5672;
  wire w5673;
  wire w5674;
  wire w5675;
  wire w5676;
  wire w5677;
  wire w5678;
  wire w5679;
  wire w5680;
  wire w5681;
  wire w5682;
  wire w5683;
  wire w5684;
  wire w5685;
  wire w5686;
  wire w5687;
  wire w5688;
  wire w5689;
  wire w5690;
  wire w5691;
  wire w5692;
  wire w5693;
  wire w5694;
  wire w5695;
  wire w5696;
  wire w5697;
  wire w5698;
  wire w5699;
  wire w5700;
  wire w5701;
  wire w5702;
  wire w5703;
  wire w5704;
  wire w5705;
  wire w5707;
  wire w5708;
  wire w5709;
  wire w5710;
  wire w5711;
  wire w5712;
  wire w5713;
  wire w5714;
  wire w5715;
  wire w5716;
  wire w5717;
  wire w5718;
  wire w5719;
  wire w5720;
  wire w5721;
  wire w5722;
  wire w5723;
  wire w5724;
  wire w5725;
  wire w5726;
  wire w5727;
  wire w5728;
  wire w5729;
  wire w5730;
  wire w5731;
  wire w5732;
  wire w5733;
  wire w5734;
  wire w5735;
  wire w5736;
  wire w5737;
  wire w5738;
  wire w5739;
  wire w5740;
  wire w5741;
  wire w5742;
  wire w5743;
  wire w5744;
  wire w5745;
  wire w5746;
  wire w5747;
  wire w5748;
  wire w5749;
  wire w5750;
  wire w5751;
  wire w5752;
  wire w5753;
  wire w5754;
  wire w5755;
  wire w5756;
  wire w5757;
  wire w5758;
  wire w5759;
  wire w5760;
  wire w5761;
  wire w5762;
  wire w5763;
  wire w5764;
  wire w5765;
  wire w5766;
  wire w5767;
  wire w5768;
  wire w5769;
  wire w5770;
  wire w5771;
  wire w5772;
  wire w5773;
  wire w5774;
  wire w5775;
  wire w5776;
  wire w5777;
  wire w5778;
  wire w5779;
  wire w5780;
  wire w5781;
  wire w5782;
  wire w5783;
  wire w5784;
  wire w5785;
  wire w5786;
  wire w5787;
  wire w5788;
  wire w5789;
  wire w5790;
  wire w5791;
  wire w5792;
  wire w5793;
  wire w5794;
  wire w5795;
  wire w5796;
  wire w5797;
  wire w5798;
  wire w5799;
  wire w5800;
  wire w5801;
  wire w5802;
  wire w5803;
  wire w5804;
  wire w5805;
  wire w5806;
  wire w5807;
  wire w5808;
  wire w5809;
  wire w5810;
  wire w5811;
  wire w5812;
  wire w5813;
  wire w5814;
  wire w5815;
  wire w5816;
  wire w5817;
  wire w5818;
  wire w5819;
  wire w5821;
  wire w5822;
  wire w5823;
  wire w5824;
  wire w5825;
  wire w5826;
  wire w5827;
  wire w5828;
  wire w5829;
  wire w5830;
  wire w5831;
  wire w5832;
  wire w5833;
  wire w5834;
  wire w5835;
  wire w5836;
  wire w5837;
  wire w5838;
  wire w5839;
  wire w5840;
  wire w5841;
  wire w5842;
  wire w5843;
  wire w5844;
  wire w5845;
  wire w5846;
  wire w5847;
  wire w5848;
  wire w5849;
  wire w5850;
  wire w5851;
  wire w5852;
  wire w5853;
  wire w5854;
  wire w5855;
  wire w5856;
  wire w5857;
  wire w5858;
  wire w5859;
  wire w5860;
  wire w5861;
  wire w5862;
  wire w5863;
  wire w5864;
  wire w5865;
  wire w5866;
  wire w5867;
  wire w5868;
  wire w5869;
  wire w5870;
  wire w5871;
  wire w5872;
  wire w5873;
  wire w5874;
  wire w5875;
  wire w5876;
  wire w5877;
  wire w5878;
  wire w5879;
  wire w5880;
  wire w5881;
  wire w5882;
  wire w5883;
  wire w5884;
  wire w5885;
  wire w5886;
  wire w5887;
  wire w5888;
  wire w5889;
  wire w5890;
  wire w5891;
  wire w5892;
  wire w5893;
  wire w5894;
  wire w5895;
  wire w5896;
  wire w5897;
  wire w5898;
  wire w5899;
  wire w5900;
  wire w5901;
  wire w5902;
  wire w5903;
  wire w5904;
  wire w5905;
  wire w5906;
  wire w5907;
  wire w5908;
  wire w5909;
  wire w5910;
  wire w5911;
  wire w5912;
  wire w5913;
  wire w5914;
  wire w5915;
  wire w5916;
  wire w5917;
  wire w5918;
  wire w5919;
  wire w5920;
  wire w5921;
  wire w5922;
  wire w5923;
  wire w5924;
  wire w5925;
  wire w5926;
  wire w5927;
  wire w5928;
  wire w5929;
  wire w5930;
  wire w5931;
  wire w5932;
  wire w5933;
  wire w5935;
  wire w5936;
  wire w5937;
  wire w5938;
  wire w5939;
  wire w5940;
  wire w5941;
  wire w5942;
  wire w5943;
  wire w5944;
  wire w5945;
  wire w5946;
  wire w5947;
  wire w5948;
  wire w5949;
  wire w5950;
  wire w5951;
  wire w5952;
  wire w5953;
  wire w5954;
  wire w5955;
  wire w5956;
  wire w5957;
  wire w5958;
  wire w5959;
  wire w5960;
  wire w5961;
  wire w5962;
  wire w5963;
  wire w5964;
  wire w5965;
  wire w5966;
  wire w5967;
  wire w5968;
  wire w5969;
  wire w5970;
  wire w5971;
  wire w5972;
  wire w5973;
  wire w5974;
  wire w5975;
  wire w5976;
  wire w5977;
  wire w5978;
  wire w5979;
  wire w5980;
  wire w5981;
  wire w5982;
  wire w5983;
  wire w5984;
  wire w5985;
  wire w5986;
  wire w5987;
  wire w5988;
  wire w5989;
  wire w5990;
  wire w5991;
  wire w5992;
  wire w5993;
  wire w5994;
  wire w5995;
  wire w5996;
  wire w5997;
  wire w5998;
  wire w5999;
  wire w6000;
  wire w6001;
  wire w6002;
  wire w6003;
  wire w6004;
  wire w6005;
  wire w6006;
  wire w6007;
  wire w6008;
  wire w6009;
  wire w6010;
  wire w6011;
  wire w6012;
  wire w6013;
  wire w6014;
  wire w6015;
  wire w6016;
  wire w6017;
  wire w6018;
  wire w6019;
  wire w6020;
  wire w6021;
  wire w6022;
  wire w6023;
  wire w6024;
  wire w6025;
  wire w6026;
  wire w6027;
  wire w6028;
  wire w6029;
  wire w6030;
  wire w6031;
  wire w6032;
  wire w6033;
  wire w6034;
  wire w6035;
  wire w6036;
  wire w6037;
  wire w6038;
  wire w6039;
  wire w6040;
  wire w6041;
  wire w6042;
  wire w6043;
  wire w6044;
  wire w6045;
  wire w6046;
  wire w6047;
  wire w6049;
  wire w6050;
  wire w6051;
  wire w6052;
  wire w6053;
  wire w6054;
  wire w6055;
  wire w6056;
  wire w6057;
  wire w6058;
  wire w6059;
  wire w6060;
  wire w6061;
  wire w6062;
  wire w6063;
  wire w6064;
  wire w6065;
  wire w6066;
  wire w6067;
  wire w6068;
  wire w6069;
  wire w6070;
  wire w6071;
  wire w6072;
  wire w6073;
  wire w6074;
  wire w6075;
  wire w6076;
  wire w6077;
  wire w6078;
  wire w6079;
  wire w6080;
  wire w6081;
  wire w6082;
  wire w6083;
  wire w6084;
  wire w6085;
  wire w6086;
  wire w6087;
  wire w6088;
  wire w6089;
  wire w6090;
  wire w6091;
  wire w6092;
  wire w6093;
  wire w6094;
  wire w6095;
  wire w6096;
  wire w6097;
  wire w6098;
  wire w6099;
  wire w6100;
  wire w6101;
  wire w6102;
  wire w6103;
  wire w6104;
  wire w6105;
  wire w6106;
  wire w6107;
  wire w6108;
  wire w6109;
  wire w6110;
  wire w6111;
  wire w6112;
  wire w6113;
  wire w6114;
  wire w6115;
  wire w6116;
  wire w6117;
  wire w6118;
  wire w6119;
  wire w6120;
  wire w6121;
  wire w6122;
  wire w6123;
  wire w6124;
  wire w6125;
  wire w6126;
  wire w6127;
  wire w6128;
  wire w6129;
  wire w6130;
  wire w6131;
  wire w6132;
  wire w6133;
  wire w6134;
  wire w6135;
  wire w6136;
  wire w6137;
  wire w6138;
  wire w6139;
  wire w6140;
  wire w6141;
  wire w6142;
  wire w6143;
  wire w6144;
  wire w6145;
  wire w6146;
  wire w6147;
  wire w6148;
  wire w6149;
  wire w6150;
  wire w6151;
  wire w6152;
  wire w6153;
  wire w6154;
  wire w6155;
  wire w6156;
  wire w6157;
  wire w6158;
  wire w6159;
  wire w6160;
  wire w6161;
  wire w6163;
  wire w6164;
  wire w6165;
  wire w6166;
  wire w6167;
  wire w6168;
  wire w6169;
  wire w6170;
  wire w6171;
  wire w6172;
  wire w6173;
  wire w6174;
  wire w6175;
  wire w6176;
  wire w6177;
  wire w6178;
  wire w6179;
  wire w6180;
  wire w6181;
  wire w6182;
  wire w6183;
  wire w6184;
  wire w6185;
  wire w6186;
  wire w6187;
  wire w6188;
  wire w6189;
  wire w6190;
  wire w6191;
  wire w6192;
  wire w6193;
  wire w6194;
  wire w6195;
  wire w6196;
  wire w6197;
  wire w6198;
  wire w6199;
  wire w6200;
  wire w6201;
  wire w6202;
  wire w6203;
  wire w6204;
  wire w6205;
  wire w6206;
  wire w6207;
  wire w6208;
  wire w6209;
  wire w6210;
  wire w6211;
  wire w6212;
  wire w6213;
  wire w6214;
  wire w6215;
  wire w6216;
  wire w6217;
  wire w6218;
  wire w6219;
  wire w6220;
  wire w6221;
  wire w6222;
  wire w6223;
  wire w6224;
  wire w6225;
  wire w6226;
  wire w6227;
  wire w6228;
  wire w6229;
  wire w6230;
  wire w6231;
  wire w6232;
  wire w6233;
  wire w6234;
  wire w6235;
  wire w6236;
  wire w6237;
  wire w6238;
  wire w6239;
  wire w6240;
  wire w6241;
  wire w6242;
  wire w6243;
  wire w6244;
  wire w6245;
  wire w6246;
  wire w6247;
  wire w6248;
  wire w6249;
  wire w6250;
  wire w6251;
  wire w6252;
  wire w6253;
  wire w6254;
  wire w6255;
  wire w6256;
  wire w6257;
  wire w6258;
  wire w6259;
  wire w6260;
  wire w6261;
  wire w6262;
  wire w6263;
  wire w6264;
  wire w6265;
  wire w6266;
  wire w6267;
  wire w6268;
  wire w6269;
  wire w6270;
  wire w6271;
  wire w6272;
  wire w6273;
  wire w6274;
  wire w6275;
  wire w6277;
  wire w6278;
  wire w6279;
  wire w6280;
  wire w6281;
  wire w6282;
  wire w6283;
  wire w6284;
  wire w6285;
  wire w6286;
  wire w6287;
  wire w6288;
  wire w6289;
  wire w6290;
  wire w6291;
  wire w6292;
  wire w6293;
  wire w6294;
  wire w6295;
  wire w6296;
  wire w6297;
  wire w6298;
  wire w6299;
  wire w6300;
  wire w6301;
  wire w6302;
  wire w6303;
  wire w6304;
  wire w6305;
  wire w6306;
  wire w6307;
  wire w6308;
  wire w6309;
  wire w6310;
  wire w6311;
  wire w6312;
  wire w6313;
  wire w6314;
  wire w6315;
  wire w6316;
  wire w6317;
  wire w6318;
  wire w6319;
  wire w6320;
  wire w6321;
  wire w6322;
  wire w6323;
  wire w6324;
  wire w6325;
  wire w6326;
  wire w6327;
  wire w6328;
  wire w6329;
  wire w6330;
  wire w6331;
  wire w6332;
  wire w6333;
  wire w6334;
  wire w6335;
  wire w6336;
  wire w6337;
  wire w6338;
  wire w6339;
  wire w6340;
  wire w6341;
  wire w6342;
  wire w6343;
  wire w6344;
  wire w6345;
  wire w6346;
  wire w6347;
  wire w6348;
  wire w6349;
  wire w6350;
  wire w6351;
  wire w6352;
  wire w6353;
  wire w6354;
  wire w6355;
  wire w6356;
  wire w6357;
  wire w6358;
  wire w6359;
  wire w6360;
  wire w6361;
  wire w6362;
  wire w6363;
  wire w6364;
  wire w6365;
  wire w6366;
  wire w6367;
  wire w6368;
  wire w6369;
  wire w6370;
  wire w6371;
  wire w6372;
  wire w6373;
  wire w6374;
  wire w6375;
  wire w6376;
  wire w6377;
  wire w6378;
  wire w6379;
  wire w6380;
  wire w6381;
  wire w6382;
  wire w6383;
  wire w6384;
  wire w6385;
  wire w6386;
  wire w6387;
  wire w6388;
  wire w6389;
  wire w6391;
  wire w6392;
  wire w6393;
  wire w6394;
  wire w6395;
  wire w6396;
  wire w6397;
  wire w6398;
  wire w6399;
  wire w6400;
  wire w6401;
  wire w6402;
  wire w6403;
  wire w6404;
  wire w6405;
  wire w6406;
  wire w6407;
  wire w6408;
  wire w6409;
  wire w6410;
  wire w6411;
  wire w6412;
  wire w6413;
  wire w6414;
  wire w6415;
  wire w6416;
  wire w6417;
  wire w6418;
  wire w6419;
  wire w6420;
  wire w6421;
  wire w6422;
  wire w6423;
  wire w6424;
  wire w6425;
  wire w6426;
  wire w6427;
  wire w6428;
  wire w6429;
  wire w6430;
  wire w6431;
  wire w6432;
  wire w6433;
  wire w6434;
  wire w6435;
  wire w6436;
  wire w6437;
  wire w6438;
  wire w6439;
  wire w6440;
  wire w6441;
  wire w6442;
  wire w6443;
  wire w6444;
  wire w6445;
  wire w6446;
  wire w6447;
  wire w6448;
  wire w6449;
  wire w6450;
  wire w6451;
  wire w6452;
  wire w6453;
  wire w6454;
  wire w6455;
  wire w6456;
  wire w6457;
  wire w6458;
  wire w6459;
  wire w6460;
  wire w6461;
  wire w6462;
  wire w6463;
  wire w6464;
  wire w6465;
  wire w6466;
  wire w6467;
  wire w6468;
  wire w6469;
  wire w6470;
  wire w6471;
  wire w6472;
  wire w6473;
  wire w6474;
  wire w6475;
  wire w6476;
  wire w6477;
  wire w6478;
  wire w6479;
  wire w6480;
  wire w6481;
  wire w6482;
  wire w6483;
  wire w6484;
  wire w6485;
  wire w6486;
  wire w6487;
  wire w6488;
  wire w6489;
  wire w6490;
  wire w6491;
  wire w6492;
  wire w6493;
  wire w6494;
  wire w6495;
  wire w6496;
  wire w6497;
  wire w6498;
  wire w6499;
  wire w6500;
  wire w6501;
  wire w6502;
  wire w6503;
  wire w6505;
  wire w6506;
  wire w6507;
  wire w6508;
  wire w6509;
  wire w6510;
  wire w6511;
  wire w6512;
  wire w6513;
  wire w6514;
  wire w6515;
  wire w6516;
  wire w6517;
  wire w6518;
  wire w6519;
  wire w6520;
  wire w6521;
  wire w6522;
  wire w6523;
  wire w6524;
  wire w6525;
  wire w6526;
  wire w6527;
  wire w6528;
  wire w6529;
  wire w6530;
  wire w6531;
  wire w6532;
  wire w6533;
  wire w6534;
  wire w6535;
  wire w6536;
  wire w6537;
  wire w6538;
  wire w6539;
  wire w6540;
  wire w6541;
  wire w6542;
  wire w6543;
  wire w6544;
  wire w6545;
  wire w6546;
  wire w6547;
  wire w6548;
  wire w6549;
  wire w6550;
  wire w6551;
  wire w6552;
  wire w6553;
  wire w6554;
  wire w6555;
  wire w6556;
  wire w6557;
  wire w6558;
  wire w6559;
  wire w6560;
  wire w6561;
  wire w6562;
  wire w6563;
  wire w6564;
  wire w6565;
  wire w6566;
  wire w6567;
  wire w6568;
  wire w6569;
  wire w6570;
  wire w6571;
  wire w6572;
  wire w6573;
  wire w6574;
  wire w6575;
  wire w6576;
  wire w6577;
  wire w6578;
  wire w6579;
  wire w6580;
  wire w6581;
  wire w6582;
  wire w6583;
  wire w6584;
  wire w6585;
  wire w6586;
  wire w6587;
  wire w6588;
  wire w6589;
  wire w6590;
  wire w6591;
  wire w6592;
  wire w6593;
  wire w6594;
  wire w6595;
  wire w6596;
  wire w6597;
  wire w6598;
  wire w6599;
  wire w6600;
  wire w6601;
  wire w6602;
  wire w6603;
  wire w6604;
  wire w6605;
  wire w6606;
  wire w6607;
  wire w6608;
  wire w6609;
  wire w6610;
  wire w6611;
  wire w6612;
  wire w6613;
  wire w6614;
  wire w6615;
  wire w6616;
  wire w6617;
  wire w6619;
  wire w6620;
  wire w6621;
  wire w6622;
  wire w6623;
  wire w6624;
  wire w6625;
  wire w6626;
  wire w6627;
  wire w6628;
  wire w6629;
  wire w6630;
  wire w6631;
  wire w6632;
  wire w6633;
  wire w6634;
  wire w6635;
  wire w6636;
  wire w6637;
  wire w6638;
  wire w6639;
  wire w6640;
  wire w6641;
  wire w6642;
  wire w6643;
  wire w6644;
  wire w6645;
  wire w6646;
  wire w6647;
  wire w6648;
  wire w6649;
  wire w6650;
  wire w6651;
  wire w6652;
  wire w6653;
  wire w6654;
  wire w6655;
  wire w6656;
  wire w6657;
  wire w6658;
  wire w6659;
  wire w6660;
  wire w6661;
  wire w6662;
  wire w6663;
  wire w6664;
  wire w6665;
  wire w6666;
  wire w6667;
  wire w6668;
  wire w6669;
  wire w6670;
  wire w6671;
  wire w6672;
  wire w6673;
  wire w6674;
  wire w6675;
  wire w6676;
  wire w6677;
  wire w6678;
  wire w6679;
  wire w6680;
  wire w6681;
  wire w6682;
  wire w6683;
  wire w6684;
  wire w6685;
  wire w6686;
  wire w6687;
  wire w6688;
  wire w6689;
  wire w6690;
  wire w6691;
  wire w6692;
  wire w6693;
  wire w6694;
  wire w6695;
  wire w6696;
  wire w6697;
  wire w6698;
  wire w6699;
  wire w6700;
  wire w6701;
  wire w6702;
  wire w6703;
  wire w6704;
  wire w6705;
  wire w6706;
  wire w6707;
  wire w6708;
  wire w6709;
  wire w6710;
  wire w6711;
  wire w6712;
  wire w6713;
  wire w6714;
  wire w6715;
  wire w6716;
  wire w6717;
  wire w6718;
  wire w6719;
  wire w6720;
  wire w6721;
  wire w6722;
  wire w6723;
  wire w6724;
  wire w6725;
  wire w6726;
  wire w6727;
  wire w6728;
  wire w6729;
  wire w6730;
  wire w6731;
  wire w6733;
  wire w6734;
  wire w6735;
  wire w6736;
  wire w6737;
  wire w6738;
  wire w6739;
  wire w6740;
  wire w6741;
  wire w6742;
  wire w6743;
  wire w6744;
  wire w6745;
  wire w6746;
  wire w6747;
  wire w6748;
  wire w6749;
  wire w6750;
  wire w6751;
  wire w6752;
  wire w6753;
  wire w6754;
  wire w6755;
  wire w6756;
  wire w6757;
  wire w6758;
  wire w6759;
  wire w6760;
  wire w6761;
  wire w6762;
  wire w6763;
  wire w6764;
  wire w6765;
  wire w6766;
  wire w6767;
  wire w6768;
  wire w6769;
  wire w6770;
  wire w6771;
  wire w6772;
  wire w6773;
  wire w6774;
  wire w6775;
  wire w6776;
  wire w6777;
  wire w6778;
  wire w6779;
  wire w6780;
  wire w6781;
  wire w6782;
  wire w6783;
  wire w6784;
  wire w6785;
  wire w6786;
  wire w6787;
  wire w6788;
  wire w6789;
  wire w6790;
  wire w6791;
  wire w6792;
  wire w6793;
  wire w6794;
  wire w6795;
  wire w6796;
  wire w6797;
  wire w6798;
  wire w6799;
  wire w6800;
  wire w6801;
  wire w6802;
  wire w6803;
  wire w6804;
  wire w6805;
  wire w6806;
  wire w6807;
  wire w6808;
  wire w6809;
  wire w6810;
  wire w6811;
  wire w6812;
  wire w6813;
  wire w6814;
  wire w6815;
  wire w6816;
  wire w6817;
  wire w6818;
  wire w6819;
  wire w6820;
  wire w6821;
  wire w6822;
  wire w6823;
  wire w6824;
  wire w6825;
  wire w6826;
  wire w6827;
  wire w6828;
  wire w6829;
  wire w6830;
  wire w6831;
  wire w6832;
  wire w6833;
  wire w6834;
  wire w6835;
  wire w6836;
  wire w6837;
  wire w6838;
  wire w6839;
  wire w6840;
  wire w6841;
  wire w6842;
  wire w6843;
  wire w6844;
  wire w6845;
  wire w6847;
  wire w6848;
  wire w6849;
  wire w6850;
  wire w6851;
  wire w6852;
  wire w6853;
  wire w6854;
  wire w6855;
  wire w6856;
  wire w6857;
  wire w6858;
  wire w6859;
  wire w6860;
  wire w6861;
  wire w6862;
  wire w6863;
  wire w6864;
  wire w6865;
  wire w6866;
  wire w6867;
  wire w6868;
  wire w6869;
  wire w6870;
  wire w6871;
  wire w6872;
  wire w6873;
  wire w6874;
  wire w6875;
  wire w6876;
  wire w6877;
  wire w6878;
  wire w6879;
  wire w6880;
  wire w6881;
  wire w6882;
  wire w6883;
  wire w6884;
  wire w6885;
  wire w6886;
  wire w6887;
  wire w6888;
  wire w6889;
  wire w6890;
  wire w6891;
  wire w6892;
  wire w6893;
  wire w6894;
  wire w6895;
  wire w6896;
  wire w6897;
  wire w6898;
  wire w6899;
  wire w6900;
  wire w6901;
  wire w6902;
  wire w6903;
  wire w6904;
  wire w6905;
  wire w6906;
  wire w6907;
  wire w6908;
  wire w6909;
  wire w6910;
  wire w6911;
  wire w6912;
  wire w6913;
  wire w6914;
  wire w6915;
  wire w6916;
  wire w6917;
  wire w6918;
  wire w6919;
  wire w6920;
  wire w6921;
  wire w6922;
  wire w6923;
  wire w6924;
  wire w6925;
  wire w6926;
  wire w6927;
  wire w6928;
  wire w6929;
  wire w6930;
  wire w6931;
  wire w6932;
  wire w6933;
  wire w6934;
  wire w6935;
  wire w6936;
  wire w6937;
  wire w6938;
  wire w6939;
  wire w6940;
  wire w6941;
  wire w6942;
  wire w6943;
  wire w6944;
  wire w6945;
  wire w6946;
  wire w6947;
  wire w6948;
  wire w6949;
  wire w6950;
  wire w6951;
  wire w6952;
  wire w6953;
  wire w6954;
  wire w6955;
  wire w6956;
  wire w6957;
  wire w6958;
  wire w6959;
  wire w6961;
  wire w6962;
  wire w6963;
  wire w6964;
  wire w6965;
  wire w6966;
  wire w6967;
  wire w6968;
  wire w6969;
  wire w6970;
  wire w6971;
  wire w6972;
  wire w6973;
  wire w6974;
  wire w6975;
  wire w6976;
  wire w6977;
  wire w6978;
  wire w6979;
  wire w6980;
  wire w6981;
  wire w6982;
  wire w6983;
  wire w6984;
  wire w6985;
  wire w6986;
  wire w6987;
  wire w6988;
  wire w6989;
  wire w6990;
  wire w6991;
  wire w6992;
  wire w6993;
  wire w6994;
  wire w6995;
  wire w6996;
  wire w6997;
  wire w6998;
  wire w6999;
  wire w7000;
  wire w7001;
  wire w7002;
  wire w7003;
  wire w7004;
  wire w7005;
  wire w7006;
  wire w7007;
  wire w7008;
  wire w7009;
  wire w7010;
  wire w7011;
  wire w7012;
  wire w7013;
  wire w7014;
  wire w7015;
  wire w7016;
  wire w7017;
  wire w7018;
  wire w7019;
  wire w7020;
  wire w7021;
  wire w7022;
  wire w7023;
  wire w7024;
  wire w7025;
  wire w7026;
  wire w7027;
  wire w7028;
  wire w7029;
  wire w7030;
  wire w7031;
  wire w7032;
  wire w7033;
  wire w7034;
  wire w7035;
  wire w7036;
  wire w7037;
  wire w7038;
  wire w7039;
  wire w7040;
  wire w7041;
  wire w7042;
  wire w7043;
  wire w7044;
  wire w7045;
  wire w7046;
  wire w7047;
  wire w7048;
  wire w7049;
  wire w7050;
  wire w7051;
  wire w7052;
  wire w7053;
  wire w7054;
  wire w7055;
  wire w7056;
  wire w7057;
  wire w7058;
  wire w7059;
  wire w7060;
  wire w7061;
  wire w7062;
  wire w7063;
  wire w7064;
  wire w7065;
  wire w7066;
  wire w7067;
  wire w7068;
  wire w7069;
  wire w7070;
  wire w7071;
  wire w7072;
  wire w7073;
  wire w7075;
  wire w7076;
  wire w7077;
  wire w7078;
  wire w7079;
  wire w7080;
  wire w7081;
  wire w7082;
  wire w7083;
  wire w7084;
  wire w7085;
  wire w7086;
  wire w7087;
  wire w7088;
  wire w7089;
  wire w7090;
  wire w7091;
  wire w7092;
  wire w7093;
  wire w7094;
  wire w7095;
  wire w7096;
  wire w7097;
  wire w7098;
  wire w7099;
  wire w7100;
  wire w7101;
  wire w7102;
  wire w7103;
  wire w7104;
  wire w7105;
  wire w7106;
  wire w7107;
  wire w7108;
  wire w7109;
  wire w7110;
  wire w7111;
  wire w7112;
  wire w7113;
  wire w7114;
  wire w7115;
  wire w7116;
  wire w7117;
  wire w7118;
  wire w7119;
  wire w7120;
  wire w7121;
  wire w7122;
  wire w7123;
  wire w7124;
  wire w7125;
  wire w7126;
  wire w7127;
  wire w7128;
  wire w7129;
  wire w7130;
  wire w7131;
  wire w7132;
  wire w7133;
  wire w7134;
  wire w7135;
  wire w7136;
  wire w7137;
  wire w7138;
  wire w7139;
  wire w7140;
  wire w7141;
  wire w7142;
  wire w7143;
  wire w7144;
  wire w7145;
  wire w7146;
  wire w7147;
  wire w7148;
  wire w7149;
  wire w7150;
  wire w7151;
  wire w7152;
  wire w7153;
  wire w7154;
  wire w7155;
  wire w7156;
  wire w7157;
  wire w7158;
  wire w7159;
  wire w7160;
  wire w7161;
  wire w7162;
  wire w7163;
  wire w7164;
  wire w7165;
  wire w7166;
  wire w7167;
  wire w7168;
  wire w7169;
  wire w7170;
  wire w7171;
  wire w7172;
  wire w7173;
  wire w7174;
  wire w7175;
  wire w7176;
  wire w7177;
  wire w7178;
  wire w7179;
  wire w7180;
  wire w7181;
  wire w7182;
  wire w7183;
  wire w7184;
  wire w7185;
  wire w7186;
  wire w7187;
  wire w7189;
  wire w7190;
  wire w7191;
  wire w7192;
  wire w7193;
  wire w7194;
  wire w7195;
  wire w7196;
  wire w7197;
  wire w7198;
  wire w7199;
  wire w7200;
  wire w7201;
  wire w7202;
  wire w7203;
  wire w7204;
  wire w7205;
  wire w7206;
  wire w7207;
  wire w7208;
  wire w7209;
  wire w7210;
  wire w7211;
  wire w7212;
  wire w7213;
  wire w7214;
  wire w7215;
  wire w7216;
  wire w7217;
  wire w7218;
  wire w7219;
  wire w7220;
  wire w7221;
  wire w7222;
  wire w7223;
  wire w7224;
  wire w7225;
  wire w7226;
  wire w7227;
  wire w7228;
  wire w7229;
  wire w7230;
  wire w7231;
  wire w7232;
  wire w7233;
  wire w7234;
  wire w7235;
  wire w7236;
  wire w7237;
  wire w7238;
  wire w7239;
  wire w7240;
  wire w7241;
  wire w7242;
  wire w7243;
  wire w7244;
  wire w7245;
  wire w7246;
  wire w7247;
  wire w7248;
  wire w7249;
  wire w7250;
  wire w7251;
  wire w7252;
  wire w7253;
  wire w7254;
  wire w7255;
  wire w7256;
  wire w7257;
  wire w7258;
  wire w7259;
  wire w7260;
  wire w7261;
  wire w7262;
  wire w7263;
  wire w7264;
  wire w7265;
  wire w7266;
  wire w7267;
  wire w7268;
  wire w7269;
  wire w7270;
  wire w7271;
  wire w7272;
  wire w7273;
  wire w7274;
  wire w7275;
  wire w7276;
  wire w7277;
  wire w7278;
  wire w7279;
  wire w7280;
  wire w7281;
  wire w7282;
  wire w7283;
  wire w7284;
  wire w7285;
  wire w7286;
  wire w7287;
  wire w7288;
  wire w7289;
  wire w7290;
  wire w7291;
  wire w7292;
  wire w7293;
  wire w7294;
  wire w7295;
  wire w7296;
  wire w7297;
  wire w7298;
  wire w7299;
  wire w7300;
  wire w7301;
  wire w7303;
  wire w7304;
  wire w7305;
  wire w7306;
  wire w7307;
  wire w7308;
  wire w7309;
  wire w7310;
  wire w7311;
  wire w7312;
  wire w7313;
  wire w7314;
  wire w7315;
  wire w7316;
  wire w7317;
  wire w7318;
  wire w7319;
  wire w7320;
  wire w7321;
  wire w7322;
  wire w7323;
  wire w7324;
  wire w7325;
  wire w7326;
  wire w7327;
  wire w7328;
  wire w7329;
  wire w7330;
  wire w7331;
  wire w7332;
  wire w7333;
  wire w7334;
  wire w7335;
  wire w7336;
  wire w7337;
  wire w7338;
  wire w7339;
  wire w7340;
  wire w7341;
  wire w7342;
  wire w7343;
  wire w7344;
  wire w7345;
  wire w7346;
  wire w7347;
  wire w7348;
  wire w7349;
  wire w7350;
  wire w7351;
  wire w7352;
  wire w7353;
  wire w7354;
  wire w7355;
  wire w7356;
  wire w7357;
  wire w7358;
  wire w7359;
  wire w7360;
  wire w7361;
  wire w7362;
  wire w7363;
  wire w7364;
  wire w7365;
  wire w7366;
  wire w7367;
  wire w7368;
  wire w7369;
  wire w7370;
  wire w7371;
  wire w7372;
  wire w7373;
  wire w7374;
  wire w7375;
  wire w7376;
  wire w7377;
  wire w7378;
  wire w7379;
  wire w7380;
  wire w7381;
  wire w7382;
  wire w7383;
  wire w7384;
  wire w7385;
  wire w7386;
  wire w7387;
  wire w7388;
  wire w7389;
  wire w7390;
  wire w7391;
  wire w7392;
  wire w7393;
  wire w7394;
  wire w7395;
  wire w7396;
  wire w7397;
  wire w7398;
  wire w7399;
  wire w7400;
  wire w7401;
  wire w7402;
  wire w7403;
  wire w7404;
  wire w7405;
  wire w7406;
  wire w7407;
  wire w7408;
  wire w7409;
  wire w7410;
  wire w7411;
  wire w7412;
  wire w7413;
  wire w7414;
  wire w7415;
  wire w7417;
  wire w7418;
  wire w7419;
  wire w7420;
  wire w7421;
  wire w7422;
  wire w7423;
  wire w7424;
  wire w7425;
  wire w7426;
  wire w7427;
  wire w7428;
  wire w7429;
  wire w7430;
  wire w7431;
  wire w7432;
  wire w7433;
  wire w7434;
  wire w7435;
  wire w7436;
  wire w7437;
  wire w7438;
  wire w7439;
  wire w7440;
  wire w7441;
  wire w7442;
  wire w7443;
  wire w7444;
  wire w7445;
  wire w7446;
  wire w7447;
  wire w7448;
  wire w7449;
  wire w7450;
  wire w7451;
  wire w7452;
  wire w7453;
  wire w7454;
  wire w7455;
  wire w7456;
  wire w7457;
  wire w7458;
  wire w7459;
  wire w7460;
  wire w7461;
  wire w7462;
  wire w7463;
  wire w7464;
  wire w7465;
  wire w7466;
  wire w7467;
  wire w7468;
  wire w7469;
  wire w7470;
  wire w7471;
  wire w7472;
  wire w7473;
  wire w7474;
  wire w7475;
  wire w7476;
  wire w7477;
  wire w7478;
  wire w7479;
  wire w7480;
  wire w7481;
  wire w7482;
  wire w7483;
  wire w7484;
  wire w7485;
  wire w7486;
  wire w7487;
  wire w7488;
  wire w7489;
  wire w7490;
  wire w7491;
  wire w7492;
  wire w7493;
  wire w7494;
  wire w7495;
  wire w7496;
  wire w7497;
  wire w7498;
  wire w7499;
  wire w7500;
  wire w7501;
  wire w7502;
  wire w7503;
  wire w7504;
  wire w7505;
  wire w7506;
  wire w7507;
  wire w7508;
  wire w7509;
  wire w7510;
  wire w7511;
  wire w7512;
  wire w7513;
  wire w7514;
  wire w7515;
  wire w7516;
  wire w7517;
  wire w7518;
  wire w7519;
  wire w7520;
  wire w7521;
  wire w7522;
  wire w7523;
  wire w7524;
  wire w7525;
  wire w7526;
  wire w7527;
  wire w7528;
  wire w7529;
  wire w7531;
  wire w7532;
  wire w7533;
  wire w7534;
  wire w7535;
  wire w7536;
  wire w7537;
  wire w7538;
  wire w7539;
  wire w7540;
  wire w7541;
  wire w7542;
  wire w7543;
  wire w7544;
  wire w7545;
  wire w7546;
  wire w7547;
  wire w7548;
  wire w7549;
  wire w7550;
  wire w7551;
  wire w7552;
  wire w7553;
  wire w7554;
  wire w7555;
  wire w7556;
  wire w7557;
  wire w7558;
  wire w7559;
  wire w7560;
  wire w7561;
  wire w7562;
  wire w7563;
  wire w7564;
  wire w7565;
  wire w7566;
  wire w7567;
  wire w7568;
  wire w7569;
  wire w7570;
  wire w7571;
  wire w7572;
  wire w7573;
  wire w7574;
  wire w7575;
  wire w7576;
  wire w7577;
  wire w7578;
  wire w7579;
  wire w7580;
  wire w7581;
  wire w7582;
  wire w7583;
  wire w7584;
  wire w7585;
  wire w7586;
  wire w7587;
  wire w7588;
  wire w7589;
  wire w7590;
  wire w7591;
  wire w7592;
  wire w7593;
  wire w7594;
  wire w7595;
  wire w7596;
  wire w7597;
  wire w7598;
  wire w7599;
  wire w7600;
  wire w7601;
  wire w7602;
  wire w7603;
  wire w7604;
  wire w7605;
  wire w7606;
  wire w7607;
  wire w7608;
  wire w7609;
  wire w7610;
  wire w7611;
  wire w7612;
  wire w7613;
  wire w7614;
  wire w7615;
  wire w7616;
  wire w7617;
  wire w7618;
  wire w7619;
  wire w7620;
  wire w7621;
  wire w7622;
  wire w7623;
  wire w7624;
  wire w7625;
  wire w7626;
  wire w7627;
  wire w7628;
  wire w7629;
  wire w7630;
  wire w7631;
  wire w7632;
  wire w7633;
  wire w7634;
  wire w7635;
  wire w7636;
  wire w7637;
  wire w7638;
  wire w7639;
  wire w7640;
  wire w7641;
  wire w7642;
  wire w7643;
  wire w7645;
  wire w7646;
  wire w7647;
  wire w7648;
  wire w7649;
  wire w7650;
  wire w7651;
  wire w7652;
  wire w7653;
  wire w7654;
  wire w7655;
  wire w7656;
  wire w7657;
  wire w7658;
  wire w7659;
  wire w7660;
  wire w7661;
  wire w7662;
  wire w7663;
  wire w7664;
  wire w7665;
  wire w7666;
  wire w7667;
  wire w7668;
  wire w7669;
  wire w7670;
  wire w7671;
  wire w7672;
  wire w7673;
  wire w7674;
  wire w7675;
  wire w7676;
  wire w7677;
  wire w7678;
  wire w7679;
  wire w7680;
  wire w7681;
  wire w7682;
  wire w7683;
  wire w7684;
  wire w7685;
  wire w7686;
  wire w7687;
  wire w7688;
  wire w7689;
  wire w7690;
  wire w7691;
  wire w7692;
  wire w7693;
  wire w7694;
  wire w7695;
  wire w7696;
  wire w7697;
  wire w7698;
  wire w7699;
  wire w7700;
  wire w7701;
  wire w7702;
  wire w7703;
  wire w7704;
  wire w7705;
  wire w7706;
  wire w7707;
  wire w7708;
  wire w7709;
  wire w7710;
  wire w7711;
  wire w7712;
  wire w7713;
  wire w7714;
  wire w7715;
  wire w7716;
  wire w7717;
  wire w7718;
  wire w7719;
  wire w7720;
  wire w7721;
  wire w7722;
  wire w7723;
  wire w7724;
  wire w7725;
  wire w7726;
  wire w7727;
  wire w7728;
  wire w7729;
  wire w7730;
  wire w7731;
  wire w7732;
  wire w7733;
  wire w7734;
  wire w7735;
  wire w7736;
  wire w7737;
  wire w7738;
  wire w7739;
  wire w7740;
  wire w7741;
  wire w7742;
  wire w7743;
  wire w7744;
  wire w7745;
  wire w7746;
  wire w7747;
  wire w7748;
  wire w7749;
  wire w7750;
  wire w7751;
  wire w7752;
  wire w7753;
  wire w7754;
  wire w7755;
  wire w7756;
  wire w7757;
  wire w7759;
  wire w7760;
  wire w7761;
  wire w7762;
  wire w7763;
  wire w7764;
  wire w7765;
  wire w7766;
  wire w7767;
  wire w7768;
  wire w7769;
  wire w7770;
  wire w7771;
  wire w7772;
  wire w7773;
  wire w7774;
  wire w7775;
  wire w7776;
  wire w7777;
  wire w7778;
  wire w7779;
  wire w7780;
  wire w7781;
  wire w7782;
  wire w7783;
  wire w7784;
  wire w7785;
  wire w7786;
  wire w7787;
  wire w7788;
  wire w7789;
  wire w7790;
  wire w7791;
  wire w7792;
  wire w7793;
  wire w7794;
  wire w7795;
  wire w7796;
  wire w7797;
  wire w7798;
  wire w7799;
  wire w7800;
  wire w7801;
  wire w7802;
  wire w7803;
  wire w7804;
  wire w7805;
  wire w7806;
  wire w7807;
  wire w7808;
  wire w7809;
  wire w7810;
  wire w7811;
  wire w7812;
  wire w7813;
  wire w7814;
  wire w7815;
  wire w7816;
  wire w7817;
  wire w7818;
  wire w7819;
  wire w7820;
  wire w7821;
  wire w7822;
  wire w7823;
  wire w7824;
  wire w7825;
  wire w7826;
  wire w7827;
  wire w7828;
  wire w7829;
  wire w7830;
  wire w7831;
  wire w7832;
  wire w7833;
  wire w7834;
  wire w7835;
  wire w7836;
  wire w7837;
  wire w7838;
  wire w7839;
  wire w7840;
  wire w7841;
  wire w7842;
  wire w7843;
  wire w7844;
  wire w7845;
  wire w7846;
  wire w7847;
  wire w7848;
  wire w7849;
  wire w7850;
  wire w7851;
  wire w7852;
  wire w7853;
  wire w7854;
  wire w7855;
  wire w7856;
  wire w7857;
  wire w7858;
  wire w7859;
  wire w7860;
  wire w7861;
  wire w7862;
  wire w7863;
  wire w7864;
  wire w7865;
  wire w7866;
  wire w7867;
  wire w7868;
  wire w7869;
  wire w7870;
  wire w7871;
  wire w7873;
  wire w7874;
  wire w7875;
  wire w7876;
  wire w7877;
  wire w7878;
  wire w7879;
  wire w7880;
  wire w7881;
  wire w7882;
  wire w7883;
  wire w7884;
  wire w7885;
  wire w7886;
  wire w7887;
  wire w7888;
  wire w7889;
  wire w7890;
  wire w7891;
  wire w7892;
  wire w7893;
  wire w7894;
  wire w7895;
  wire w7896;
  wire w7897;
  wire w7898;
  wire w7899;
  wire w7900;
  wire w7901;
  wire w7902;
  wire w7903;
  wire w7904;
  wire w7905;
  wire w7906;
  wire w7907;
  wire w7908;
  wire w7909;
  wire w7910;
  wire w7911;
  wire w7912;
  wire w7913;
  wire w7914;
  wire w7915;
  wire w7916;
  wire w7917;
  wire w7918;
  wire w7919;
  wire w7920;
  wire w7921;
  wire w7922;
  wire w7923;
  wire w7924;
  wire w7925;
  wire w7926;
  wire w7927;
  wire w7928;
  wire w7929;
  wire w7930;
  wire w7931;
  wire w7932;
  wire w7933;
  wire w7934;
  wire w7935;
  wire w7936;
  wire w7937;
  wire w7938;
  wire w7939;
  wire w7940;
  wire w7941;
  wire w7942;
  wire w7943;
  wire w7944;
  wire w7945;
  wire w7946;
  wire w7947;
  wire w7948;
  wire w7949;
  wire w7950;
  wire w7951;
  wire w7952;
  wire w7953;
  wire w7954;
  wire w7955;
  wire w7956;
  wire w7957;
  wire w7958;
  wire w7959;
  wire w7960;
  wire w7961;
  wire w7962;
  wire w7963;
  wire w7964;
  wire w7965;
  wire w7966;
  wire w7967;
  wire w7968;
  wire w7969;
  wire w7970;
  wire w7971;
  wire w7972;
  wire w7973;
  wire w7974;
  wire w7975;
  wire w7976;
  wire w7977;
  wire w7978;
  wire w7979;
  wire w7980;
  wire w7981;
  wire w7982;
  wire w7983;
  wire w7984;
  wire w7985;
  wire w7987;
  wire w7988;
  wire w7989;
  wire w7990;
  wire w7991;
  wire w7992;
  wire w7993;
  wire w7994;
  wire w7995;
  wire w7996;
  wire w7997;
  wire w7998;
  wire w7999;
  wire w8000;
  wire w8001;
  wire w8002;
  wire w8003;
  wire w8004;
  wire w8005;
  wire w8006;
  wire w8007;
  wire w8008;
  wire w8009;
  wire w8010;
  wire w8011;
  wire w8012;
  wire w8013;
  wire w8014;
  wire w8015;
  wire w8016;
  wire w8017;
  wire w8018;
  wire w8019;
  wire w8020;
  wire w8021;
  wire w8022;
  wire w8023;
  wire w8024;
  wire w8025;
  wire w8026;
  wire w8027;
  wire w8028;
  wire w8029;
  wire w8030;
  wire w8031;
  wire w8032;
  wire w8033;
  wire w8034;
  wire w8035;
  wire w8036;
  wire w8037;
  wire w8038;
  wire w8039;
  wire w8040;
  wire w8041;
  wire w8042;
  wire w8043;
  wire w8044;
  wire w8045;
  wire w8046;
  wire w8047;
  wire w8048;
  wire w8049;
  wire w8050;
  wire w8051;
  wire w8052;
  wire w8053;
  wire w8054;
  wire w8055;
  wire w8056;
  wire w8057;
  wire w8058;
  wire w8059;
  wire w8060;
  wire w8061;
  wire w8062;
  wire w8063;
  wire w8064;
  wire w8065;
  wire w8066;
  wire w8067;
  wire w8068;
  wire w8069;
  wire w8070;
  wire w8071;
  wire w8072;
  wire w8073;
  wire w8074;
  wire w8075;
  wire w8076;
  wire w8077;
  wire w8078;
  wire w8079;
  wire w8080;
  wire w8081;
  wire w8082;
  wire w8083;
  wire w8084;
  wire w8085;
  wire w8086;
  wire w8087;
  wire w8088;
  wire w8089;
  wire w8090;
  wire w8091;
  wire w8092;
  wire w8093;
  wire w8094;
  wire w8095;
  wire w8096;
  wire w8097;
  wire w8098;
  wire w8099;
  wire w8101;
  wire w8102;
  wire w8103;
  wire w8104;
  wire w8105;
  wire w8106;
  wire w8107;
  wire w8108;
  wire w8109;
  wire w8110;
  wire w8111;
  wire w8112;
  wire w8113;
  wire w8114;
  wire w8115;
  wire w8116;
  wire w8117;
  wire w8118;
  wire w8119;
  wire w8120;
  wire w8121;
  wire w8122;
  wire w8123;
  wire w8124;
  wire w8125;
  wire w8126;
  wire w8127;
  wire w8128;
  wire w8129;
  wire w8130;
  wire w8131;
  wire w8132;
  wire w8133;
  wire w8134;
  wire w8135;
  wire w8136;
  wire w8137;
  wire w8138;
  wire w8139;
  wire w8140;
  wire w8141;
  wire w8142;
  wire w8143;
  wire w8144;
  wire w8145;
  wire w8146;
  wire w8147;
  wire w8148;
  wire w8149;
  wire w8150;
  wire w8151;
  wire w8152;
  wire w8153;
  wire w8154;
  wire w8155;
  wire w8156;
  wire w8157;
  wire w8158;
  wire w8159;
  wire w8160;
  wire w8161;
  wire w8162;
  wire w8163;
  wire w8164;
  wire w8165;
  wire w8166;
  wire w8167;
  wire w8168;
  wire w8169;
  wire w8170;
  wire w8171;
  wire w8172;
  wire w8173;
  wire w8174;
  wire w8175;
  wire w8176;
  wire w8177;
  wire w8178;
  wire w8179;
  wire w8180;
  wire w8181;
  wire w8182;
  wire w8183;
  wire w8184;
  wire w8185;
  wire w8186;
  wire w8187;
  wire w8188;
  wire w8189;
  wire w8190;
  wire w8191;
  wire w8192;
  wire w8193;
  wire w8194;
  wire w8195;
  wire w8196;
  wire w8197;
  wire w8198;
  wire w8199;
  wire w8200;
  wire w8201;
  wire w8202;
  wire w8203;
  wire w8204;
  wire w8205;
  wire w8206;
  wire w8207;
  wire w8208;
  wire w8209;
  wire w8210;
  wire w8211;
  wire w8212;
  wire w8213;
  wire w8215;
  wire w8216;
  wire w8217;
  wire w8218;
  wire w8219;
  wire w8220;
  wire w8221;
  wire w8222;
  wire w8223;
  wire w8224;
  wire w8225;
  wire w8226;
  wire w8227;
  wire w8228;
  wire w8229;
  wire w8230;
  wire w8231;
  wire w8232;
  wire w8233;
  wire w8234;
  wire w8235;
  wire w8236;
  wire w8237;
  wire w8238;
  wire w8239;
  wire w8240;
  wire w8241;
  wire w8242;
  wire w8243;
  wire w8244;
  wire w8245;
  wire w8246;
  wire w8247;
  wire w8248;
  wire w8249;
  wire w8250;
  wire w8251;
  wire w8252;
  wire w8253;
  wire w8254;
  wire w8255;
  wire w8256;
  wire w8257;
  wire w8258;
  wire w8259;
  wire w8260;
  wire w8261;
  wire w8262;
  wire w8263;
  wire w8264;
  wire w8265;
  wire w8266;
  wire w8267;
  wire w8268;
  wire w8269;
  wire w8270;
  wire w8271;
  wire w8272;
  wire w8273;
  wire w8274;
  wire w8275;
  wire w8276;
  wire w8277;
  wire w8278;
  wire w8279;
  wire w8280;
  wire w8281;
  wire w8282;
  wire w8283;
  wire w8284;
  wire w8285;
  wire w8286;
  wire w8287;
  wire w8288;
  wire w8289;
  wire w8290;
  wire w8291;
  wire w8292;
  wire w8293;
  wire w8294;
  wire w8295;
  wire w8296;
  wire w8297;
  wire w8298;
  wire w8299;
  wire w8300;
  wire w8301;
  wire w8302;
  wire w8303;
  wire w8304;
  wire w8305;
  wire w8306;
  wire w8307;
  wire w8308;
  wire w8309;
  wire w8310;
  wire w8311;
  wire w8312;
  wire w8313;
  wire w8314;
  wire w8315;
  wire w8316;
  wire w8317;
  wire w8318;
  wire w8319;
  wire w8320;
  wire w8321;
  wire w8322;
  wire w8323;
  wire w8324;
  wire w8325;
  wire w8326;
  wire w8327;
  wire w8329;
  wire w8330;
  wire w8331;
  wire w8332;
  wire w8333;
  wire w8334;
  wire w8335;
  wire w8336;
  wire w8337;
  wire w8338;
  wire w8339;
  wire w8340;
  wire w8341;
  wire w8342;
  wire w8343;
  wire w8344;
  wire w8345;
  wire w8346;
  wire w8347;
  wire w8348;
  wire w8349;
  wire w8350;
  wire w8351;
  wire w8352;
  wire w8353;
  wire w8354;
  wire w8355;
  wire w8356;
  wire w8357;
  wire w8358;
  wire w8359;
  wire w8360;
  wire w8361;
  wire w8362;
  wire w8363;
  wire w8364;
  wire w8365;
  wire w8366;
  wire w8367;
  wire w8368;
  wire w8369;
  wire w8370;
  wire w8371;
  wire w8372;
  wire w8373;
  wire w8374;
  wire w8375;
  wire w8376;
  wire w8377;
  wire w8378;
  wire w8379;
  wire w8380;
  wire w8381;
  wire w8382;
  wire w8383;
  wire w8384;
  wire w8385;
  wire w8386;
  wire w8387;
  wire w8388;
  wire w8389;
  wire w8390;
  wire w8391;
  wire w8392;
  wire w8393;
  wire w8394;
  wire w8395;
  wire w8396;
  wire w8397;
  wire w8398;
  wire w8399;
  wire w8400;
  wire w8401;
  wire w8402;
  wire w8403;
  wire w8404;
  wire w8405;
  wire w8406;
  wire w8407;
  wire w8408;
  wire w8409;
  wire w8410;
  wire w8411;
  wire w8412;
  wire w8413;
  wire w8414;
  wire w8415;
  wire w8416;
  wire w8417;
  wire w8418;
  wire w8419;
  wire w8420;
  wire w8421;
  wire w8422;
  wire w8423;
  wire w8424;
  wire w8425;
  wire w8426;
  wire w8427;
  wire w8428;
  wire w8429;
  wire w8430;
  wire w8431;
  wire w8432;
  wire w8433;
  wire w8434;
  wire w8435;
  wire w8436;
  wire w8437;
  wire w8438;
  wire w8439;
  wire w8440;
  wire w8441;
  wire w8443;
  wire w8444;
  wire w8445;
  wire w8446;
  wire w8447;
  wire w8448;
  wire w8449;
  wire w8450;
  wire w8451;
  wire w8452;
  wire w8453;
  wire w8454;
  wire w8455;
  wire w8456;
  wire w8457;
  wire w8458;
  wire w8459;
  wire w8460;
  wire w8461;
  wire w8462;
  wire w8463;
  wire w8464;
  wire w8465;
  wire w8466;
  wire w8467;
  wire w8468;
  wire w8469;
  wire w8470;
  wire w8471;
  wire w8472;
  wire w8473;
  wire w8474;
  wire w8475;
  wire w8476;
  wire w8477;
  wire w8478;
  wire w8479;
  wire w8480;
  wire w8481;
  wire w8482;
  wire w8483;
  wire w8484;
  wire w8485;
  wire w8486;
  wire w8487;
  wire w8488;
  wire w8489;
  wire w8490;
  wire w8491;
  wire w8492;
  wire w8493;
  wire w8494;
  wire w8495;
  wire w8496;
  wire w8497;
  wire w8498;
  wire w8499;
  wire w8500;
  wire w8501;
  wire w8502;
  wire w8503;
  wire w8504;
  wire w8505;
  wire w8506;
  wire w8507;
  wire w8508;
  wire w8509;
  wire w8510;
  wire w8511;
  wire w8512;
  wire w8513;
  wire w8514;
  wire w8515;
  wire w8516;
  wire w8517;
  wire w8518;
  wire w8519;
  wire w8520;
  wire w8521;
  wire w8522;
  wire w8523;
  wire w8524;
  wire w8525;
  wire w8526;
  wire w8527;
  wire w8528;
  wire w8529;
  wire w8530;
  wire w8531;
  wire w8532;
  wire w8533;
  wire w8534;
  wire w8535;
  wire w8536;
  wire w8537;
  wire w8538;
  wire w8539;
  wire w8540;
  wire w8541;
  wire w8542;
  wire w8543;
  wire w8544;
  wire w8545;
  wire w8546;
  wire w8547;
  wire w8548;
  wire w8549;
  wire w8550;
  wire w8551;
  wire w8552;
  wire w8553;
  wire w8554;
  wire w8555;
  wire w8557;
  wire w8558;
  wire w8559;
  wire w8560;
  wire w8561;
  wire w8562;
  wire w8563;
  wire w8564;
  wire w8565;
  wire w8566;
  wire w8567;
  wire w8568;
  wire w8569;
  wire w8570;
  wire w8571;
  wire w8572;
  wire w8573;
  wire w8574;
  wire w8575;
  wire w8576;
  wire w8577;
  wire w8578;
  wire w8579;
  wire w8580;
  wire w8581;
  wire w8582;
  wire w8583;
  wire w8584;
  wire w8585;
  wire w8586;
  wire w8587;
  wire w8588;
  wire w8589;
  wire w8590;
  wire w8591;
  wire w8592;
  wire w8593;
  wire w8594;
  wire w8595;
  wire w8596;
  wire w8597;
  wire w8598;
  wire w8599;
  wire w8600;
  wire w8601;
  wire w8602;
  wire w8603;
  wire w8604;
  wire w8605;
  wire w8606;
  wire w8607;
  wire w8608;
  wire w8609;
  wire w8610;
  wire w8611;
  wire w8612;
  wire w8613;
  wire w8614;
  wire w8615;
  wire w8616;
  wire w8617;
  wire w8618;
  wire w8619;
  wire w8620;
  wire w8621;
  wire w8622;
  wire w8623;
  wire w8624;
  wire w8625;
  wire w8626;
  wire w8627;
  wire w8628;
  wire w8629;
  wire w8630;
  wire w8631;
  wire w8632;
  wire w8633;
  wire w8634;
  wire w8635;
  wire w8636;
  wire w8637;
  wire w8638;
  wire w8639;
  wire w8640;
  wire w8641;
  wire w8642;
  wire w8643;
  wire w8644;
  wire w8645;
  wire w8646;
  wire w8647;
  wire w8648;
  wire w8649;
  wire w8650;
  wire w8651;
  wire w8652;
  wire w8653;
  wire w8654;
  wire w8655;
  wire w8656;
  wire w8657;
  wire w8658;
  wire w8659;
  wire w8660;
  wire w8661;
  wire w8662;
  wire w8663;
  wire w8664;
  wire w8665;
  wire w8666;
  wire w8667;
  wire w8668;
  wire w8669;
  wire w8671;
  wire w8672;
  wire w8673;
  wire w8674;
  wire w8675;
  wire w8676;
  wire w8677;
  wire w8678;
  wire w8679;
  wire w8680;
  wire w8681;
  wire w8682;
  wire w8683;
  wire w8684;
  wire w8685;
  wire w8686;
  wire w8687;
  wire w8688;
  wire w8689;
  wire w8690;
  wire w8691;
  wire w8692;
  wire w8693;
  wire w8694;
  wire w8695;
  wire w8696;
  wire w8697;
  wire w8698;
  wire w8699;
  wire w8700;
  wire w8701;
  wire w8702;
  wire w8703;
  wire w8704;
  wire w8705;
  wire w8706;
  wire w8707;
  wire w8708;
  wire w8709;
  wire w8710;
  wire w8711;
  wire w8712;
  wire w8713;
  wire w8714;
  wire w8715;
  wire w8716;
  wire w8717;
  wire w8718;
  wire w8719;
  wire w8720;
  wire w8721;
  wire w8722;
  wire w8723;
  wire w8724;
  wire w8725;
  wire w8726;
  wire w8727;
  wire w8728;
  wire w8729;
  wire w8730;
  wire w8731;
  wire w8732;
  wire w8733;
  wire w8734;
  wire w8735;
  wire w8736;
  wire w8737;
  wire w8738;
  wire w8739;
  wire w8740;
  wire w8741;
  wire w8742;
  wire w8743;
  wire w8744;
  wire w8745;
  wire w8746;
  wire w8747;
  wire w8748;
  wire w8749;
  wire w8750;
  wire w8751;
  wire w8752;
  wire w8753;
  wire w8754;
  wire w8755;
  wire w8756;
  wire w8757;
  wire w8758;
  wire w8759;
  wire w8760;
  wire w8761;
  wire w8762;
  wire w8763;
  wire w8764;
  wire w8765;
  wire w8766;
  wire w8767;
  wire w8768;
  wire w8769;
  wire w8770;
  wire w8771;
  wire w8772;
  wire w8773;
  wire w8774;
  wire w8775;
  wire w8776;
  wire w8777;
  wire w8778;
  wire w8779;
  wire w8780;
  wire w8781;
  wire w8782;
  wire w8783;
  wire w8785;
  wire w8786;
  wire w8787;
  wire w8788;
  wire w8789;
  wire w8790;
  wire w8791;
  wire w8792;
  wire w8793;
  wire w8794;
  wire w8795;
  wire w8796;
  wire w8797;
  wire w8798;
  wire w8799;
  wire w8800;
  wire w8801;
  wire w8802;
  wire w8803;
  wire w8804;
  wire w8805;
  wire w8806;
  wire w8807;
  wire w8808;
  wire w8809;
  wire w8810;
  wire w8811;
  wire w8812;
  wire w8813;
  wire w8814;
  wire w8815;
  wire w8816;
  wire w8817;
  wire w8818;
  wire w8819;
  wire w8820;
  wire w8821;
  wire w8822;
  wire w8823;
  wire w8824;
  wire w8825;
  wire w8826;
  wire w8827;
  wire w8828;
  wire w8829;
  wire w8830;
  wire w8831;
  wire w8832;
  wire w8833;
  wire w8834;
  wire w8835;
  wire w8836;
  wire w8837;
  wire w8838;
  wire w8839;
  wire w8840;
  wire w8841;
  wire w8842;
  wire w8843;
  wire w8844;
  wire w8845;
  wire w8846;
  wire w8847;
  wire w8848;
  wire w8849;
  wire w8850;
  wire w8851;
  wire w8852;
  wire w8853;
  wire w8854;
  wire w8855;
  wire w8856;
  wire w8857;
  wire w8858;
  wire w8859;
  wire w8860;
  wire w8861;
  wire w8862;
  wire w8863;
  wire w8864;
  wire w8865;
  wire w8866;
  wire w8867;
  wire w8868;
  wire w8869;
  wire w8870;
  wire w8871;
  wire w8872;
  wire w8873;
  wire w8874;
  wire w8875;
  wire w8876;
  wire w8877;
  wire w8878;
  wire w8879;
  wire w8880;
  wire w8881;
  wire w8882;
  wire w8883;
  wire w8884;
  wire w8885;
  wire w8886;
  wire w8887;
  wire w8888;
  wire w8889;
  wire w8890;
  wire w8891;
  wire w8892;
  wire w8893;
  wire w8894;
  wire w8895;
  wire w8896;
  wire w8897;
  wire w8899;
  wire w8900;
  wire w8901;
  wire w8902;
  wire w8903;
  wire w8904;
  wire w8905;
  wire w8906;
  wire w8907;
  wire w8908;
  wire w8909;
  wire w8910;
  wire w8911;
  wire w8912;
  wire w8913;
  wire w8914;
  wire w8915;
  wire w8916;
  wire w8917;
  wire w8918;
  wire w8919;
  wire w8920;
  wire w8921;
  wire w8922;
  wire w8923;
  wire w8924;
  wire w8925;
  wire w8926;
  wire w8927;
  wire w8928;
  wire w8929;
  wire w8930;
  wire w8931;
  wire w8932;
  wire w8933;
  wire w8934;
  wire w8935;
  wire w8936;
  wire w8937;
  wire w8938;
  wire w8939;
  wire w8940;
  wire w8941;
  wire w8942;
  wire w8943;
  wire w8944;
  wire w8945;
  wire w8946;
  wire w8947;
  wire w8948;
  wire w8949;
  wire w8950;
  wire w8951;
  wire w8952;
  wire w8953;
  wire w8954;
  wire w8955;
  wire w8956;
  wire w8957;
  wire w8958;
  wire w8959;
  wire w8960;
  wire w8961;
  wire w8962;
  wire w8963;
  wire w8964;
  wire w8965;
  wire w8966;
  wire w8967;
  wire w8968;
  wire w8969;
  wire w8970;
  wire w8971;
  wire w8972;
  wire w8973;
  wire w8974;
  wire w8975;
  wire w8976;
  wire w8977;
  wire w8978;
  wire w8979;
  wire w8980;
  wire w8981;
  wire w8982;
  wire w8983;
  wire w8984;
  wire w8985;
  wire w8986;
  wire w8987;
  wire w8988;
  wire w8989;
  wire w8990;
  wire w8991;
  wire w8992;
  wire w8993;
  wire w8994;
  wire w8995;
  wire w8996;
  wire w8997;
  wire w8998;
  wire w8999;
  wire w9000;
  wire w9001;
  wire w9002;
  wire w9003;
  wire w9004;
  wire w9005;
  wire w9006;
  wire w9007;
  wire w9008;
  wire w9009;
  wire w9010;
  wire w9011;
  wire w9013;
  wire w9014;
  wire w9015;
  wire w9016;
  wire w9017;
  wire w9018;
  wire w9019;
  wire w9020;
  wire w9021;
  wire w9022;
  wire w9023;
  wire w9024;
  wire w9025;
  wire w9026;
  wire w9027;
  wire w9028;
  wire w9029;
  wire w9030;
  wire w9031;
  wire w9032;
  wire w9033;
  wire w9034;
  wire w9035;
  wire w9036;
  wire w9037;
  wire w9038;
  wire w9039;
  wire w9040;
  wire w9041;
  wire w9042;
  wire w9043;
  wire w9044;
  wire w9045;
  wire w9046;
  wire w9047;
  wire w9048;
  wire w9049;
  wire w9050;
  wire w9051;
  wire w9052;
  wire w9053;
  wire w9054;
  wire w9055;
  wire w9056;
  wire w9057;
  wire w9058;
  wire w9059;
  wire w9060;
  wire w9061;
  wire w9062;
  wire w9063;
  wire w9064;
  wire w9065;
  wire w9066;
  wire w9067;
  wire w9068;
  wire w9069;
  wire w9070;
  wire w9071;
  wire w9072;
  wire w9073;
  wire w9074;
  wire w9075;
  wire w9076;
  wire w9077;
  wire w9078;
  wire w9079;
  wire w9080;
  wire w9081;
  wire w9082;
  wire w9083;
  wire w9084;
  wire w9085;
  wire w9086;
  wire w9087;
  wire w9088;
  wire w9089;
  wire w9090;
  wire w9091;
  wire w9092;
  wire w9093;
  wire w9094;
  wire w9095;
  wire w9096;
  wire w9097;
  wire w9098;
  wire w9099;
  wire w9100;
  wire w9101;
  wire w9102;
  wire w9103;
  wire w9104;
  wire w9105;
  wire w9106;
  wire w9107;
  wire w9108;
  wire w9109;
  wire w9110;
  wire w9111;
  wire w9112;
  wire w9113;
  wire w9114;
  wire w9115;
  wire w9116;
  wire w9117;
  wire w9118;
  wire w9119;
  wire w9120;
  wire w9121;
  wire w9122;
  wire w9123;
  wire w9124;
  wire w9125;
  wire w9127;
  wire w9128;
  wire w9129;
  wire w9130;
  wire w9131;
  wire w9132;
  wire w9133;
  wire w9134;
  wire w9135;
  wire w9136;
  wire w9137;
  wire w9138;
  wire w9139;
  wire w9140;
  wire w9141;
  wire w9142;
  wire w9143;
  wire w9144;
  wire w9145;
  wire w9146;
  wire w9147;
  wire w9148;
  wire w9149;
  wire w9150;
  wire w9151;
  wire w9152;
  wire w9153;
  wire w9154;
  wire w9155;
  wire w9156;
  wire w9157;
  wire w9158;
  wire w9159;
  wire w9160;
  wire w9161;
  wire w9162;
  wire w9163;
  wire w9164;
  wire w9165;
  wire w9166;
  wire w9167;
  wire w9168;
  wire w9169;
  wire w9170;
  wire w9171;
  wire w9172;
  wire w9173;
  wire w9174;
  wire w9175;
  wire w9176;
  wire w9177;
  wire w9178;
  wire w9179;
  wire w9180;
  wire w9181;
  wire w9182;
  wire w9183;
  wire w9184;
  wire w9185;
  wire w9186;
  wire w9187;
  wire w9188;
  wire w9189;
  wire w9190;
  wire w9191;
  wire w9192;
  wire w9193;
  wire w9194;
  wire w9195;
  wire w9196;
  wire w9197;
  wire w9198;
  wire w9199;
  wire w9200;
  wire w9201;
  wire w9202;
  wire w9203;
  wire w9204;
  wire w9205;
  wire w9206;
  wire w9207;
  wire w9208;
  wire w9209;
  wire w9210;
  wire w9211;
  wire w9212;
  wire w9213;
  wire w9214;
  wire w9215;
  wire w9216;
  wire w9217;
  wire w9218;
  wire w9219;
  wire w9220;
  wire w9221;
  wire w9222;
  wire w9223;
  wire w9224;
  wire w9225;
  wire w9226;
  wire w9227;
  wire w9228;
  wire w9229;
  wire w9230;
  wire w9231;
  wire w9232;
  wire w9233;
  wire w9234;
  wire w9235;
  wire w9236;
  wire w9237;
  wire w9238;
  wire w9239;
  wire w9241;
  wire w9242;
  wire w9243;
  wire w9244;
  wire w9245;
  wire w9246;
  wire w9247;
  wire w9248;
  wire w9249;
  wire w9250;
  wire w9251;
  wire w9252;
  wire w9253;
  wire w9254;
  wire w9255;
  wire w9256;
  wire w9257;
  wire w9258;
  wire w9259;
  wire w9260;
  wire w9261;
  wire w9262;
  wire w9263;
  wire w9264;
  wire w9265;
  wire w9266;
  wire w9267;
  wire w9268;
  wire w9269;
  wire w9270;
  wire w9271;
  wire w9272;
  wire w9273;
  wire w9274;
  wire w9275;
  wire w9276;
  wire w9277;
  wire w9278;
  wire w9279;
  wire w9280;
  wire w9281;
  wire w9282;
  wire w9283;
  wire w9284;
  wire w9285;
  wire w9286;
  wire w9287;
  wire w9288;
  wire w9289;
  wire w9290;
  wire w9291;
  wire w9292;
  wire w9293;
  wire w9294;
  wire w9295;
  wire w9296;
  wire w9297;
  wire w9298;
  wire w9299;
  wire w9300;
  wire w9301;
  wire w9302;
  wire w9303;
  wire w9304;
  wire w9305;
  wire w9306;
  wire w9307;
  wire w9308;
  wire w9309;
  wire w9310;
  wire w9311;
  wire w9312;
  wire w9313;
  wire w9314;
  wire w9315;
  wire w9316;
  wire w9317;
  wire w9318;
  wire w9319;
  wire w9320;
  wire w9321;
  wire w9322;
  wire w9323;
  wire w9324;
  wire w9325;
  wire w9326;
  wire w9327;
  wire w9328;
  wire w9329;
  wire w9330;
  wire w9331;
  wire w9332;
  wire w9333;
  wire w9334;
  wire w9335;
  wire w9336;
  wire w9337;
  wire w9338;
  wire w9339;
  wire w9340;
  wire w9341;
  wire w9342;
  wire w9343;
  wire w9344;
  wire w9345;
  wire w9346;
  wire w9347;
  wire w9348;
  wire w9349;
  wire w9350;
  wire w9351;
  wire w9352;
  wire w9353;
  wire w9355;
  wire w9356;
  wire w9357;
  wire w9358;
  wire w9359;
  wire w9360;
  wire w9361;
  wire w9362;
  wire w9363;
  wire w9364;
  wire w9365;
  wire w9366;
  wire w9367;
  wire w9368;
  wire w9369;
  wire w9370;
  wire w9371;
  wire w9372;
  wire w9373;
  wire w9374;
  wire w9375;
  wire w9376;
  wire w9377;
  wire w9378;
  wire w9379;
  wire w9380;
  wire w9381;
  wire w9382;
  wire w9383;
  wire w9384;
  wire w9385;
  wire w9386;
  wire w9387;
  wire w9388;
  wire w9389;
  wire w9390;
  wire w9391;
  wire w9392;
  wire w9393;
  wire w9394;
  wire w9395;
  wire w9396;
  wire w9397;
  wire w9398;
  wire w9399;
  wire w9400;
  wire w9401;
  wire w9402;
  wire w9403;
  wire w9404;
  wire w9405;
  wire w9406;
  wire w9407;
  wire w9408;
  wire w9409;
  wire w9410;
  wire w9411;
  wire w9412;
  wire w9413;
  wire w9414;
  wire w9415;
  wire w9416;
  wire w9417;
  wire w9418;
  wire w9419;
  wire w9420;
  wire w9421;
  wire w9422;
  wire w9423;
  wire w9424;
  wire w9425;
  wire w9426;
  wire w9427;
  wire w9428;
  wire w9429;
  wire w9430;
  wire w9431;
  wire w9432;
  wire w9433;
  wire w9434;
  wire w9435;
  wire w9436;
  wire w9437;
  wire w9438;
  wire w9439;
  wire w9440;
  wire w9441;
  wire w9442;
  wire w9443;
  wire w9444;
  wire w9445;
  wire w9446;
  wire w9447;
  wire w9448;
  wire w9449;
  wire w9450;
  wire w9451;
  wire w9452;
  wire w9453;
  wire w9454;
  wire w9455;
  wire w9456;
  wire w9457;
  wire w9458;
  wire w9459;
  wire w9460;
  wire w9461;
  wire w9462;
  wire w9463;
  wire w9464;
  wire w9465;
  wire w9466;
  wire w9467;
  wire w9469;
  wire w9470;
  wire w9471;
  wire w9472;
  wire w9473;
  wire w9474;
  wire w9475;
  wire w9476;
  wire w9477;
  wire w9478;
  wire w9479;
  wire w9480;
  wire w9481;
  wire w9482;
  wire w9483;
  wire w9484;
  wire w9485;
  wire w9486;
  wire w9487;
  wire w9488;
  wire w9489;
  wire w9490;
  wire w9491;
  wire w9492;
  wire w9493;
  wire w9494;
  wire w9495;
  wire w9496;
  wire w9497;
  wire w9498;
  wire w9499;
  wire w9500;
  wire w9501;
  wire w9502;
  wire w9503;
  wire w9504;
  wire w9505;
  wire w9506;
  wire w9507;
  wire w9508;
  wire w9509;
  wire w9510;
  wire w9511;
  wire w9512;
  wire w9513;
  wire w9514;
  wire w9515;
  wire w9516;
  wire w9517;
  wire w9518;
  wire w9519;
  wire w9520;
  wire w9521;
  wire w9522;
  wire w9523;
  wire w9524;
  wire w9525;
  wire w9526;
  wire w9527;
  wire w9528;
  wire w9529;
  wire w9530;
  wire w9531;
  wire w9532;
  wire w9533;
  wire w9534;
  wire w9535;
  wire w9536;
  wire w9537;
  wire w9538;
  wire w9539;
  wire w9540;
  wire w9541;
  wire w9542;
  wire w9543;
  wire w9544;
  wire w9545;
  wire w9546;
  wire w9547;
  wire w9548;
  wire w9549;
  wire w9550;
  wire w9551;
  wire w9552;
  wire w9553;
  wire w9554;
  wire w9555;
  wire w9556;
  wire w9557;
  wire w9558;
  wire w9559;
  wire w9560;
  wire w9561;
  wire w9562;
  wire w9563;
  wire w9564;
  wire w9565;
  wire w9566;
  wire w9567;
  wire w9568;
  wire w9569;
  wire w9570;
  wire w9571;
  wire w9572;
  wire w9573;
  wire w9574;
  wire w9575;
  wire w9576;
  wire w9577;
  wire w9578;
  wire w9579;
  wire w9580;
  wire w9581;
  wire w9583;
  wire w9584;
  wire w9585;
  wire w9586;
  wire w9587;
  wire w9588;
  wire w9589;
  wire w9590;
  wire w9591;
  wire w9592;
  wire w9593;
  wire w9594;
  wire w9595;
  wire w9596;
  wire w9597;
  wire w9598;
  wire w9599;
  wire w9600;
  wire w9601;
  wire w9602;
  wire w9603;
  wire w9604;
  wire w9605;
  wire w9606;
  wire w9607;
  wire w9608;
  wire w9609;
  wire w9610;
  wire w9611;
  wire w9612;
  wire w9613;
  wire w9614;
  wire w9615;
  wire w9616;
  wire w9617;
  wire w9618;
  wire w9619;
  wire w9620;
  wire w9621;
  wire w9622;
  wire w9623;
  wire w9624;
  wire w9625;
  wire w9626;
  wire w9627;
  wire w9628;
  wire w9629;
  wire w9630;
  wire w9631;
  wire w9632;
  wire w9633;
  wire w9634;
  wire w9635;
  wire w9636;
  wire w9637;
  wire w9638;
  wire w9639;
  wire w9640;
  wire w9641;
  wire w9642;
  wire w9643;
  wire w9644;
  wire w9645;
  wire w9646;
  wire w9647;
  wire w9648;
  wire w9649;
  wire w9650;
  wire w9651;
  wire w9652;
  wire w9653;
  wire w9654;
  wire w9655;
  wire w9656;
  wire w9657;
  wire w9658;
  wire w9659;
  wire w9660;
  wire w9661;
  wire w9662;
  wire w9663;
  wire w9664;
  wire w9665;
  wire w9666;
  wire w9667;
  wire w9668;
  wire w9669;
  wire w9670;
  wire w9671;
  wire w9672;
  wire w9673;
  wire w9674;
  wire w9675;
  wire w9676;
  wire w9677;
  wire w9678;
  wire w9679;
  wire w9680;
  wire w9681;
  wire w9682;
  wire w9683;
  wire w9684;
  wire w9685;
  wire w9686;
  wire w9687;
  wire w9688;
  wire w9689;
  wire w9690;
  wire w9691;
  wire w9692;
  wire w9693;
  wire w9694;
  wire w9695;
  wire w9697;
  wire w9698;
  wire w9699;
  wire w9700;
  wire w9701;
  wire w9702;
  wire w9703;
  wire w9704;
  wire w9705;
  wire w9706;
  wire w9707;
  wire w9708;
  wire w9709;
  wire w9710;
  wire w9711;
  wire w9712;
  wire w9713;
  wire w9714;
  wire w9715;
  wire w9716;
  wire w9717;
  wire w9718;
  wire w9719;
  wire w9720;
  wire w9721;
  wire w9722;
  wire w9723;
  wire w9724;
  wire w9725;
  wire w9726;
  wire w9727;
  wire w9728;
  wire w9729;
  wire w9730;
  wire w9731;
  wire w9732;
  wire w9733;
  wire w9734;
  wire w9735;
  wire w9736;
  wire w9737;
  wire w9738;
  wire w9739;
  wire w9740;
  wire w9741;
  wire w9742;
  wire w9743;
  wire w9744;
  wire w9745;
  wire w9746;
  wire w9747;
  wire w9748;
  wire w9749;
  wire w9750;
  wire w9751;
  wire w9752;
  wire w9753;
  wire w9754;
  wire w9755;
  wire w9756;
  wire w9757;
  wire w9758;
  wire w9759;
  wire w9760;
  wire w9761;
  wire w9762;
  wire w9763;
  wire w9764;
  wire w9765;
  wire w9766;
  wire w9767;
  wire w9768;
  wire w9769;
  wire w9770;
  wire w9771;
  wire w9772;
  wire w9773;
  wire w9774;
  wire w9775;
  wire w9776;
  wire w9777;
  wire w9778;
  wire w9779;
  wire w9780;
  wire w9781;
  wire w9782;
  wire w9783;
  wire w9784;
  wire w9785;
  wire w9786;
  wire w9787;
  wire w9788;
  wire w9789;
  wire w9790;
  wire w9791;
  wire w9792;
  wire w9793;
  wire w9794;
  wire w9795;
  wire w9796;
  wire w9797;
  wire w9798;
  wire w9799;
  wire w9800;
  wire w9801;
  wire w9802;
  wire w9803;
  wire w9804;
  wire w9805;
  wire w9806;
  wire w9807;
  wire w9808;
  wire w9809;
  wire w9811;
  wire w9812;
  wire w9813;
  wire w9814;
  wire w9815;
  wire w9816;
  wire w9817;
  wire w9818;
  wire w9819;
  wire w9820;
  wire w9821;
  wire w9822;
  wire w9823;
  wire w9824;
  wire w9825;
  wire w9826;
  wire w9827;
  wire w9828;
  wire w9829;
  wire w9830;
  wire w9831;
  wire w9832;
  wire w9833;
  wire w9834;
  wire w9835;
  wire w9836;
  wire w9837;
  wire w9838;
  wire w9839;
  wire w9840;
  wire w9841;
  wire w9842;
  wire w9843;
  wire w9844;
  wire w9845;
  wire w9846;
  wire w9847;
  wire w9848;
  wire w9849;
  wire w9850;
  wire w9851;
  wire w9852;
  wire w9853;
  wire w9854;
  wire w9855;
  wire w9856;
  wire w9857;
  wire w9858;
  wire w9859;
  wire w9860;
  wire w9861;
  wire w9862;
  wire w9863;
  wire w9864;
  wire w9865;
  wire w9866;
  wire w9867;
  wire w9868;
  wire w9869;
  wire w9870;
  wire w9871;
  wire w9872;
  wire w9873;
  wire w9874;
  wire w9875;
  wire w9876;
  wire w9877;
  wire w9878;
  wire w9879;
  wire w9880;
  wire w9881;
  wire w9882;
  wire w9883;
  wire w9884;
  wire w9885;
  wire w9886;
  wire w9887;
  wire w9888;
  wire w9889;
  wire w9890;
  wire w9891;
  wire w9892;
  wire w9893;
  wire w9894;
  wire w9895;
  wire w9896;
  wire w9897;
  wire w9898;
  wire w9899;
  wire w9900;
  wire w9901;
  wire w9902;
  wire w9903;
  wire w9904;
  wire w9905;
  wire w9906;
  wire w9907;
  wire w9908;
  wire w9909;
  wire w9910;
  wire w9911;
  wire w9912;
  wire w9913;
  wire w9914;
  wire w9915;
  wire w9916;
  wire w9917;
  wire w9918;
  wire w9919;
  wire w9920;
  wire w9921;
  wire w9922;
  wire w9923;
  wire w9925;
  wire w9926;
  wire w9927;
  wire w9928;
  wire w9929;
  wire w9930;
  wire w9931;
  wire w9932;
  wire w9933;
  wire w9934;
  wire w9935;
  wire w9936;
  wire w9937;
  wire w9938;
  wire w9939;
  wire w9940;
  wire w9941;
  wire w9942;
  wire w9943;
  wire w9944;
  wire w9945;
  wire w9946;
  wire w9947;
  wire w9948;
  wire w9949;
  wire w9950;
  wire w9951;
  wire w9952;
  wire w9953;
  wire w9954;
  wire w9955;
  wire w9956;
  wire w9957;
  wire w9958;
  wire w9959;
  wire w9960;
  wire w9961;
  wire w9962;
  wire w9963;
  wire w9964;
  wire w9965;
  wire w9966;
  wire w9967;
  wire w9968;
  wire w9969;
  wire w9970;
  wire w9971;
  wire w9972;
  wire w9973;
  wire w9974;
  wire w9975;
  wire w9976;
  wire w9977;
  wire w9978;
  wire w9979;
  wire w9980;
  wire w9981;
  wire w9982;
  wire w9983;
  wire w9984;
  wire w9985;
  wire w9986;
  wire w9987;
  wire w9988;
  wire w9989;
  wire w9990;
  wire w9991;
  wire w9992;
  wire w9993;
  wire w9994;
  wire w9995;
  wire w9996;
  wire w9997;
  wire w9998;
  wire w9999;
  wire w10000;
  wire w10001;
  wire w10002;
  wire w10003;
  wire w10004;
  wire w10005;
  wire w10006;
  wire w10007;
  wire w10008;
  wire w10009;
  wire w10010;
  wire w10011;
  wire w10012;
  wire w10013;
  wire w10014;
  wire w10015;
  wire w10016;
  wire w10017;
  wire w10018;
  wire w10019;
  wire w10020;
  wire w10021;
  wire w10022;
  wire w10023;
  wire w10024;
  wire w10025;
  wire w10026;
  wire w10027;
  wire w10028;
  wire w10029;
  wire w10030;
  wire w10031;
  wire w10032;
  wire w10033;
  wire w10034;
  wire w10035;
  wire w10036;
  wire w10037;
  wire w10039;
  wire w10040;
  wire w10041;
  wire w10042;
  wire w10043;
  wire w10044;
  wire w10045;
  wire w10046;
  wire w10047;
  wire w10048;
  wire w10049;
  wire w10050;
  wire w10051;
  wire w10052;
  wire w10053;
  wire w10054;
  wire w10055;
  wire w10056;
  wire w10057;
  wire w10058;
  wire w10059;
  wire w10060;
  wire w10061;
  wire w10062;
  wire w10063;
  wire w10064;
  wire w10065;
  wire w10066;
  wire w10067;
  wire w10068;
  wire w10069;
  wire w10070;
  wire w10071;
  wire w10072;
  wire w10073;
  wire w10074;
  wire w10075;
  wire w10076;
  wire w10077;
  wire w10078;
  wire w10079;
  wire w10080;
  wire w10081;
  wire w10082;
  wire w10083;
  wire w10084;
  wire w10085;
  wire w10086;
  wire w10087;
  wire w10088;
  wire w10089;
  wire w10090;
  wire w10091;
  wire w10092;
  wire w10093;
  wire w10094;
  wire w10095;
  wire w10096;
  wire w10097;
  wire w10098;
  wire w10099;
  wire w10100;
  wire w10101;
  wire w10102;
  wire w10103;
  wire w10104;
  wire w10105;
  wire w10106;
  wire w10107;
  wire w10108;
  wire w10109;
  wire w10110;
  wire w10111;
  wire w10112;
  wire w10113;
  wire w10114;
  wire w10115;
  wire w10116;
  wire w10117;
  wire w10118;
  wire w10119;
  wire w10120;
  wire w10121;
  wire w10122;
  wire w10123;
  wire w10124;
  wire w10125;
  wire w10126;
  wire w10127;
  wire w10128;
  wire w10129;
  wire w10130;
  wire w10131;
  wire w10132;
  wire w10133;
  wire w10134;
  wire w10135;
  wire w10136;
  wire w10137;
  wire w10138;
  wire w10139;
  wire w10140;
  wire w10141;
  wire w10142;
  wire w10143;
  wire w10144;
  wire w10145;
  wire w10146;
  wire w10147;
  wire w10148;
  wire w10149;
  wire w10150;
  wire w10151;
  wire w10153;
  wire w10154;
  wire w10155;
  wire w10156;
  wire w10157;
  wire w10158;
  wire w10159;
  wire w10160;
  wire w10161;
  wire w10162;
  wire w10163;
  wire w10164;
  wire w10165;
  wire w10166;
  wire w10167;
  wire w10168;
  wire w10169;
  wire w10170;
  wire w10171;
  wire w10172;
  wire w10173;
  wire w10174;
  wire w10175;
  wire w10176;
  wire w10177;
  wire w10178;
  wire w10179;
  wire w10180;
  wire w10181;
  wire w10182;
  wire w10183;
  wire w10184;
  wire w10185;
  wire w10186;
  wire w10187;
  wire w10188;
  wire w10189;
  wire w10190;
  wire w10191;
  wire w10192;
  wire w10193;
  wire w10194;
  wire w10195;
  wire w10196;
  wire w10197;
  wire w10198;
  wire w10199;
  wire w10200;
  wire w10201;
  wire w10202;
  wire w10203;
  wire w10204;
  wire w10205;
  wire w10206;
  wire w10207;
  wire w10208;
  wire w10209;
  wire w10210;
  wire w10211;
  wire w10212;
  wire w10213;
  wire w10214;
  wire w10215;
  wire w10216;
  wire w10217;
  wire w10218;
  wire w10219;
  wire w10220;
  wire w10221;
  wire w10222;
  wire w10223;
  wire w10224;
  wire w10225;
  wire w10226;
  wire w10227;
  wire w10228;
  wire w10229;
  wire w10230;
  wire w10231;
  wire w10232;
  wire w10233;
  wire w10234;
  wire w10235;
  wire w10236;
  wire w10237;
  wire w10238;
  wire w10239;
  wire w10240;
  wire w10241;
  wire w10242;
  wire w10243;
  wire w10244;
  wire w10245;
  wire w10246;
  wire w10247;
  wire w10248;
  wire w10249;
  wire w10250;
  wire w10251;
  wire w10252;
  wire w10253;
  wire w10254;
  wire w10255;
  wire w10256;
  wire w10257;
  wire w10258;
  wire w10259;
  wire w10260;
  wire w10261;
  wire w10262;
  wire w10263;
  wire w10264;
  wire w10265;
  wire w10267;
  wire w10268;
  wire w10269;
  wire w10270;
  wire w10271;
  wire w10272;
  wire w10273;
  wire w10274;
  wire w10275;
  wire w10276;
  wire w10277;
  wire w10278;
  wire w10279;
  wire w10280;
  wire w10281;
  wire w10282;
  wire w10283;
  wire w10284;
  wire w10285;
  wire w10286;
  wire w10287;
  wire w10288;
  wire w10289;
  wire w10290;
  wire w10291;
  wire w10292;
  wire w10293;
  wire w10294;
  wire w10295;
  wire w10296;
  wire w10297;
  wire w10298;
  wire w10299;
  wire w10300;
  wire w10301;
  wire w10302;
  wire w10303;
  wire w10304;
  wire w10305;
  wire w10306;
  wire w10307;
  wire w10308;
  wire w10309;
  wire w10310;
  wire w10311;
  wire w10312;
  wire w10313;
  wire w10314;
  wire w10315;
  wire w10316;
  wire w10317;
  wire w10318;
  wire w10319;
  wire w10320;
  wire w10321;
  wire w10322;
  wire w10323;
  wire w10324;
  wire w10325;
  wire w10326;
  wire w10327;
  wire w10328;
  wire w10329;
  wire w10330;
  wire w10331;
  wire w10332;
  wire w10333;
  wire w10334;
  wire w10335;
  wire w10336;
  wire w10337;
  wire w10338;
  wire w10339;
  wire w10340;
  wire w10341;
  wire w10342;
  wire w10343;
  wire w10344;
  wire w10345;
  wire w10346;
  wire w10347;
  wire w10348;
  wire w10349;
  wire w10350;
  wire w10351;
  wire w10352;
  wire w10353;
  wire w10354;
  wire w10355;
  wire w10356;
  wire w10357;
  wire w10358;
  wire w10359;
  wire w10360;
  wire w10361;
  wire w10362;
  wire w10363;
  wire w10364;
  wire w10365;
  wire w10366;
  wire w10367;
  wire w10368;
  wire w10369;
  wire w10370;
  wire w10371;
  wire w10372;
  wire w10373;
  wire w10374;
  wire w10375;
  wire w10376;
  wire w10377;
  wire w10378;
  wire w10379;
  wire w10381;
  wire w10382;
  wire w10383;
  wire w10384;
  wire w10385;
  wire w10386;
  wire w10387;
  wire w10388;
  wire w10389;
  wire w10390;
  wire w10391;
  wire w10392;
  wire w10393;
  wire w10394;
  wire w10395;
  wire w10396;
  wire w10397;
  wire w10398;
  wire w10399;
  wire w10400;
  wire w10401;
  wire w10402;
  wire w10403;
  wire w10404;
  wire w10405;
  wire w10406;
  wire w10407;
  wire w10408;
  wire w10409;
  wire w10410;
  wire w10411;
  wire w10412;
  wire w10413;
  wire w10414;
  wire w10415;
  wire w10416;
  wire w10417;
  wire w10418;
  wire w10419;
  wire w10420;
  wire w10421;
  wire w10422;
  wire w10423;
  wire w10424;
  wire w10425;
  wire w10426;
  wire w10427;
  wire w10428;
  wire w10429;
  wire w10430;
  wire w10431;
  wire w10432;
  wire w10433;
  wire w10434;
  wire w10435;
  wire w10436;
  wire w10437;
  wire w10438;
  wire w10439;
  wire w10440;
  wire w10441;
  wire w10442;
  wire w10443;
  wire w10444;
  wire w10445;
  wire w10446;
  wire w10447;
  wire w10448;
  wire w10449;
  wire w10450;
  wire w10451;
  wire w10452;
  wire w10453;
  wire w10454;
  wire w10455;
  wire w10456;
  wire w10457;
  wire w10458;
  wire w10459;
  wire w10460;
  wire w10461;
  wire w10462;
  wire w10463;
  wire w10464;
  wire w10465;
  wire w10466;
  wire w10467;
  wire w10468;
  wire w10469;
  wire w10470;
  wire w10471;
  wire w10472;
  wire w10473;
  wire w10474;
  wire w10475;
  wire w10476;
  wire w10477;
  wire w10478;
  wire w10479;
  wire w10480;
  wire w10481;
  wire w10482;
  wire w10483;
  wire w10484;
  wire w10485;
  wire w10486;
  wire w10487;
  wire w10488;
  wire w10489;
  wire w10490;
  wire w10491;
  wire w10492;
  wire w10493;
  wire w10495;
  wire w10496;
  wire w10497;
  wire w10498;
  wire w10499;
  wire w10500;
  wire w10501;
  wire w10502;
  wire w10503;
  wire w10504;
  wire w10505;
  wire w10506;
  wire w10507;
  wire w10508;
  wire w10509;
  wire w10510;
  wire w10511;
  wire w10512;
  wire w10513;
  wire w10514;
  wire w10515;
  wire w10516;
  wire w10517;
  wire w10518;
  wire w10519;
  wire w10520;
  wire w10521;
  wire w10522;
  wire w10523;
  wire w10524;
  wire w10525;
  wire w10526;
  wire w10527;
  wire w10528;
  wire w10529;
  wire w10530;
  wire w10531;
  wire w10532;
  wire w10533;
  wire w10534;
  wire w10535;
  wire w10536;
  wire w10537;
  wire w10538;
  wire w10539;
  wire w10540;
  wire w10541;
  wire w10542;
  wire w10543;
  wire w10544;
  wire w10545;
  wire w10546;
  wire w10547;
  wire w10548;
  wire w10549;
  wire w10550;
  wire w10551;
  wire w10552;
  wire w10553;
  wire w10554;
  wire w10555;
  wire w10556;
  wire w10557;
  wire w10558;
  wire w10559;
  wire w10560;
  wire w10561;
  wire w10562;
  wire w10563;
  wire w10564;
  wire w10565;
  wire w10566;
  wire w10567;
  wire w10568;
  wire w10569;
  wire w10570;
  wire w10571;
  wire w10572;
  wire w10573;
  wire w10574;
  wire w10575;
  wire w10576;
  wire w10577;
  wire w10578;
  wire w10579;
  wire w10580;
  wire w10581;
  wire w10582;
  wire w10583;
  wire w10584;
  wire w10585;
  wire w10586;
  wire w10587;
  wire w10588;
  wire w10589;
  wire w10590;
  wire w10591;
  wire w10592;
  wire w10593;
  wire w10594;
  wire w10595;
  wire w10596;
  wire w10597;
  wire w10598;
  wire w10599;
  wire w10600;
  wire w10601;
  wire w10602;
  wire w10603;
  wire w10604;
  wire w10605;
  wire w10606;
  wire w10607;
  wire w10609;
  wire w10611;
  wire w10613;
  wire w10615;
  wire w10617;
  wire w10619;
  wire w10621;
  wire w10623;
  wire w10625;
  wire w10627;
  wire w10629;
  wire w10631;
  wire w10633;
  wire w10635;
  wire w10637;
  wire w10639;
  wire w10641;
  wire w10643;
  wire w10645;
  wire w10647;
  wire w10649;
  wire w10651;
  wire w10653;
  wire w10655;
  wire w10657;
  wire w10659;
  wire w10661;
  wire w10663;
  wire w10665;
  wire w10667;
  wire w10669;
  wire w10671;
  wire w10673;
  wire w10675;
  wire w10677;
  wire w10679;
  wire w10681;
  wire w10683;
  wire w10685;
  wire w10687;
  wire w10689;
  wire w10691;
  wire w10693;
  wire w10695;
  wire w10697;
  wire w10699;
  wire w10701;
  wire w10703;
  wire w10705;
  wire w10707;
  wire w10709;
  wire w10711;
  wire w10713;
  wire w10715;
  wire w10717;
  wire w10719;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w3655);
  FullAdder U1 (w3655, IN2[0], IN2[1], w3656, w3657);
  FullAdder U2 (w3657, IN3[0], IN3[1], w3658, w3659);
  FullAdder U3 (w3659, IN4[0], IN4[1], w3660, w3661);
  FullAdder U4 (w3661, IN5[0], IN5[1], w3662, w3663);
  FullAdder U5 (w3663, IN6[0], IN6[1], w3664, w3665);
  FullAdder U6 (w3665, IN7[0], IN7[1], w3666, w3667);
  FullAdder U7 (w3667, IN8[0], IN8[1], w3668, w3669);
  FullAdder U8 (w3669, IN9[0], IN9[1], w3670, w3671);
  FullAdder U9 (w3671, IN10[0], IN10[1], w3672, w3673);
  FullAdder U10 (w3673, IN11[0], IN11[1], w3674, w3675);
  FullAdder U11 (w3675, IN12[0], IN12[1], w3676, w3677);
  FullAdder U12 (w3677, IN13[0], IN13[1], w3678, w3679);
  FullAdder U13 (w3679, IN14[0], IN14[1], w3680, w3681);
  FullAdder U14 (w3681, IN15[0], IN15[1], w3682, w3683);
  FullAdder U15 (w3683, IN16[0], IN16[1], w3684, w3685);
  FullAdder U16 (w3685, IN17[0], IN17[1], w3686, w3687);
  FullAdder U17 (w3687, IN18[0], IN18[1], w3688, w3689);
  FullAdder U18 (w3689, IN19[0], IN19[1], w3690, w3691);
  FullAdder U19 (w3691, IN20[0], IN20[1], w3692, w3693);
  FullAdder U20 (w3693, IN21[0], IN21[1], w3694, w3695);
  FullAdder U21 (w3695, IN22[0], IN22[1], w3696, w3697);
  FullAdder U22 (w3697, IN23[0], IN23[1], w3698, w3699);
  FullAdder U23 (w3699, IN24[0], IN24[1], w3700, w3701);
  FullAdder U24 (w3701, IN25[0], IN25[1], w3702, w3703);
  FullAdder U25 (w3703, IN26[0], IN26[1], w3704, w3705);
  FullAdder U26 (w3705, IN27[0], IN27[1], w3706, w3707);
  FullAdder U27 (w3707, IN28[0], IN28[1], w3708, w3709);
  FullAdder U28 (w3709, IN29[0], IN29[1], w3710, w3711);
  FullAdder U29 (w3711, IN30[0], IN30[1], w3712, w3713);
  FullAdder U30 (w3713, IN31[0], IN31[1], w3714, w3715);
  FullAdder U31 (w3715, IN32[0], IN32[1], w3716, w3717);
  FullAdder U32 (w3717, IN33[0], IN33[1], w3718, w3719);
  FullAdder U33 (w3719, IN34[0], IN34[1], w3720, w3721);
  FullAdder U34 (w3721, IN35[0], IN35[1], w3722, w3723);
  FullAdder U35 (w3723, IN36[0], IN36[1], w3724, w3725);
  FullAdder U36 (w3725, IN37[0], IN37[1], w3726, w3727);
  FullAdder U37 (w3727, IN38[0], IN38[1], w3728, w3729);
  FullAdder U38 (w3729, IN39[0], IN39[1], w3730, w3731);
  FullAdder U39 (w3731, IN40[0], IN40[1], w3732, w3733);
  FullAdder U40 (w3733, IN41[0], IN41[1], w3734, w3735);
  FullAdder U41 (w3735, IN42[0], IN42[1], w3736, w3737);
  FullAdder U42 (w3737, IN43[0], IN43[1], w3738, w3739);
  FullAdder U43 (w3739, IN44[0], IN44[1], w3740, w3741);
  FullAdder U44 (w3741, IN45[0], IN45[1], w3742, w3743);
  FullAdder U45 (w3743, IN46[0], IN46[1], w3744, w3745);
  FullAdder U46 (w3745, IN47[0], IN47[1], w3746, w3747);
  FullAdder U47 (w3747, IN48[0], IN48[1], w3748, w3749);
  FullAdder U48 (w3749, IN49[0], IN49[1], w3750, w3751);
  FullAdder U49 (w3751, IN50[0], IN50[1], w3752, w3753);
  FullAdder U50 (w3753, IN51[0], IN51[1], w3754, w3755);
  FullAdder U51 (w3755, IN52[0], IN52[1], w3756, w3757);
  FullAdder U52 (w3757, IN53[0], IN53[1], w3758, w3759);
  FullAdder U53 (w3759, IN54[0], IN54[1], w3760, w3761);
  FullAdder U54 (w3761, IN55[0], IN55[1], w3762, w3763);
  FullAdder U55 (w3763, IN56[0], IN56[1], w3764, w3765);
  FullAdder U56 (w3765, IN57[0], IN57[1], w3766, w3767);
  HalfAdder U57 (w3656, IN2[2], Out1[2], w3769);
  FullAdder U58 (w3769, w3658, IN3[2], w3770, w3771);
  FullAdder U59 (w3771, w3660, IN4[2], w3772, w3773);
  FullAdder U60 (w3773, w3662, IN5[2], w3774, w3775);
  FullAdder U61 (w3775, w3664, IN6[2], w3776, w3777);
  FullAdder U62 (w3777, w3666, IN7[2], w3778, w3779);
  FullAdder U63 (w3779, w3668, IN8[2], w3780, w3781);
  FullAdder U64 (w3781, w3670, IN9[2], w3782, w3783);
  FullAdder U65 (w3783, w3672, IN10[2], w3784, w3785);
  FullAdder U66 (w3785, w3674, IN11[2], w3786, w3787);
  FullAdder U67 (w3787, w3676, IN12[2], w3788, w3789);
  FullAdder U68 (w3789, w3678, IN13[2], w3790, w3791);
  FullAdder U69 (w3791, w3680, IN14[2], w3792, w3793);
  FullAdder U70 (w3793, w3682, IN15[2], w3794, w3795);
  FullAdder U71 (w3795, w3684, IN16[2], w3796, w3797);
  FullAdder U72 (w3797, w3686, IN17[2], w3798, w3799);
  FullAdder U73 (w3799, w3688, IN18[2], w3800, w3801);
  FullAdder U74 (w3801, w3690, IN19[2], w3802, w3803);
  FullAdder U75 (w3803, w3692, IN20[2], w3804, w3805);
  FullAdder U76 (w3805, w3694, IN21[2], w3806, w3807);
  FullAdder U77 (w3807, w3696, IN22[2], w3808, w3809);
  FullAdder U78 (w3809, w3698, IN23[2], w3810, w3811);
  FullAdder U79 (w3811, w3700, IN24[2], w3812, w3813);
  FullAdder U80 (w3813, w3702, IN25[2], w3814, w3815);
  FullAdder U81 (w3815, w3704, IN26[2], w3816, w3817);
  FullAdder U82 (w3817, w3706, IN27[2], w3818, w3819);
  FullAdder U83 (w3819, w3708, IN28[2], w3820, w3821);
  FullAdder U84 (w3821, w3710, IN29[2], w3822, w3823);
  FullAdder U85 (w3823, w3712, IN30[2], w3824, w3825);
  FullAdder U86 (w3825, w3714, IN31[2], w3826, w3827);
  FullAdder U87 (w3827, w3716, IN32[2], w3828, w3829);
  FullAdder U88 (w3829, w3718, IN33[2], w3830, w3831);
  FullAdder U89 (w3831, w3720, IN34[2], w3832, w3833);
  FullAdder U90 (w3833, w3722, IN35[2], w3834, w3835);
  FullAdder U91 (w3835, w3724, IN36[2], w3836, w3837);
  FullAdder U92 (w3837, w3726, IN37[2], w3838, w3839);
  FullAdder U93 (w3839, w3728, IN38[2], w3840, w3841);
  FullAdder U94 (w3841, w3730, IN39[2], w3842, w3843);
  FullAdder U95 (w3843, w3732, IN40[2], w3844, w3845);
  FullAdder U96 (w3845, w3734, IN41[2], w3846, w3847);
  FullAdder U97 (w3847, w3736, IN42[2], w3848, w3849);
  FullAdder U98 (w3849, w3738, IN43[2], w3850, w3851);
  FullAdder U99 (w3851, w3740, IN44[2], w3852, w3853);
  FullAdder U100 (w3853, w3742, IN45[2], w3854, w3855);
  FullAdder U101 (w3855, w3744, IN46[2], w3856, w3857);
  FullAdder U102 (w3857, w3746, IN47[2], w3858, w3859);
  FullAdder U103 (w3859, w3748, IN48[2], w3860, w3861);
  FullAdder U104 (w3861, w3750, IN49[2], w3862, w3863);
  FullAdder U105 (w3863, w3752, IN50[2], w3864, w3865);
  FullAdder U106 (w3865, w3754, IN51[2], w3866, w3867);
  FullAdder U107 (w3867, w3756, IN52[2], w3868, w3869);
  FullAdder U108 (w3869, w3758, IN53[2], w3870, w3871);
  FullAdder U109 (w3871, w3760, IN54[2], w3872, w3873);
  FullAdder U110 (w3873, w3762, IN55[2], w3874, w3875);
  FullAdder U111 (w3875, w3764, IN56[2], w3876, w3877);
  FullAdder U112 (w3877, w3766, IN57[2], w3878, w3879);
  FullAdder U113 (w3879, w3767, IN58[0], w3880, w3881);
  HalfAdder U114 (w3770, IN3[3], Out1[3], w3883);
  FullAdder U115 (w3883, w3772, IN4[3], w3884, w3885);
  FullAdder U116 (w3885, w3774, IN5[3], w3886, w3887);
  FullAdder U117 (w3887, w3776, IN6[3], w3888, w3889);
  FullAdder U118 (w3889, w3778, IN7[3], w3890, w3891);
  FullAdder U119 (w3891, w3780, IN8[3], w3892, w3893);
  FullAdder U120 (w3893, w3782, IN9[3], w3894, w3895);
  FullAdder U121 (w3895, w3784, IN10[3], w3896, w3897);
  FullAdder U122 (w3897, w3786, IN11[3], w3898, w3899);
  FullAdder U123 (w3899, w3788, IN12[3], w3900, w3901);
  FullAdder U124 (w3901, w3790, IN13[3], w3902, w3903);
  FullAdder U125 (w3903, w3792, IN14[3], w3904, w3905);
  FullAdder U126 (w3905, w3794, IN15[3], w3906, w3907);
  FullAdder U127 (w3907, w3796, IN16[3], w3908, w3909);
  FullAdder U128 (w3909, w3798, IN17[3], w3910, w3911);
  FullAdder U129 (w3911, w3800, IN18[3], w3912, w3913);
  FullAdder U130 (w3913, w3802, IN19[3], w3914, w3915);
  FullAdder U131 (w3915, w3804, IN20[3], w3916, w3917);
  FullAdder U132 (w3917, w3806, IN21[3], w3918, w3919);
  FullAdder U133 (w3919, w3808, IN22[3], w3920, w3921);
  FullAdder U134 (w3921, w3810, IN23[3], w3922, w3923);
  FullAdder U135 (w3923, w3812, IN24[3], w3924, w3925);
  FullAdder U136 (w3925, w3814, IN25[3], w3926, w3927);
  FullAdder U137 (w3927, w3816, IN26[3], w3928, w3929);
  FullAdder U138 (w3929, w3818, IN27[3], w3930, w3931);
  FullAdder U139 (w3931, w3820, IN28[3], w3932, w3933);
  FullAdder U140 (w3933, w3822, IN29[3], w3934, w3935);
  FullAdder U141 (w3935, w3824, IN30[3], w3936, w3937);
  FullAdder U142 (w3937, w3826, IN31[3], w3938, w3939);
  FullAdder U143 (w3939, w3828, IN32[3], w3940, w3941);
  FullAdder U144 (w3941, w3830, IN33[3], w3942, w3943);
  FullAdder U145 (w3943, w3832, IN34[3], w3944, w3945);
  FullAdder U146 (w3945, w3834, IN35[3], w3946, w3947);
  FullAdder U147 (w3947, w3836, IN36[3], w3948, w3949);
  FullAdder U148 (w3949, w3838, IN37[3], w3950, w3951);
  FullAdder U149 (w3951, w3840, IN38[3], w3952, w3953);
  FullAdder U150 (w3953, w3842, IN39[3], w3954, w3955);
  FullAdder U151 (w3955, w3844, IN40[3], w3956, w3957);
  FullAdder U152 (w3957, w3846, IN41[3], w3958, w3959);
  FullAdder U153 (w3959, w3848, IN42[3], w3960, w3961);
  FullAdder U154 (w3961, w3850, IN43[3], w3962, w3963);
  FullAdder U155 (w3963, w3852, IN44[3], w3964, w3965);
  FullAdder U156 (w3965, w3854, IN45[3], w3966, w3967);
  FullAdder U157 (w3967, w3856, IN46[3], w3968, w3969);
  FullAdder U158 (w3969, w3858, IN47[3], w3970, w3971);
  FullAdder U159 (w3971, w3860, IN48[3], w3972, w3973);
  FullAdder U160 (w3973, w3862, IN49[3], w3974, w3975);
  FullAdder U161 (w3975, w3864, IN50[3], w3976, w3977);
  FullAdder U162 (w3977, w3866, IN51[3], w3978, w3979);
  FullAdder U163 (w3979, w3868, IN52[3], w3980, w3981);
  FullAdder U164 (w3981, w3870, IN53[3], w3982, w3983);
  FullAdder U165 (w3983, w3872, IN54[3], w3984, w3985);
  FullAdder U166 (w3985, w3874, IN55[3], w3986, w3987);
  FullAdder U167 (w3987, w3876, IN56[3], w3988, w3989);
  FullAdder U168 (w3989, w3878, IN57[3], w3990, w3991);
  FullAdder U169 (w3991, w3880, IN58[1], w3992, w3993);
  FullAdder U170 (w3993, w3881, IN59[0], w3994, w3995);
  HalfAdder U171 (w3884, IN4[4], Out1[4], w3997);
  FullAdder U172 (w3997, w3886, IN5[4], w3998, w3999);
  FullAdder U173 (w3999, w3888, IN6[4], w4000, w4001);
  FullAdder U174 (w4001, w3890, IN7[4], w4002, w4003);
  FullAdder U175 (w4003, w3892, IN8[4], w4004, w4005);
  FullAdder U176 (w4005, w3894, IN9[4], w4006, w4007);
  FullAdder U177 (w4007, w3896, IN10[4], w4008, w4009);
  FullAdder U178 (w4009, w3898, IN11[4], w4010, w4011);
  FullAdder U179 (w4011, w3900, IN12[4], w4012, w4013);
  FullAdder U180 (w4013, w3902, IN13[4], w4014, w4015);
  FullAdder U181 (w4015, w3904, IN14[4], w4016, w4017);
  FullAdder U182 (w4017, w3906, IN15[4], w4018, w4019);
  FullAdder U183 (w4019, w3908, IN16[4], w4020, w4021);
  FullAdder U184 (w4021, w3910, IN17[4], w4022, w4023);
  FullAdder U185 (w4023, w3912, IN18[4], w4024, w4025);
  FullAdder U186 (w4025, w3914, IN19[4], w4026, w4027);
  FullAdder U187 (w4027, w3916, IN20[4], w4028, w4029);
  FullAdder U188 (w4029, w3918, IN21[4], w4030, w4031);
  FullAdder U189 (w4031, w3920, IN22[4], w4032, w4033);
  FullAdder U190 (w4033, w3922, IN23[4], w4034, w4035);
  FullAdder U191 (w4035, w3924, IN24[4], w4036, w4037);
  FullAdder U192 (w4037, w3926, IN25[4], w4038, w4039);
  FullAdder U193 (w4039, w3928, IN26[4], w4040, w4041);
  FullAdder U194 (w4041, w3930, IN27[4], w4042, w4043);
  FullAdder U195 (w4043, w3932, IN28[4], w4044, w4045);
  FullAdder U196 (w4045, w3934, IN29[4], w4046, w4047);
  FullAdder U197 (w4047, w3936, IN30[4], w4048, w4049);
  FullAdder U198 (w4049, w3938, IN31[4], w4050, w4051);
  FullAdder U199 (w4051, w3940, IN32[4], w4052, w4053);
  FullAdder U200 (w4053, w3942, IN33[4], w4054, w4055);
  FullAdder U201 (w4055, w3944, IN34[4], w4056, w4057);
  FullAdder U202 (w4057, w3946, IN35[4], w4058, w4059);
  FullAdder U203 (w4059, w3948, IN36[4], w4060, w4061);
  FullAdder U204 (w4061, w3950, IN37[4], w4062, w4063);
  FullAdder U205 (w4063, w3952, IN38[4], w4064, w4065);
  FullAdder U206 (w4065, w3954, IN39[4], w4066, w4067);
  FullAdder U207 (w4067, w3956, IN40[4], w4068, w4069);
  FullAdder U208 (w4069, w3958, IN41[4], w4070, w4071);
  FullAdder U209 (w4071, w3960, IN42[4], w4072, w4073);
  FullAdder U210 (w4073, w3962, IN43[4], w4074, w4075);
  FullAdder U211 (w4075, w3964, IN44[4], w4076, w4077);
  FullAdder U212 (w4077, w3966, IN45[4], w4078, w4079);
  FullAdder U213 (w4079, w3968, IN46[4], w4080, w4081);
  FullAdder U214 (w4081, w3970, IN47[4], w4082, w4083);
  FullAdder U215 (w4083, w3972, IN48[4], w4084, w4085);
  FullAdder U216 (w4085, w3974, IN49[4], w4086, w4087);
  FullAdder U217 (w4087, w3976, IN50[4], w4088, w4089);
  FullAdder U218 (w4089, w3978, IN51[4], w4090, w4091);
  FullAdder U219 (w4091, w3980, IN52[4], w4092, w4093);
  FullAdder U220 (w4093, w3982, IN53[4], w4094, w4095);
  FullAdder U221 (w4095, w3984, IN54[4], w4096, w4097);
  FullAdder U222 (w4097, w3986, IN55[4], w4098, w4099);
  FullAdder U223 (w4099, w3988, IN56[4], w4100, w4101);
  FullAdder U224 (w4101, w3990, IN57[4], w4102, w4103);
  FullAdder U225 (w4103, w3992, IN58[2], w4104, w4105);
  FullAdder U226 (w4105, w3994, IN59[1], w4106, w4107);
  FullAdder U227 (w4107, w3995, IN60[0], w4108, w4109);
  HalfAdder U228 (w3998, IN5[5], Out1[5], w4111);
  FullAdder U229 (w4111, w4000, IN6[5], w4112, w4113);
  FullAdder U230 (w4113, w4002, IN7[5], w4114, w4115);
  FullAdder U231 (w4115, w4004, IN8[5], w4116, w4117);
  FullAdder U232 (w4117, w4006, IN9[5], w4118, w4119);
  FullAdder U233 (w4119, w4008, IN10[5], w4120, w4121);
  FullAdder U234 (w4121, w4010, IN11[5], w4122, w4123);
  FullAdder U235 (w4123, w4012, IN12[5], w4124, w4125);
  FullAdder U236 (w4125, w4014, IN13[5], w4126, w4127);
  FullAdder U237 (w4127, w4016, IN14[5], w4128, w4129);
  FullAdder U238 (w4129, w4018, IN15[5], w4130, w4131);
  FullAdder U239 (w4131, w4020, IN16[5], w4132, w4133);
  FullAdder U240 (w4133, w4022, IN17[5], w4134, w4135);
  FullAdder U241 (w4135, w4024, IN18[5], w4136, w4137);
  FullAdder U242 (w4137, w4026, IN19[5], w4138, w4139);
  FullAdder U243 (w4139, w4028, IN20[5], w4140, w4141);
  FullAdder U244 (w4141, w4030, IN21[5], w4142, w4143);
  FullAdder U245 (w4143, w4032, IN22[5], w4144, w4145);
  FullAdder U246 (w4145, w4034, IN23[5], w4146, w4147);
  FullAdder U247 (w4147, w4036, IN24[5], w4148, w4149);
  FullAdder U248 (w4149, w4038, IN25[5], w4150, w4151);
  FullAdder U249 (w4151, w4040, IN26[5], w4152, w4153);
  FullAdder U250 (w4153, w4042, IN27[5], w4154, w4155);
  FullAdder U251 (w4155, w4044, IN28[5], w4156, w4157);
  FullAdder U252 (w4157, w4046, IN29[5], w4158, w4159);
  FullAdder U253 (w4159, w4048, IN30[5], w4160, w4161);
  FullAdder U254 (w4161, w4050, IN31[5], w4162, w4163);
  FullAdder U255 (w4163, w4052, IN32[5], w4164, w4165);
  FullAdder U256 (w4165, w4054, IN33[5], w4166, w4167);
  FullAdder U257 (w4167, w4056, IN34[5], w4168, w4169);
  FullAdder U258 (w4169, w4058, IN35[5], w4170, w4171);
  FullAdder U259 (w4171, w4060, IN36[5], w4172, w4173);
  FullAdder U260 (w4173, w4062, IN37[5], w4174, w4175);
  FullAdder U261 (w4175, w4064, IN38[5], w4176, w4177);
  FullAdder U262 (w4177, w4066, IN39[5], w4178, w4179);
  FullAdder U263 (w4179, w4068, IN40[5], w4180, w4181);
  FullAdder U264 (w4181, w4070, IN41[5], w4182, w4183);
  FullAdder U265 (w4183, w4072, IN42[5], w4184, w4185);
  FullAdder U266 (w4185, w4074, IN43[5], w4186, w4187);
  FullAdder U267 (w4187, w4076, IN44[5], w4188, w4189);
  FullAdder U268 (w4189, w4078, IN45[5], w4190, w4191);
  FullAdder U269 (w4191, w4080, IN46[5], w4192, w4193);
  FullAdder U270 (w4193, w4082, IN47[5], w4194, w4195);
  FullAdder U271 (w4195, w4084, IN48[5], w4196, w4197);
  FullAdder U272 (w4197, w4086, IN49[5], w4198, w4199);
  FullAdder U273 (w4199, w4088, IN50[5], w4200, w4201);
  FullAdder U274 (w4201, w4090, IN51[5], w4202, w4203);
  FullAdder U275 (w4203, w4092, IN52[5], w4204, w4205);
  FullAdder U276 (w4205, w4094, IN53[5], w4206, w4207);
  FullAdder U277 (w4207, w4096, IN54[5], w4208, w4209);
  FullAdder U278 (w4209, w4098, IN55[5], w4210, w4211);
  FullAdder U279 (w4211, w4100, IN56[5], w4212, w4213);
  FullAdder U280 (w4213, w4102, IN57[5], w4214, w4215);
  FullAdder U281 (w4215, w4104, IN58[3], w4216, w4217);
  FullAdder U282 (w4217, w4106, IN59[2], w4218, w4219);
  FullAdder U283 (w4219, w4108, IN60[1], w4220, w4221);
  FullAdder U284 (w4221, w4109, IN61[0], w4222, w4223);
  HalfAdder U285 (w4112, IN6[6], Out1[6], w4225);
  FullAdder U286 (w4225, w4114, IN7[6], w4226, w4227);
  FullAdder U287 (w4227, w4116, IN8[6], w4228, w4229);
  FullAdder U288 (w4229, w4118, IN9[6], w4230, w4231);
  FullAdder U289 (w4231, w4120, IN10[6], w4232, w4233);
  FullAdder U290 (w4233, w4122, IN11[6], w4234, w4235);
  FullAdder U291 (w4235, w4124, IN12[6], w4236, w4237);
  FullAdder U292 (w4237, w4126, IN13[6], w4238, w4239);
  FullAdder U293 (w4239, w4128, IN14[6], w4240, w4241);
  FullAdder U294 (w4241, w4130, IN15[6], w4242, w4243);
  FullAdder U295 (w4243, w4132, IN16[6], w4244, w4245);
  FullAdder U296 (w4245, w4134, IN17[6], w4246, w4247);
  FullAdder U297 (w4247, w4136, IN18[6], w4248, w4249);
  FullAdder U298 (w4249, w4138, IN19[6], w4250, w4251);
  FullAdder U299 (w4251, w4140, IN20[6], w4252, w4253);
  FullAdder U300 (w4253, w4142, IN21[6], w4254, w4255);
  FullAdder U301 (w4255, w4144, IN22[6], w4256, w4257);
  FullAdder U302 (w4257, w4146, IN23[6], w4258, w4259);
  FullAdder U303 (w4259, w4148, IN24[6], w4260, w4261);
  FullAdder U304 (w4261, w4150, IN25[6], w4262, w4263);
  FullAdder U305 (w4263, w4152, IN26[6], w4264, w4265);
  FullAdder U306 (w4265, w4154, IN27[6], w4266, w4267);
  FullAdder U307 (w4267, w4156, IN28[6], w4268, w4269);
  FullAdder U308 (w4269, w4158, IN29[6], w4270, w4271);
  FullAdder U309 (w4271, w4160, IN30[6], w4272, w4273);
  FullAdder U310 (w4273, w4162, IN31[6], w4274, w4275);
  FullAdder U311 (w4275, w4164, IN32[6], w4276, w4277);
  FullAdder U312 (w4277, w4166, IN33[6], w4278, w4279);
  FullAdder U313 (w4279, w4168, IN34[6], w4280, w4281);
  FullAdder U314 (w4281, w4170, IN35[6], w4282, w4283);
  FullAdder U315 (w4283, w4172, IN36[6], w4284, w4285);
  FullAdder U316 (w4285, w4174, IN37[6], w4286, w4287);
  FullAdder U317 (w4287, w4176, IN38[6], w4288, w4289);
  FullAdder U318 (w4289, w4178, IN39[6], w4290, w4291);
  FullAdder U319 (w4291, w4180, IN40[6], w4292, w4293);
  FullAdder U320 (w4293, w4182, IN41[6], w4294, w4295);
  FullAdder U321 (w4295, w4184, IN42[6], w4296, w4297);
  FullAdder U322 (w4297, w4186, IN43[6], w4298, w4299);
  FullAdder U323 (w4299, w4188, IN44[6], w4300, w4301);
  FullAdder U324 (w4301, w4190, IN45[6], w4302, w4303);
  FullAdder U325 (w4303, w4192, IN46[6], w4304, w4305);
  FullAdder U326 (w4305, w4194, IN47[6], w4306, w4307);
  FullAdder U327 (w4307, w4196, IN48[6], w4308, w4309);
  FullAdder U328 (w4309, w4198, IN49[6], w4310, w4311);
  FullAdder U329 (w4311, w4200, IN50[6], w4312, w4313);
  FullAdder U330 (w4313, w4202, IN51[6], w4314, w4315);
  FullAdder U331 (w4315, w4204, IN52[6], w4316, w4317);
  FullAdder U332 (w4317, w4206, IN53[6], w4318, w4319);
  FullAdder U333 (w4319, w4208, IN54[6], w4320, w4321);
  FullAdder U334 (w4321, w4210, IN55[6], w4322, w4323);
  FullAdder U335 (w4323, w4212, IN56[6], w4324, w4325);
  FullAdder U336 (w4325, w4214, IN57[6], w4326, w4327);
  FullAdder U337 (w4327, w4216, IN58[4], w4328, w4329);
  FullAdder U338 (w4329, w4218, IN59[3], w4330, w4331);
  FullAdder U339 (w4331, w4220, IN60[2], w4332, w4333);
  FullAdder U340 (w4333, w4222, IN61[1], w4334, w4335);
  FullAdder U341 (w4335, w4223, IN62[0], w4336, w4337);
  HalfAdder U342 (w4226, IN7[7], Out1[7], w4339);
  FullAdder U343 (w4339, w4228, IN8[7], w4340, w4341);
  FullAdder U344 (w4341, w4230, IN9[7], w4342, w4343);
  FullAdder U345 (w4343, w4232, IN10[7], w4344, w4345);
  FullAdder U346 (w4345, w4234, IN11[7], w4346, w4347);
  FullAdder U347 (w4347, w4236, IN12[7], w4348, w4349);
  FullAdder U348 (w4349, w4238, IN13[7], w4350, w4351);
  FullAdder U349 (w4351, w4240, IN14[7], w4352, w4353);
  FullAdder U350 (w4353, w4242, IN15[7], w4354, w4355);
  FullAdder U351 (w4355, w4244, IN16[7], w4356, w4357);
  FullAdder U352 (w4357, w4246, IN17[7], w4358, w4359);
  FullAdder U353 (w4359, w4248, IN18[7], w4360, w4361);
  FullAdder U354 (w4361, w4250, IN19[7], w4362, w4363);
  FullAdder U355 (w4363, w4252, IN20[7], w4364, w4365);
  FullAdder U356 (w4365, w4254, IN21[7], w4366, w4367);
  FullAdder U357 (w4367, w4256, IN22[7], w4368, w4369);
  FullAdder U358 (w4369, w4258, IN23[7], w4370, w4371);
  FullAdder U359 (w4371, w4260, IN24[7], w4372, w4373);
  FullAdder U360 (w4373, w4262, IN25[7], w4374, w4375);
  FullAdder U361 (w4375, w4264, IN26[7], w4376, w4377);
  FullAdder U362 (w4377, w4266, IN27[7], w4378, w4379);
  FullAdder U363 (w4379, w4268, IN28[7], w4380, w4381);
  FullAdder U364 (w4381, w4270, IN29[7], w4382, w4383);
  FullAdder U365 (w4383, w4272, IN30[7], w4384, w4385);
  FullAdder U366 (w4385, w4274, IN31[7], w4386, w4387);
  FullAdder U367 (w4387, w4276, IN32[7], w4388, w4389);
  FullAdder U368 (w4389, w4278, IN33[7], w4390, w4391);
  FullAdder U369 (w4391, w4280, IN34[7], w4392, w4393);
  FullAdder U370 (w4393, w4282, IN35[7], w4394, w4395);
  FullAdder U371 (w4395, w4284, IN36[7], w4396, w4397);
  FullAdder U372 (w4397, w4286, IN37[7], w4398, w4399);
  FullAdder U373 (w4399, w4288, IN38[7], w4400, w4401);
  FullAdder U374 (w4401, w4290, IN39[7], w4402, w4403);
  FullAdder U375 (w4403, w4292, IN40[7], w4404, w4405);
  FullAdder U376 (w4405, w4294, IN41[7], w4406, w4407);
  FullAdder U377 (w4407, w4296, IN42[7], w4408, w4409);
  FullAdder U378 (w4409, w4298, IN43[7], w4410, w4411);
  FullAdder U379 (w4411, w4300, IN44[7], w4412, w4413);
  FullAdder U380 (w4413, w4302, IN45[7], w4414, w4415);
  FullAdder U381 (w4415, w4304, IN46[7], w4416, w4417);
  FullAdder U382 (w4417, w4306, IN47[7], w4418, w4419);
  FullAdder U383 (w4419, w4308, IN48[7], w4420, w4421);
  FullAdder U384 (w4421, w4310, IN49[7], w4422, w4423);
  FullAdder U385 (w4423, w4312, IN50[7], w4424, w4425);
  FullAdder U386 (w4425, w4314, IN51[7], w4426, w4427);
  FullAdder U387 (w4427, w4316, IN52[7], w4428, w4429);
  FullAdder U388 (w4429, w4318, IN53[7], w4430, w4431);
  FullAdder U389 (w4431, w4320, IN54[7], w4432, w4433);
  FullAdder U390 (w4433, w4322, IN55[7], w4434, w4435);
  FullAdder U391 (w4435, w4324, IN56[7], w4436, w4437);
  FullAdder U392 (w4437, w4326, IN57[7], w4438, w4439);
  FullAdder U393 (w4439, w4328, IN58[5], w4440, w4441);
  FullAdder U394 (w4441, w4330, IN59[4], w4442, w4443);
  FullAdder U395 (w4443, w4332, IN60[3], w4444, w4445);
  FullAdder U396 (w4445, w4334, IN61[2], w4446, w4447);
  FullAdder U397 (w4447, w4336, IN62[1], w4448, w4449);
  FullAdder U398 (w4449, w4337, IN63[0], w4450, w4451);
  HalfAdder U399 (w4340, IN8[8], Out1[8], w4453);
  FullAdder U400 (w4453, w4342, IN9[8], w4454, w4455);
  FullAdder U401 (w4455, w4344, IN10[8], w4456, w4457);
  FullAdder U402 (w4457, w4346, IN11[8], w4458, w4459);
  FullAdder U403 (w4459, w4348, IN12[8], w4460, w4461);
  FullAdder U404 (w4461, w4350, IN13[8], w4462, w4463);
  FullAdder U405 (w4463, w4352, IN14[8], w4464, w4465);
  FullAdder U406 (w4465, w4354, IN15[8], w4466, w4467);
  FullAdder U407 (w4467, w4356, IN16[8], w4468, w4469);
  FullAdder U408 (w4469, w4358, IN17[8], w4470, w4471);
  FullAdder U409 (w4471, w4360, IN18[8], w4472, w4473);
  FullAdder U410 (w4473, w4362, IN19[8], w4474, w4475);
  FullAdder U411 (w4475, w4364, IN20[8], w4476, w4477);
  FullAdder U412 (w4477, w4366, IN21[8], w4478, w4479);
  FullAdder U413 (w4479, w4368, IN22[8], w4480, w4481);
  FullAdder U414 (w4481, w4370, IN23[8], w4482, w4483);
  FullAdder U415 (w4483, w4372, IN24[8], w4484, w4485);
  FullAdder U416 (w4485, w4374, IN25[8], w4486, w4487);
  FullAdder U417 (w4487, w4376, IN26[8], w4488, w4489);
  FullAdder U418 (w4489, w4378, IN27[8], w4490, w4491);
  FullAdder U419 (w4491, w4380, IN28[8], w4492, w4493);
  FullAdder U420 (w4493, w4382, IN29[8], w4494, w4495);
  FullAdder U421 (w4495, w4384, IN30[8], w4496, w4497);
  FullAdder U422 (w4497, w4386, IN31[8], w4498, w4499);
  FullAdder U423 (w4499, w4388, IN32[8], w4500, w4501);
  FullAdder U424 (w4501, w4390, IN33[8], w4502, w4503);
  FullAdder U425 (w4503, w4392, IN34[8], w4504, w4505);
  FullAdder U426 (w4505, w4394, IN35[8], w4506, w4507);
  FullAdder U427 (w4507, w4396, IN36[8], w4508, w4509);
  FullAdder U428 (w4509, w4398, IN37[8], w4510, w4511);
  FullAdder U429 (w4511, w4400, IN38[8], w4512, w4513);
  FullAdder U430 (w4513, w4402, IN39[8], w4514, w4515);
  FullAdder U431 (w4515, w4404, IN40[8], w4516, w4517);
  FullAdder U432 (w4517, w4406, IN41[8], w4518, w4519);
  FullAdder U433 (w4519, w4408, IN42[8], w4520, w4521);
  FullAdder U434 (w4521, w4410, IN43[8], w4522, w4523);
  FullAdder U435 (w4523, w4412, IN44[8], w4524, w4525);
  FullAdder U436 (w4525, w4414, IN45[8], w4526, w4527);
  FullAdder U437 (w4527, w4416, IN46[8], w4528, w4529);
  FullAdder U438 (w4529, w4418, IN47[8], w4530, w4531);
  FullAdder U439 (w4531, w4420, IN48[8], w4532, w4533);
  FullAdder U440 (w4533, w4422, IN49[8], w4534, w4535);
  FullAdder U441 (w4535, w4424, IN50[8], w4536, w4537);
  FullAdder U442 (w4537, w4426, IN51[8], w4538, w4539);
  FullAdder U443 (w4539, w4428, IN52[8], w4540, w4541);
  FullAdder U444 (w4541, w4430, IN53[8], w4542, w4543);
  FullAdder U445 (w4543, w4432, IN54[8], w4544, w4545);
  FullAdder U446 (w4545, w4434, IN55[8], w4546, w4547);
  FullAdder U447 (w4547, w4436, IN56[8], w4548, w4549);
  FullAdder U448 (w4549, w4438, IN57[8], w4550, w4551);
  FullAdder U449 (w4551, w4440, IN58[6], w4552, w4553);
  FullAdder U450 (w4553, w4442, IN59[5], w4554, w4555);
  FullAdder U451 (w4555, w4444, IN60[4], w4556, w4557);
  FullAdder U452 (w4557, w4446, IN61[3], w4558, w4559);
  FullAdder U453 (w4559, w4448, IN62[2], w4560, w4561);
  FullAdder U454 (w4561, w4450, IN63[1], w4562, w4563);
  FullAdder U455 (w4563, w4451, IN64[0], w4564, w4565);
  HalfAdder U456 (w4454, IN9[9], Out1[9], w4567);
  FullAdder U457 (w4567, w4456, IN10[9], w4568, w4569);
  FullAdder U458 (w4569, w4458, IN11[9], w4570, w4571);
  FullAdder U459 (w4571, w4460, IN12[9], w4572, w4573);
  FullAdder U460 (w4573, w4462, IN13[9], w4574, w4575);
  FullAdder U461 (w4575, w4464, IN14[9], w4576, w4577);
  FullAdder U462 (w4577, w4466, IN15[9], w4578, w4579);
  FullAdder U463 (w4579, w4468, IN16[9], w4580, w4581);
  FullAdder U464 (w4581, w4470, IN17[9], w4582, w4583);
  FullAdder U465 (w4583, w4472, IN18[9], w4584, w4585);
  FullAdder U466 (w4585, w4474, IN19[9], w4586, w4587);
  FullAdder U467 (w4587, w4476, IN20[9], w4588, w4589);
  FullAdder U468 (w4589, w4478, IN21[9], w4590, w4591);
  FullAdder U469 (w4591, w4480, IN22[9], w4592, w4593);
  FullAdder U470 (w4593, w4482, IN23[9], w4594, w4595);
  FullAdder U471 (w4595, w4484, IN24[9], w4596, w4597);
  FullAdder U472 (w4597, w4486, IN25[9], w4598, w4599);
  FullAdder U473 (w4599, w4488, IN26[9], w4600, w4601);
  FullAdder U474 (w4601, w4490, IN27[9], w4602, w4603);
  FullAdder U475 (w4603, w4492, IN28[9], w4604, w4605);
  FullAdder U476 (w4605, w4494, IN29[9], w4606, w4607);
  FullAdder U477 (w4607, w4496, IN30[9], w4608, w4609);
  FullAdder U478 (w4609, w4498, IN31[9], w4610, w4611);
  FullAdder U479 (w4611, w4500, IN32[9], w4612, w4613);
  FullAdder U480 (w4613, w4502, IN33[9], w4614, w4615);
  FullAdder U481 (w4615, w4504, IN34[9], w4616, w4617);
  FullAdder U482 (w4617, w4506, IN35[9], w4618, w4619);
  FullAdder U483 (w4619, w4508, IN36[9], w4620, w4621);
  FullAdder U484 (w4621, w4510, IN37[9], w4622, w4623);
  FullAdder U485 (w4623, w4512, IN38[9], w4624, w4625);
  FullAdder U486 (w4625, w4514, IN39[9], w4626, w4627);
  FullAdder U487 (w4627, w4516, IN40[9], w4628, w4629);
  FullAdder U488 (w4629, w4518, IN41[9], w4630, w4631);
  FullAdder U489 (w4631, w4520, IN42[9], w4632, w4633);
  FullAdder U490 (w4633, w4522, IN43[9], w4634, w4635);
  FullAdder U491 (w4635, w4524, IN44[9], w4636, w4637);
  FullAdder U492 (w4637, w4526, IN45[9], w4638, w4639);
  FullAdder U493 (w4639, w4528, IN46[9], w4640, w4641);
  FullAdder U494 (w4641, w4530, IN47[9], w4642, w4643);
  FullAdder U495 (w4643, w4532, IN48[9], w4644, w4645);
  FullAdder U496 (w4645, w4534, IN49[9], w4646, w4647);
  FullAdder U497 (w4647, w4536, IN50[9], w4648, w4649);
  FullAdder U498 (w4649, w4538, IN51[9], w4650, w4651);
  FullAdder U499 (w4651, w4540, IN52[9], w4652, w4653);
  FullAdder U500 (w4653, w4542, IN53[9], w4654, w4655);
  FullAdder U501 (w4655, w4544, IN54[9], w4656, w4657);
  FullAdder U502 (w4657, w4546, IN55[9], w4658, w4659);
  FullAdder U503 (w4659, w4548, IN56[9], w4660, w4661);
  FullAdder U504 (w4661, w4550, IN57[9], w4662, w4663);
  FullAdder U505 (w4663, w4552, IN58[7], w4664, w4665);
  FullAdder U506 (w4665, w4554, IN59[6], w4666, w4667);
  FullAdder U507 (w4667, w4556, IN60[5], w4668, w4669);
  FullAdder U508 (w4669, w4558, IN61[4], w4670, w4671);
  FullAdder U509 (w4671, w4560, IN62[3], w4672, w4673);
  FullAdder U510 (w4673, w4562, IN63[2], w4674, w4675);
  FullAdder U511 (w4675, w4564, IN64[1], w4676, w4677);
  FullAdder U512 (w4677, w4565, IN65[0], w4678, w4679);
  HalfAdder U513 (w4568, IN10[10], Out1[10], w4681);
  FullAdder U514 (w4681, w4570, IN11[10], w4682, w4683);
  FullAdder U515 (w4683, w4572, IN12[10], w4684, w4685);
  FullAdder U516 (w4685, w4574, IN13[10], w4686, w4687);
  FullAdder U517 (w4687, w4576, IN14[10], w4688, w4689);
  FullAdder U518 (w4689, w4578, IN15[10], w4690, w4691);
  FullAdder U519 (w4691, w4580, IN16[10], w4692, w4693);
  FullAdder U520 (w4693, w4582, IN17[10], w4694, w4695);
  FullAdder U521 (w4695, w4584, IN18[10], w4696, w4697);
  FullAdder U522 (w4697, w4586, IN19[10], w4698, w4699);
  FullAdder U523 (w4699, w4588, IN20[10], w4700, w4701);
  FullAdder U524 (w4701, w4590, IN21[10], w4702, w4703);
  FullAdder U525 (w4703, w4592, IN22[10], w4704, w4705);
  FullAdder U526 (w4705, w4594, IN23[10], w4706, w4707);
  FullAdder U527 (w4707, w4596, IN24[10], w4708, w4709);
  FullAdder U528 (w4709, w4598, IN25[10], w4710, w4711);
  FullAdder U529 (w4711, w4600, IN26[10], w4712, w4713);
  FullAdder U530 (w4713, w4602, IN27[10], w4714, w4715);
  FullAdder U531 (w4715, w4604, IN28[10], w4716, w4717);
  FullAdder U532 (w4717, w4606, IN29[10], w4718, w4719);
  FullAdder U533 (w4719, w4608, IN30[10], w4720, w4721);
  FullAdder U534 (w4721, w4610, IN31[10], w4722, w4723);
  FullAdder U535 (w4723, w4612, IN32[10], w4724, w4725);
  FullAdder U536 (w4725, w4614, IN33[10], w4726, w4727);
  FullAdder U537 (w4727, w4616, IN34[10], w4728, w4729);
  FullAdder U538 (w4729, w4618, IN35[10], w4730, w4731);
  FullAdder U539 (w4731, w4620, IN36[10], w4732, w4733);
  FullAdder U540 (w4733, w4622, IN37[10], w4734, w4735);
  FullAdder U541 (w4735, w4624, IN38[10], w4736, w4737);
  FullAdder U542 (w4737, w4626, IN39[10], w4738, w4739);
  FullAdder U543 (w4739, w4628, IN40[10], w4740, w4741);
  FullAdder U544 (w4741, w4630, IN41[10], w4742, w4743);
  FullAdder U545 (w4743, w4632, IN42[10], w4744, w4745);
  FullAdder U546 (w4745, w4634, IN43[10], w4746, w4747);
  FullAdder U547 (w4747, w4636, IN44[10], w4748, w4749);
  FullAdder U548 (w4749, w4638, IN45[10], w4750, w4751);
  FullAdder U549 (w4751, w4640, IN46[10], w4752, w4753);
  FullAdder U550 (w4753, w4642, IN47[10], w4754, w4755);
  FullAdder U551 (w4755, w4644, IN48[10], w4756, w4757);
  FullAdder U552 (w4757, w4646, IN49[10], w4758, w4759);
  FullAdder U553 (w4759, w4648, IN50[10], w4760, w4761);
  FullAdder U554 (w4761, w4650, IN51[10], w4762, w4763);
  FullAdder U555 (w4763, w4652, IN52[10], w4764, w4765);
  FullAdder U556 (w4765, w4654, IN53[10], w4766, w4767);
  FullAdder U557 (w4767, w4656, IN54[10], w4768, w4769);
  FullAdder U558 (w4769, w4658, IN55[10], w4770, w4771);
  FullAdder U559 (w4771, w4660, IN56[10], w4772, w4773);
  FullAdder U560 (w4773, w4662, IN57[10], w4774, w4775);
  FullAdder U561 (w4775, w4664, IN58[8], w4776, w4777);
  FullAdder U562 (w4777, w4666, IN59[7], w4778, w4779);
  FullAdder U563 (w4779, w4668, IN60[6], w4780, w4781);
  FullAdder U564 (w4781, w4670, IN61[5], w4782, w4783);
  FullAdder U565 (w4783, w4672, IN62[4], w4784, w4785);
  FullAdder U566 (w4785, w4674, IN63[3], w4786, w4787);
  FullAdder U567 (w4787, w4676, IN64[2], w4788, w4789);
  FullAdder U568 (w4789, w4678, IN65[1], w4790, w4791);
  FullAdder U569 (w4791, w4679, IN66[0], w4792, w4793);
  HalfAdder U570 (w4682, IN11[11], Out1[11], w4795);
  FullAdder U571 (w4795, w4684, IN12[11], w4796, w4797);
  FullAdder U572 (w4797, w4686, IN13[11], w4798, w4799);
  FullAdder U573 (w4799, w4688, IN14[11], w4800, w4801);
  FullAdder U574 (w4801, w4690, IN15[11], w4802, w4803);
  FullAdder U575 (w4803, w4692, IN16[11], w4804, w4805);
  FullAdder U576 (w4805, w4694, IN17[11], w4806, w4807);
  FullAdder U577 (w4807, w4696, IN18[11], w4808, w4809);
  FullAdder U578 (w4809, w4698, IN19[11], w4810, w4811);
  FullAdder U579 (w4811, w4700, IN20[11], w4812, w4813);
  FullAdder U580 (w4813, w4702, IN21[11], w4814, w4815);
  FullAdder U581 (w4815, w4704, IN22[11], w4816, w4817);
  FullAdder U582 (w4817, w4706, IN23[11], w4818, w4819);
  FullAdder U583 (w4819, w4708, IN24[11], w4820, w4821);
  FullAdder U584 (w4821, w4710, IN25[11], w4822, w4823);
  FullAdder U585 (w4823, w4712, IN26[11], w4824, w4825);
  FullAdder U586 (w4825, w4714, IN27[11], w4826, w4827);
  FullAdder U587 (w4827, w4716, IN28[11], w4828, w4829);
  FullAdder U588 (w4829, w4718, IN29[11], w4830, w4831);
  FullAdder U589 (w4831, w4720, IN30[11], w4832, w4833);
  FullAdder U590 (w4833, w4722, IN31[11], w4834, w4835);
  FullAdder U591 (w4835, w4724, IN32[11], w4836, w4837);
  FullAdder U592 (w4837, w4726, IN33[11], w4838, w4839);
  FullAdder U593 (w4839, w4728, IN34[11], w4840, w4841);
  FullAdder U594 (w4841, w4730, IN35[11], w4842, w4843);
  FullAdder U595 (w4843, w4732, IN36[11], w4844, w4845);
  FullAdder U596 (w4845, w4734, IN37[11], w4846, w4847);
  FullAdder U597 (w4847, w4736, IN38[11], w4848, w4849);
  FullAdder U598 (w4849, w4738, IN39[11], w4850, w4851);
  FullAdder U599 (w4851, w4740, IN40[11], w4852, w4853);
  FullAdder U600 (w4853, w4742, IN41[11], w4854, w4855);
  FullAdder U601 (w4855, w4744, IN42[11], w4856, w4857);
  FullAdder U602 (w4857, w4746, IN43[11], w4858, w4859);
  FullAdder U603 (w4859, w4748, IN44[11], w4860, w4861);
  FullAdder U604 (w4861, w4750, IN45[11], w4862, w4863);
  FullAdder U605 (w4863, w4752, IN46[11], w4864, w4865);
  FullAdder U606 (w4865, w4754, IN47[11], w4866, w4867);
  FullAdder U607 (w4867, w4756, IN48[11], w4868, w4869);
  FullAdder U608 (w4869, w4758, IN49[11], w4870, w4871);
  FullAdder U609 (w4871, w4760, IN50[11], w4872, w4873);
  FullAdder U610 (w4873, w4762, IN51[11], w4874, w4875);
  FullAdder U611 (w4875, w4764, IN52[11], w4876, w4877);
  FullAdder U612 (w4877, w4766, IN53[11], w4878, w4879);
  FullAdder U613 (w4879, w4768, IN54[11], w4880, w4881);
  FullAdder U614 (w4881, w4770, IN55[11], w4882, w4883);
  FullAdder U615 (w4883, w4772, IN56[11], w4884, w4885);
  FullAdder U616 (w4885, w4774, IN57[11], w4886, w4887);
  FullAdder U617 (w4887, w4776, IN58[9], w4888, w4889);
  FullAdder U618 (w4889, w4778, IN59[8], w4890, w4891);
  FullAdder U619 (w4891, w4780, IN60[7], w4892, w4893);
  FullAdder U620 (w4893, w4782, IN61[6], w4894, w4895);
  FullAdder U621 (w4895, w4784, IN62[5], w4896, w4897);
  FullAdder U622 (w4897, w4786, IN63[4], w4898, w4899);
  FullAdder U623 (w4899, w4788, IN64[3], w4900, w4901);
  FullAdder U624 (w4901, w4790, IN65[2], w4902, w4903);
  FullAdder U625 (w4903, w4792, IN66[1], w4904, w4905);
  FullAdder U626 (w4905, w4793, IN67[0], w4906, w4907);
  HalfAdder U627 (w4796, IN12[12], Out1[12], w4909);
  FullAdder U628 (w4909, w4798, IN13[12], w4910, w4911);
  FullAdder U629 (w4911, w4800, IN14[12], w4912, w4913);
  FullAdder U630 (w4913, w4802, IN15[12], w4914, w4915);
  FullAdder U631 (w4915, w4804, IN16[12], w4916, w4917);
  FullAdder U632 (w4917, w4806, IN17[12], w4918, w4919);
  FullAdder U633 (w4919, w4808, IN18[12], w4920, w4921);
  FullAdder U634 (w4921, w4810, IN19[12], w4922, w4923);
  FullAdder U635 (w4923, w4812, IN20[12], w4924, w4925);
  FullAdder U636 (w4925, w4814, IN21[12], w4926, w4927);
  FullAdder U637 (w4927, w4816, IN22[12], w4928, w4929);
  FullAdder U638 (w4929, w4818, IN23[12], w4930, w4931);
  FullAdder U639 (w4931, w4820, IN24[12], w4932, w4933);
  FullAdder U640 (w4933, w4822, IN25[12], w4934, w4935);
  FullAdder U641 (w4935, w4824, IN26[12], w4936, w4937);
  FullAdder U642 (w4937, w4826, IN27[12], w4938, w4939);
  FullAdder U643 (w4939, w4828, IN28[12], w4940, w4941);
  FullAdder U644 (w4941, w4830, IN29[12], w4942, w4943);
  FullAdder U645 (w4943, w4832, IN30[12], w4944, w4945);
  FullAdder U646 (w4945, w4834, IN31[12], w4946, w4947);
  FullAdder U647 (w4947, w4836, IN32[12], w4948, w4949);
  FullAdder U648 (w4949, w4838, IN33[12], w4950, w4951);
  FullAdder U649 (w4951, w4840, IN34[12], w4952, w4953);
  FullAdder U650 (w4953, w4842, IN35[12], w4954, w4955);
  FullAdder U651 (w4955, w4844, IN36[12], w4956, w4957);
  FullAdder U652 (w4957, w4846, IN37[12], w4958, w4959);
  FullAdder U653 (w4959, w4848, IN38[12], w4960, w4961);
  FullAdder U654 (w4961, w4850, IN39[12], w4962, w4963);
  FullAdder U655 (w4963, w4852, IN40[12], w4964, w4965);
  FullAdder U656 (w4965, w4854, IN41[12], w4966, w4967);
  FullAdder U657 (w4967, w4856, IN42[12], w4968, w4969);
  FullAdder U658 (w4969, w4858, IN43[12], w4970, w4971);
  FullAdder U659 (w4971, w4860, IN44[12], w4972, w4973);
  FullAdder U660 (w4973, w4862, IN45[12], w4974, w4975);
  FullAdder U661 (w4975, w4864, IN46[12], w4976, w4977);
  FullAdder U662 (w4977, w4866, IN47[12], w4978, w4979);
  FullAdder U663 (w4979, w4868, IN48[12], w4980, w4981);
  FullAdder U664 (w4981, w4870, IN49[12], w4982, w4983);
  FullAdder U665 (w4983, w4872, IN50[12], w4984, w4985);
  FullAdder U666 (w4985, w4874, IN51[12], w4986, w4987);
  FullAdder U667 (w4987, w4876, IN52[12], w4988, w4989);
  FullAdder U668 (w4989, w4878, IN53[12], w4990, w4991);
  FullAdder U669 (w4991, w4880, IN54[12], w4992, w4993);
  FullAdder U670 (w4993, w4882, IN55[12], w4994, w4995);
  FullAdder U671 (w4995, w4884, IN56[12], w4996, w4997);
  FullAdder U672 (w4997, w4886, IN57[12], w4998, w4999);
  FullAdder U673 (w4999, w4888, IN58[10], w5000, w5001);
  FullAdder U674 (w5001, w4890, IN59[9], w5002, w5003);
  FullAdder U675 (w5003, w4892, IN60[8], w5004, w5005);
  FullAdder U676 (w5005, w4894, IN61[7], w5006, w5007);
  FullAdder U677 (w5007, w4896, IN62[6], w5008, w5009);
  FullAdder U678 (w5009, w4898, IN63[5], w5010, w5011);
  FullAdder U679 (w5011, w4900, IN64[4], w5012, w5013);
  FullAdder U680 (w5013, w4902, IN65[3], w5014, w5015);
  FullAdder U681 (w5015, w4904, IN66[2], w5016, w5017);
  FullAdder U682 (w5017, w4906, IN67[1], w5018, w5019);
  FullAdder U683 (w5019, w4907, IN68[0], w5020, w5021);
  HalfAdder U684 (w4910, IN13[13], Out1[13], w5023);
  FullAdder U685 (w5023, w4912, IN14[13], w5024, w5025);
  FullAdder U686 (w5025, w4914, IN15[13], w5026, w5027);
  FullAdder U687 (w5027, w4916, IN16[13], w5028, w5029);
  FullAdder U688 (w5029, w4918, IN17[13], w5030, w5031);
  FullAdder U689 (w5031, w4920, IN18[13], w5032, w5033);
  FullAdder U690 (w5033, w4922, IN19[13], w5034, w5035);
  FullAdder U691 (w5035, w4924, IN20[13], w5036, w5037);
  FullAdder U692 (w5037, w4926, IN21[13], w5038, w5039);
  FullAdder U693 (w5039, w4928, IN22[13], w5040, w5041);
  FullAdder U694 (w5041, w4930, IN23[13], w5042, w5043);
  FullAdder U695 (w5043, w4932, IN24[13], w5044, w5045);
  FullAdder U696 (w5045, w4934, IN25[13], w5046, w5047);
  FullAdder U697 (w5047, w4936, IN26[13], w5048, w5049);
  FullAdder U698 (w5049, w4938, IN27[13], w5050, w5051);
  FullAdder U699 (w5051, w4940, IN28[13], w5052, w5053);
  FullAdder U700 (w5053, w4942, IN29[13], w5054, w5055);
  FullAdder U701 (w5055, w4944, IN30[13], w5056, w5057);
  FullAdder U702 (w5057, w4946, IN31[13], w5058, w5059);
  FullAdder U703 (w5059, w4948, IN32[13], w5060, w5061);
  FullAdder U704 (w5061, w4950, IN33[13], w5062, w5063);
  FullAdder U705 (w5063, w4952, IN34[13], w5064, w5065);
  FullAdder U706 (w5065, w4954, IN35[13], w5066, w5067);
  FullAdder U707 (w5067, w4956, IN36[13], w5068, w5069);
  FullAdder U708 (w5069, w4958, IN37[13], w5070, w5071);
  FullAdder U709 (w5071, w4960, IN38[13], w5072, w5073);
  FullAdder U710 (w5073, w4962, IN39[13], w5074, w5075);
  FullAdder U711 (w5075, w4964, IN40[13], w5076, w5077);
  FullAdder U712 (w5077, w4966, IN41[13], w5078, w5079);
  FullAdder U713 (w5079, w4968, IN42[13], w5080, w5081);
  FullAdder U714 (w5081, w4970, IN43[13], w5082, w5083);
  FullAdder U715 (w5083, w4972, IN44[13], w5084, w5085);
  FullAdder U716 (w5085, w4974, IN45[13], w5086, w5087);
  FullAdder U717 (w5087, w4976, IN46[13], w5088, w5089);
  FullAdder U718 (w5089, w4978, IN47[13], w5090, w5091);
  FullAdder U719 (w5091, w4980, IN48[13], w5092, w5093);
  FullAdder U720 (w5093, w4982, IN49[13], w5094, w5095);
  FullAdder U721 (w5095, w4984, IN50[13], w5096, w5097);
  FullAdder U722 (w5097, w4986, IN51[13], w5098, w5099);
  FullAdder U723 (w5099, w4988, IN52[13], w5100, w5101);
  FullAdder U724 (w5101, w4990, IN53[13], w5102, w5103);
  FullAdder U725 (w5103, w4992, IN54[13], w5104, w5105);
  FullAdder U726 (w5105, w4994, IN55[13], w5106, w5107);
  FullAdder U727 (w5107, w4996, IN56[13], w5108, w5109);
  FullAdder U728 (w5109, w4998, IN57[13], w5110, w5111);
  FullAdder U729 (w5111, w5000, IN58[11], w5112, w5113);
  FullAdder U730 (w5113, w5002, IN59[10], w5114, w5115);
  FullAdder U731 (w5115, w5004, IN60[9], w5116, w5117);
  FullAdder U732 (w5117, w5006, IN61[8], w5118, w5119);
  FullAdder U733 (w5119, w5008, IN62[7], w5120, w5121);
  FullAdder U734 (w5121, w5010, IN63[6], w5122, w5123);
  FullAdder U735 (w5123, w5012, IN64[5], w5124, w5125);
  FullAdder U736 (w5125, w5014, IN65[4], w5126, w5127);
  FullAdder U737 (w5127, w5016, IN66[3], w5128, w5129);
  FullAdder U738 (w5129, w5018, IN67[2], w5130, w5131);
  FullAdder U739 (w5131, w5020, IN68[1], w5132, w5133);
  FullAdder U740 (w5133, w5021, IN69[0], w5134, w5135);
  HalfAdder U741 (w5024, IN14[14], Out1[14], w5137);
  FullAdder U742 (w5137, w5026, IN15[14], w5138, w5139);
  FullAdder U743 (w5139, w5028, IN16[14], w5140, w5141);
  FullAdder U744 (w5141, w5030, IN17[14], w5142, w5143);
  FullAdder U745 (w5143, w5032, IN18[14], w5144, w5145);
  FullAdder U746 (w5145, w5034, IN19[14], w5146, w5147);
  FullAdder U747 (w5147, w5036, IN20[14], w5148, w5149);
  FullAdder U748 (w5149, w5038, IN21[14], w5150, w5151);
  FullAdder U749 (w5151, w5040, IN22[14], w5152, w5153);
  FullAdder U750 (w5153, w5042, IN23[14], w5154, w5155);
  FullAdder U751 (w5155, w5044, IN24[14], w5156, w5157);
  FullAdder U752 (w5157, w5046, IN25[14], w5158, w5159);
  FullAdder U753 (w5159, w5048, IN26[14], w5160, w5161);
  FullAdder U754 (w5161, w5050, IN27[14], w5162, w5163);
  FullAdder U755 (w5163, w5052, IN28[14], w5164, w5165);
  FullAdder U756 (w5165, w5054, IN29[14], w5166, w5167);
  FullAdder U757 (w5167, w5056, IN30[14], w5168, w5169);
  FullAdder U758 (w5169, w5058, IN31[14], w5170, w5171);
  FullAdder U759 (w5171, w5060, IN32[14], w5172, w5173);
  FullAdder U760 (w5173, w5062, IN33[14], w5174, w5175);
  FullAdder U761 (w5175, w5064, IN34[14], w5176, w5177);
  FullAdder U762 (w5177, w5066, IN35[14], w5178, w5179);
  FullAdder U763 (w5179, w5068, IN36[14], w5180, w5181);
  FullAdder U764 (w5181, w5070, IN37[14], w5182, w5183);
  FullAdder U765 (w5183, w5072, IN38[14], w5184, w5185);
  FullAdder U766 (w5185, w5074, IN39[14], w5186, w5187);
  FullAdder U767 (w5187, w5076, IN40[14], w5188, w5189);
  FullAdder U768 (w5189, w5078, IN41[14], w5190, w5191);
  FullAdder U769 (w5191, w5080, IN42[14], w5192, w5193);
  FullAdder U770 (w5193, w5082, IN43[14], w5194, w5195);
  FullAdder U771 (w5195, w5084, IN44[14], w5196, w5197);
  FullAdder U772 (w5197, w5086, IN45[14], w5198, w5199);
  FullAdder U773 (w5199, w5088, IN46[14], w5200, w5201);
  FullAdder U774 (w5201, w5090, IN47[14], w5202, w5203);
  FullAdder U775 (w5203, w5092, IN48[14], w5204, w5205);
  FullAdder U776 (w5205, w5094, IN49[14], w5206, w5207);
  FullAdder U777 (w5207, w5096, IN50[14], w5208, w5209);
  FullAdder U778 (w5209, w5098, IN51[14], w5210, w5211);
  FullAdder U779 (w5211, w5100, IN52[14], w5212, w5213);
  FullAdder U780 (w5213, w5102, IN53[14], w5214, w5215);
  FullAdder U781 (w5215, w5104, IN54[14], w5216, w5217);
  FullAdder U782 (w5217, w5106, IN55[14], w5218, w5219);
  FullAdder U783 (w5219, w5108, IN56[14], w5220, w5221);
  FullAdder U784 (w5221, w5110, IN57[14], w5222, w5223);
  FullAdder U785 (w5223, w5112, IN58[12], w5224, w5225);
  FullAdder U786 (w5225, w5114, IN59[11], w5226, w5227);
  FullAdder U787 (w5227, w5116, IN60[10], w5228, w5229);
  FullAdder U788 (w5229, w5118, IN61[9], w5230, w5231);
  FullAdder U789 (w5231, w5120, IN62[8], w5232, w5233);
  FullAdder U790 (w5233, w5122, IN63[7], w5234, w5235);
  FullAdder U791 (w5235, w5124, IN64[6], w5236, w5237);
  FullAdder U792 (w5237, w5126, IN65[5], w5238, w5239);
  FullAdder U793 (w5239, w5128, IN66[4], w5240, w5241);
  FullAdder U794 (w5241, w5130, IN67[3], w5242, w5243);
  FullAdder U795 (w5243, w5132, IN68[2], w5244, w5245);
  FullAdder U796 (w5245, w5134, IN69[1], w5246, w5247);
  FullAdder U797 (w5247, w5135, IN70[0], w5248, w5249);
  HalfAdder U798 (w5138, IN15[15], Out1[15], w5251);
  FullAdder U799 (w5251, w5140, IN16[15], w5252, w5253);
  FullAdder U800 (w5253, w5142, IN17[15], w5254, w5255);
  FullAdder U801 (w5255, w5144, IN18[15], w5256, w5257);
  FullAdder U802 (w5257, w5146, IN19[15], w5258, w5259);
  FullAdder U803 (w5259, w5148, IN20[15], w5260, w5261);
  FullAdder U804 (w5261, w5150, IN21[15], w5262, w5263);
  FullAdder U805 (w5263, w5152, IN22[15], w5264, w5265);
  FullAdder U806 (w5265, w5154, IN23[15], w5266, w5267);
  FullAdder U807 (w5267, w5156, IN24[15], w5268, w5269);
  FullAdder U808 (w5269, w5158, IN25[15], w5270, w5271);
  FullAdder U809 (w5271, w5160, IN26[15], w5272, w5273);
  FullAdder U810 (w5273, w5162, IN27[15], w5274, w5275);
  FullAdder U811 (w5275, w5164, IN28[15], w5276, w5277);
  FullAdder U812 (w5277, w5166, IN29[15], w5278, w5279);
  FullAdder U813 (w5279, w5168, IN30[15], w5280, w5281);
  FullAdder U814 (w5281, w5170, IN31[15], w5282, w5283);
  FullAdder U815 (w5283, w5172, IN32[15], w5284, w5285);
  FullAdder U816 (w5285, w5174, IN33[15], w5286, w5287);
  FullAdder U817 (w5287, w5176, IN34[15], w5288, w5289);
  FullAdder U818 (w5289, w5178, IN35[15], w5290, w5291);
  FullAdder U819 (w5291, w5180, IN36[15], w5292, w5293);
  FullAdder U820 (w5293, w5182, IN37[15], w5294, w5295);
  FullAdder U821 (w5295, w5184, IN38[15], w5296, w5297);
  FullAdder U822 (w5297, w5186, IN39[15], w5298, w5299);
  FullAdder U823 (w5299, w5188, IN40[15], w5300, w5301);
  FullAdder U824 (w5301, w5190, IN41[15], w5302, w5303);
  FullAdder U825 (w5303, w5192, IN42[15], w5304, w5305);
  FullAdder U826 (w5305, w5194, IN43[15], w5306, w5307);
  FullAdder U827 (w5307, w5196, IN44[15], w5308, w5309);
  FullAdder U828 (w5309, w5198, IN45[15], w5310, w5311);
  FullAdder U829 (w5311, w5200, IN46[15], w5312, w5313);
  FullAdder U830 (w5313, w5202, IN47[15], w5314, w5315);
  FullAdder U831 (w5315, w5204, IN48[15], w5316, w5317);
  FullAdder U832 (w5317, w5206, IN49[15], w5318, w5319);
  FullAdder U833 (w5319, w5208, IN50[15], w5320, w5321);
  FullAdder U834 (w5321, w5210, IN51[15], w5322, w5323);
  FullAdder U835 (w5323, w5212, IN52[15], w5324, w5325);
  FullAdder U836 (w5325, w5214, IN53[15], w5326, w5327);
  FullAdder U837 (w5327, w5216, IN54[15], w5328, w5329);
  FullAdder U838 (w5329, w5218, IN55[15], w5330, w5331);
  FullAdder U839 (w5331, w5220, IN56[15], w5332, w5333);
  FullAdder U840 (w5333, w5222, IN57[15], w5334, w5335);
  FullAdder U841 (w5335, w5224, IN58[13], w5336, w5337);
  FullAdder U842 (w5337, w5226, IN59[12], w5338, w5339);
  FullAdder U843 (w5339, w5228, IN60[11], w5340, w5341);
  FullAdder U844 (w5341, w5230, IN61[10], w5342, w5343);
  FullAdder U845 (w5343, w5232, IN62[9], w5344, w5345);
  FullAdder U846 (w5345, w5234, IN63[8], w5346, w5347);
  FullAdder U847 (w5347, w5236, IN64[7], w5348, w5349);
  FullAdder U848 (w5349, w5238, IN65[6], w5350, w5351);
  FullAdder U849 (w5351, w5240, IN66[5], w5352, w5353);
  FullAdder U850 (w5353, w5242, IN67[4], w5354, w5355);
  FullAdder U851 (w5355, w5244, IN68[3], w5356, w5357);
  FullAdder U852 (w5357, w5246, IN69[2], w5358, w5359);
  FullAdder U853 (w5359, w5248, IN70[1], w5360, w5361);
  FullAdder U854 (w5361, w5249, IN71[0], w5362, w5363);
  HalfAdder U855 (w5252, IN16[16], Out1[16], w5365);
  FullAdder U856 (w5365, w5254, IN17[16], w5366, w5367);
  FullAdder U857 (w5367, w5256, IN18[16], w5368, w5369);
  FullAdder U858 (w5369, w5258, IN19[16], w5370, w5371);
  FullAdder U859 (w5371, w5260, IN20[16], w5372, w5373);
  FullAdder U860 (w5373, w5262, IN21[16], w5374, w5375);
  FullAdder U861 (w5375, w5264, IN22[16], w5376, w5377);
  FullAdder U862 (w5377, w5266, IN23[16], w5378, w5379);
  FullAdder U863 (w5379, w5268, IN24[16], w5380, w5381);
  FullAdder U864 (w5381, w5270, IN25[16], w5382, w5383);
  FullAdder U865 (w5383, w5272, IN26[16], w5384, w5385);
  FullAdder U866 (w5385, w5274, IN27[16], w5386, w5387);
  FullAdder U867 (w5387, w5276, IN28[16], w5388, w5389);
  FullAdder U868 (w5389, w5278, IN29[16], w5390, w5391);
  FullAdder U869 (w5391, w5280, IN30[16], w5392, w5393);
  FullAdder U870 (w5393, w5282, IN31[16], w5394, w5395);
  FullAdder U871 (w5395, w5284, IN32[16], w5396, w5397);
  FullAdder U872 (w5397, w5286, IN33[16], w5398, w5399);
  FullAdder U873 (w5399, w5288, IN34[16], w5400, w5401);
  FullAdder U874 (w5401, w5290, IN35[16], w5402, w5403);
  FullAdder U875 (w5403, w5292, IN36[16], w5404, w5405);
  FullAdder U876 (w5405, w5294, IN37[16], w5406, w5407);
  FullAdder U877 (w5407, w5296, IN38[16], w5408, w5409);
  FullAdder U878 (w5409, w5298, IN39[16], w5410, w5411);
  FullAdder U879 (w5411, w5300, IN40[16], w5412, w5413);
  FullAdder U880 (w5413, w5302, IN41[16], w5414, w5415);
  FullAdder U881 (w5415, w5304, IN42[16], w5416, w5417);
  FullAdder U882 (w5417, w5306, IN43[16], w5418, w5419);
  FullAdder U883 (w5419, w5308, IN44[16], w5420, w5421);
  FullAdder U884 (w5421, w5310, IN45[16], w5422, w5423);
  FullAdder U885 (w5423, w5312, IN46[16], w5424, w5425);
  FullAdder U886 (w5425, w5314, IN47[16], w5426, w5427);
  FullAdder U887 (w5427, w5316, IN48[16], w5428, w5429);
  FullAdder U888 (w5429, w5318, IN49[16], w5430, w5431);
  FullAdder U889 (w5431, w5320, IN50[16], w5432, w5433);
  FullAdder U890 (w5433, w5322, IN51[16], w5434, w5435);
  FullAdder U891 (w5435, w5324, IN52[16], w5436, w5437);
  FullAdder U892 (w5437, w5326, IN53[16], w5438, w5439);
  FullAdder U893 (w5439, w5328, IN54[16], w5440, w5441);
  FullAdder U894 (w5441, w5330, IN55[16], w5442, w5443);
  FullAdder U895 (w5443, w5332, IN56[16], w5444, w5445);
  FullAdder U896 (w5445, w5334, IN57[16], w5446, w5447);
  FullAdder U897 (w5447, w5336, IN58[14], w5448, w5449);
  FullAdder U898 (w5449, w5338, IN59[13], w5450, w5451);
  FullAdder U899 (w5451, w5340, IN60[12], w5452, w5453);
  FullAdder U900 (w5453, w5342, IN61[11], w5454, w5455);
  FullAdder U901 (w5455, w5344, IN62[10], w5456, w5457);
  FullAdder U902 (w5457, w5346, IN63[9], w5458, w5459);
  FullAdder U903 (w5459, w5348, IN64[8], w5460, w5461);
  FullAdder U904 (w5461, w5350, IN65[7], w5462, w5463);
  FullAdder U905 (w5463, w5352, IN66[6], w5464, w5465);
  FullAdder U906 (w5465, w5354, IN67[5], w5466, w5467);
  FullAdder U907 (w5467, w5356, IN68[4], w5468, w5469);
  FullAdder U908 (w5469, w5358, IN69[3], w5470, w5471);
  FullAdder U909 (w5471, w5360, IN70[2], w5472, w5473);
  FullAdder U910 (w5473, w5362, IN71[1], w5474, w5475);
  FullAdder U911 (w5475, w5363, IN72[0], w5476, w5477);
  HalfAdder U912 (w5366, IN17[17], Out1[17], w5479);
  FullAdder U913 (w5479, w5368, IN18[17], w5480, w5481);
  FullAdder U914 (w5481, w5370, IN19[17], w5482, w5483);
  FullAdder U915 (w5483, w5372, IN20[17], w5484, w5485);
  FullAdder U916 (w5485, w5374, IN21[17], w5486, w5487);
  FullAdder U917 (w5487, w5376, IN22[17], w5488, w5489);
  FullAdder U918 (w5489, w5378, IN23[17], w5490, w5491);
  FullAdder U919 (w5491, w5380, IN24[17], w5492, w5493);
  FullAdder U920 (w5493, w5382, IN25[17], w5494, w5495);
  FullAdder U921 (w5495, w5384, IN26[17], w5496, w5497);
  FullAdder U922 (w5497, w5386, IN27[17], w5498, w5499);
  FullAdder U923 (w5499, w5388, IN28[17], w5500, w5501);
  FullAdder U924 (w5501, w5390, IN29[17], w5502, w5503);
  FullAdder U925 (w5503, w5392, IN30[17], w5504, w5505);
  FullAdder U926 (w5505, w5394, IN31[17], w5506, w5507);
  FullAdder U927 (w5507, w5396, IN32[17], w5508, w5509);
  FullAdder U928 (w5509, w5398, IN33[17], w5510, w5511);
  FullAdder U929 (w5511, w5400, IN34[17], w5512, w5513);
  FullAdder U930 (w5513, w5402, IN35[17], w5514, w5515);
  FullAdder U931 (w5515, w5404, IN36[17], w5516, w5517);
  FullAdder U932 (w5517, w5406, IN37[17], w5518, w5519);
  FullAdder U933 (w5519, w5408, IN38[17], w5520, w5521);
  FullAdder U934 (w5521, w5410, IN39[17], w5522, w5523);
  FullAdder U935 (w5523, w5412, IN40[17], w5524, w5525);
  FullAdder U936 (w5525, w5414, IN41[17], w5526, w5527);
  FullAdder U937 (w5527, w5416, IN42[17], w5528, w5529);
  FullAdder U938 (w5529, w5418, IN43[17], w5530, w5531);
  FullAdder U939 (w5531, w5420, IN44[17], w5532, w5533);
  FullAdder U940 (w5533, w5422, IN45[17], w5534, w5535);
  FullAdder U941 (w5535, w5424, IN46[17], w5536, w5537);
  FullAdder U942 (w5537, w5426, IN47[17], w5538, w5539);
  FullAdder U943 (w5539, w5428, IN48[17], w5540, w5541);
  FullAdder U944 (w5541, w5430, IN49[17], w5542, w5543);
  FullAdder U945 (w5543, w5432, IN50[17], w5544, w5545);
  FullAdder U946 (w5545, w5434, IN51[17], w5546, w5547);
  FullAdder U947 (w5547, w5436, IN52[17], w5548, w5549);
  FullAdder U948 (w5549, w5438, IN53[17], w5550, w5551);
  FullAdder U949 (w5551, w5440, IN54[17], w5552, w5553);
  FullAdder U950 (w5553, w5442, IN55[17], w5554, w5555);
  FullAdder U951 (w5555, w5444, IN56[17], w5556, w5557);
  FullAdder U952 (w5557, w5446, IN57[17], w5558, w5559);
  FullAdder U953 (w5559, w5448, IN58[15], w5560, w5561);
  FullAdder U954 (w5561, w5450, IN59[14], w5562, w5563);
  FullAdder U955 (w5563, w5452, IN60[13], w5564, w5565);
  FullAdder U956 (w5565, w5454, IN61[12], w5566, w5567);
  FullAdder U957 (w5567, w5456, IN62[11], w5568, w5569);
  FullAdder U958 (w5569, w5458, IN63[10], w5570, w5571);
  FullAdder U959 (w5571, w5460, IN64[9], w5572, w5573);
  FullAdder U960 (w5573, w5462, IN65[8], w5574, w5575);
  FullAdder U961 (w5575, w5464, IN66[7], w5576, w5577);
  FullAdder U962 (w5577, w5466, IN67[6], w5578, w5579);
  FullAdder U963 (w5579, w5468, IN68[5], w5580, w5581);
  FullAdder U964 (w5581, w5470, IN69[4], w5582, w5583);
  FullAdder U965 (w5583, w5472, IN70[3], w5584, w5585);
  FullAdder U966 (w5585, w5474, IN71[2], w5586, w5587);
  FullAdder U967 (w5587, w5476, IN72[1], w5588, w5589);
  FullAdder U968 (w5589, w5477, IN73[0], w5590, w5591);
  HalfAdder U969 (w5480, IN18[18], Out1[18], w5593);
  FullAdder U970 (w5593, w5482, IN19[18], w5594, w5595);
  FullAdder U971 (w5595, w5484, IN20[18], w5596, w5597);
  FullAdder U972 (w5597, w5486, IN21[18], w5598, w5599);
  FullAdder U973 (w5599, w5488, IN22[18], w5600, w5601);
  FullAdder U974 (w5601, w5490, IN23[18], w5602, w5603);
  FullAdder U975 (w5603, w5492, IN24[18], w5604, w5605);
  FullAdder U976 (w5605, w5494, IN25[18], w5606, w5607);
  FullAdder U977 (w5607, w5496, IN26[18], w5608, w5609);
  FullAdder U978 (w5609, w5498, IN27[18], w5610, w5611);
  FullAdder U979 (w5611, w5500, IN28[18], w5612, w5613);
  FullAdder U980 (w5613, w5502, IN29[18], w5614, w5615);
  FullAdder U981 (w5615, w5504, IN30[18], w5616, w5617);
  FullAdder U982 (w5617, w5506, IN31[18], w5618, w5619);
  FullAdder U983 (w5619, w5508, IN32[18], w5620, w5621);
  FullAdder U984 (w5621, w5510, IN33[18], w5622, w5623);
  FullAdder U985 (w5623, w5512, IN34[18], w5624, w5625);
  FullAdder U986 (w5625, w5514, IN35[18], w5626, w5627);
  FullAdder U987 (w5627, w5516, IN36[18], w5628, w5629);
  FullAdder U988 (w5629, w5518, IN37[18], w5630, w5631);
  FullAdder U989 (w5631, w5520, IN38[18], w5632, w5633);
  FullAdder U990 (w5633, w5522, IN39[18], w5634, w5635);
  FullAdder U991 (w5635, w5524, IN40[18], w5636, w5637);
  FullAdder U992 (w5637, w5526, IN41[18], w5638, w5639);
  FullAdder U993 (w5639, w5528, IN42[18], w5640, w5641);
  FullAdder U994 (w5641, w5530, IN43[18], w5642, w5643);
  FullAdder U995 (w5643, w5532, IN44[18], w5644, w5645);
  FullAdder U996 (w5645, w5534, IN45[18], w5646, w5647);
  FullAdder U997 (w5647, w5536, IN46[18], w5648, w5649);
  FullAdder U998 (w5649, w5538, IN47[18], w5650, w5651);
  FullAdder U999 (w5651, w5540, IN48[18], w5652, w5653);
  FullAdder U1000 (w5653, w5542, IN49[18], w5654, w5655);
  FullAdder U1001 (w5655, w5544, IN50[18], w5656, w5657);
  FullAdder U1002 (w5657, w5546, IN51[18], w5658, w5659);
  FullAdder U1003 (w5659, w5548, IN52[18], w5660, w5661);
  FullAdder U1004 (w5661, w5550, IN53[18], w5662, w5663);
  FullAdder U1005 (w5663, w5552, IN54[18], w5664, w5665);
  FullAdder U1006 (w5665, w5554, IN55[18], w5666, w5667);
  FullAdder U1007 (w5667, w5556, IN56[18], w5668, w5669);
  FullAdder U1008 (w5669, w5558, IN57[18], w5670, w5671);
  FullAdder U1009 (w5671, w5560, IN58[16], w5672, w5673);
  FullAdder U1010 (w5673, w5562, IN59[15], w5674, w5675);
  FullAdder U1011 (w5675, w5564, IN60[14], w5676, w5677);
  FullAdder U1012 (w5677, w5566, IN61[13], w5678, w5679);
  FullAdder U1013 (w5679, w5568, IN62[12], w5680, w5681);
  FullAdder U1014 (w5681, w5570, IN63[11], w5682, w5683);
  FullAdder U1015 (w5683, w5572, IN64[10], w5684, w5685);
  FullAdder U1016 (w5685, w5574, IN65[9], w5686, w5687);
  FullAdder U1017 (w5687, w5576, IN66[8], w5688, w5689);
  FullAdder U1018 (w5689, w5578, IN67[7], w5690, w5691);
  FullAdder U1019 (w5691, w5580, IN68[6], w5692, w5693);
  FullAdder U1020 (w5693, w5582, IN69[5], w5694, w5695);
  FullAdder U1021 (w5695, w5584, IN70[4], w5696, w5697);
  FullAdder U1022 (w5697, w5586, IN71[3], w5698, w5699);
  FullAdder U1023 (w5699, w5588, IN72[2], w5700, w5701);
  FullAdder U1024 (w5701, w5590, IN73[1], w5702, w5703);
  FullAdder U1025 (w5703, w5591, IN74[0], w5704, w5705);
  HalfAdder U1026 (w5594, IN19[19], Out1[19], w5707);
  FullAdder U1027 (w5707, w5596, IN20[19], w5708, w5709);
  FullAdder U1028 (w5709, w5598, IN21[19], w5710, w5711);
  FullAdder U1029 (w5711, w5600, IN22[19], w5712, w5713);
  FullAdder U1030 (w5713, w5602, IN23[19], w5714, w5715);
  FullAdder U1031 (w5715, w5604, IN24[19], w5716, w5717);
  FullAdder U1032 (w5717, w5606, IN25[19], w5718, w5719);
  FullAdder U1033 (w5719, w5608, IN26[19], w5720, w5721);
  FullAdder U1034 (w5721, w5610, IN27[19], w5722, w5723);
  FullAdder U1035 (w5723, w5612, IN28[19], w5724, w5725);
  FullAdder U1036 (w5725, w5614, IN29[19], w5726, w5727);
  FullAdder U1037 (w5727, w5616, IN30[19], w5728, w5729);
  FullAdder U1038 (w5729, w5618, IN31[19], w5730, w5731);
  FullAdder U1039 (w5731, w5620, IN32[19], w5732, w5733);
  FullAdder U1040 (w5733, w5622, IN33[19], w5734, w5735);
  FullAdder U1041 (w5735, w5624, IN34[19], w5736, w5737);
  FullAdder U1042 (w5737, w5626, IN35[19], w5738, w5739);
  FullAdder U1043 (w5739, w5628, IN36[19], w5740, w5741);
  FullAdder U1044 (w5741, w5630, IN37[19], w5742, w5743);
  FullAdder U1045 (w5743, w5632, IN38[19], w5744, w5745);
  FullAdder U1046 (w5745, w5634, IN39[19], w5746, w5747);
  FullAdder U1047 (w5747, w5636, IN40[19], w5748, w5749);
  FullAdder U1048 (w5749, w5638, IN41[19], w5750, w5751);
  FullAdder U1049 (w5751, w5640, IN42[19], w5752, w5753);
  FullAdder U1050 (w5753, w5642, IN43[19], w5754, w5755);
  FullAdder U1051 (w5755, w5644, IN44[19], w5756, w5757);
  FullAdder U1052 (w5757, w5646, IN45[19], w5758, w5759);
  FullAdder U1053 (w5759, w5648, IN46[19], w5760, w5761);
  FullAdder U1054 (w5761, w5650, IN47[19], w5762, w5763);
  FullAdder U1055 (w5763, w5652, IN48[19], w5764, w5765);
  FullAdder U1056 (w5765, w5654, IN49[19], w5766, w5767);
  FullAdder U1057 (w5767, w5656, IN50[19], w5768, w5769);
  FullAdder U1058 (w5769, w5658, IN51[19], w5770, w5771);
  FullAdder U1059 (w5771, w5660, IN52[19], w5772, w5773);
  FullAdder U1060 (w5773, w5662, IN53[19], w5774, w5775);
  FullAdder U1061 (w5775, w5664, IN54[19], w5776, w5777);
  FullAdder U1062 (w5777, w5666, IN55[19], w5778, w5779);
  FullAdder U1063 (w5779, w5668, IN56[19], w5780, w5781);
  FullAdder U1064 (w5781, w5670, IN57[19], w5782, w5783);
  FullAdder U1065 (w5783, w5672, IN58[17], w5784, w5785);
  FullAdder U1066 (w5785, w5674, IN59[16], w5786, w5787);
  FullAdder U1067 (w5787, w5676, IN60[15], w5788, w5789);
  FullAdder U1068 (w5789, w5678, IN61[14], w5790, w5791);
  FullAdder U1069 (w5791, w5680, IN62[13], w5792, w5793);
  FullAdder U1070 (w5793, w5682, IN63[12], w5794, w5795);
  FullAdder U1071 (w5795, w5684, IN64[11], w5796, w5797);
  FullAdder U1072 (w5797, w5686, IN65[10], w5798, w5799);
  FullAdder U1073 (w5799, w5688, IN66[9], w5800, w5801);
  FullAdder U1074 (w5801, w5690, IN67[8], w5802, w5803);
  FullAdder U1075 (w5803, w5692, IN68[7], w5804, w5805);
  FullAdder U1076 (w5805, w5694, IN69[6], w5806, w5807);
  FullAdder U1077 (w5807, w5696, IN70[5], w5808, w5809);
  FullAdder U1078 (w5809, w5698, IN71[4], w5810, w5811);
  FullAdder U1079 (w5811, w5700, IN72[3], w5812, w5813);
  FullAdder U1080 (w5813, w5702, IN73[2], w5814, w5815);
  FullAdder U1081 (w5815, w5704, IN74[1], w5816, w5817);
  FullAdder U1082 (w5817, w5705, IN75[0], w5818, w5819);
  HalfAdder U1083 (w5708, IN20[20], Out1[20], w5821);
  FullAdder U1084 (w5821, w5710, IN21[20], w5822, w5823);
  FullAdder U1085 (w5823, w5712, IN22[20], w5824, w5825);
  FullAdder U1086 (w5825, w5714, IN23[20], w5826, w5827);
  FullAdder U1087 (w5827, w5716, IN24[20], w5828, w5829);
  FullAdder U1088 (w5829, w5718, IN25[20], w5830, w5831);
  FullAdder U1089 (w5831, w5720, IN26[20], w5832, w5833);
  FullAdder U1090 (w5833, w5722, IN27[20], w5834, w5835);
  FullAdder U1091 (w5835, w5724, IN28[20], w5836, w5837);
  FullAdder U1092 (w5837, w5726, IN29[20], w5838, w5839);
  FullAdder U1093 (w5839, w5728, IN30[20], w5840, w5841);
  FullAdder U1094 (w5841, w5730, IN31[20], w5842, w5843);
  FullAdder U1095 (w5843, w5732, IN32[20], w5844, w5845);
  FullAdder U1096 (w5845, w5734, IN33[20], w5846, w5847);
  FullAdder U1097 (w5847, w5736, IN34[20], w5848, w5849);
  FullAdder U1098 (w5849, w5738, IN35[20], w5850, w5851);
  FullAdder U1099 (w5851, w5740, IN36[20], w5852, w5853);
  FullAdder U1100 (w5853, w5742, IN37[20], w5854, w5855);
  FullAdder U1101 (w5855, w5744, IN38[20], w5856, w5857);
  FullAdder U1102 (w5857, w5746, IN39[20], w5858, w5859);
  FullAdder U1103 (w5859, w5748, IN40[20], w5860, w5861);
  FullAdder U1104 (w5861, w5750, IN41[20], w5862, w5863);
  FullAdder U1105 (w5863, w5752, IN42[20], w5864, w5865);
  FullAdder U1106 (w5865, w5754, IN43[20], w5866, w5867);
  FullAdder U1107 (w5867, w5756, IN44[20], w5868, w5869);
  FullAdder U1108 (w5869, w5758, IN45[20], w5870, w5871);
  FullAdder U1109 (w5871, w5760, IN46[20], w5872, w5873);
  FullAdder U1110 (w5873, w5762, IN47[20], w5874, w5875);
  FullAdder U1111 (w5875, w5764, IN48[20], w5876, w5877);
  FullAdder U1112 (w5877, w5766, IN49[20], w5878, w5879);
  FullAdder U1113 (w5879, w5768, IN50[20], w5880, w5881);
  FullAdder U1114 (w5881, w5770, IN51[20], w5882, w5883);
  FullAdder U1115 (w5883, w5772, IN52[20], w5884, w5885);
  FullAdder U1116 (w5885, w5774, IN53[20], w5886, w5887);
  FullAdder U1117 (w5887, w5776, IN54[20], w5888, w5889);
  FullAdder U1118 (w5889, w5778, IN55[20], w5890, w5891);
  FullAdder U1119 (w5891, w5780, IN56[20], w5892, w5893);
  FullAdder U1120 (w5893, w5782, IN57[20], w5894, w5895);
  FullAdder U1121 (w5895, w5784, IN58[18], w5896, w5897);
  FullAdder U1122 (w5897, w5786, IN59[17], w5898, w5899);
  FullAdder U1123 (w5899, w5788, IN60[16], w5900, w5901);
  FullAdder U1124 (w5901, w5790, IN61[15], w5902, w5903);
  FullAdder U1125 (w5903, w5792, IN62[14], w5904, w5905);
  FullAdder U1126 (w5905, w5794, IN63[13], w5906, w5907);
  FullAdder U1127 (w5907, w5796, IN64[12], w5908, w5909);
  FullAdder U1128 (w5909, w5798, IN65[11], w5910, w5911);
  FullAdder U1129 (w5911, w5800, IN66[10], w5912, w5913);
  FullAdder U1130 (w5913, w5802, IN67[9], w5914, w5915);
  FullAdder U1131 (w5915, w5804, IN68[8], w5916, w5917);
  FullAdder U1132 (w5917, w5806, IN69[7], w5918, w5919);
  FullAdder U1133 (w5919, w5808, IN70[6], w5920, w5921);
  FullAdder U1134 (w5921, w5810, IN71[5], w5922, w5923);
  FullAdder U1135 (w5923, w5812, IN72[4], w5924, w5925);
  FullAdder U1136 (w5925, w5814, IN73[3], w5926, w5927);
  FullAdder U1137 (w5927, w5816, IN74[2], w5928, w5929);
  FullAdder U1138 (w5929, w5818, IN75[1], w5930, w5931);
  FullAdder U1139 (w5931, w5819, IN76[0], w5932, w5933);
  HalfAdder U1140 (w5822, IN21[21], Out1[21], w5935);
  FullAdder U1141 (w5935, w5824, IN22[21], w5936, w5937);
  FullAdder U1142 (w5937, w5826, IN23[21], w5938, w5939);
  FullAdder U1143 (w5939, w5828, IN24[21], w5940, w5941);
  FullAdder U1144 (w5941, w5830, IN25[21], w5942, w5943);
  FullAdder U1145 (w5943, w5832, IN26[21], w5944, w5945);
  FullAdder U1146 (w5945, w5834, IN27[21], w5946, w5947);
  FullAdder U1147 (w5947, w5836, IN28[21], w5948, w5949);
  FullAdder U1148 (w5949, w5838, IN29[21], w5950, w5951);
  FullAdder U1149 (w5951, w5840, IN30[21], w5952, w5953);
  FullAdder U1150 (w5953, w5842, IN31[21], w5954, w5955);
  FullAdder U1151 (w5955, w5844, IN32[21], w5956, w5957);
  FullAdder U1152 (w5957, w5846, IN33[21], w5958, w5959);
  FullAdder U1153 (w5959, w5848, IN34[21], w5960, w5961);
  FullAdder U1154 (w5961, w5850, IN35[21], w5962, w5963);
  FullAdder U1155 (w5963, w5852, IN36[21], w5964, w5965);
  FullAdder U1156 (w5965, w5854, IN37[21], w5966, w5967);
  FullAdder U1157 (w5967, w5856, IN38[21], w5968, w5969);
  FullAdder U1158 (w5969, w5858, IN39[21], w5970, w5971);
  FullAdder U1159 (w5971, w5860, IN40[21], w5972, w5973);
  FullAdder U1160 (w5973, w5862, IN41[21], w5974, w5975);
  FullAdder U1161 (w5975, w5864, IN42[21], w5976, w5977);
  FullAdder U1162 (w5977, w5866, IN43[21], w5978, w5979);
  FullAdder U1163 (w5979, w5868, IN44[21], w5980, w5981);
  FullAdder U1164 (w5981, w5870, IN45[21], w5982, w5983);
  FullAdder U1165 (w5983, w5872, IN46[21], w5984, w5985);
  FullAdder U1166 (w5985, w5874, IN47[21], w5986, w5987);
  FullAdder U1167 (w5987, w5876, IN48[21], w5988, w5989);
  FullAdder U1168 (w5989, w5878, IN49[21], w5990, w5991);
  FullAdder U1169 (w5991, w5880, IN50[21], w5992, w5993);
  FullAdder U1170 (w5993, w5882, IN51[21], w5994, w5995);
  FullAdder U1171 (w5995, w5884, IN52[21], w5996, w5997);
  FullAdder U1172 (w5997, w5886, IN53[21], w5998, w5999);
  FullAdder U1173 (w5999, w5888, IN54[21], w6000, w6001);
  FullAdder U1174 (w6001, w5890, IN55[21], w6002, w6003);
  FullAdder U1175 (w6003, w5892, IN56[21], w6004, w6005);
  FullAdder U1176 (w6005, w5894, IN57[21], w6006, w6007);
  FullAdder U1177 (w6007, w5896, IN58[19], w6008, w6009);
  FullAdder U1178 (w6009, w5898, IN59[18], w6010, w6011);
  FullAdder U1179 (w6011, w5900, IN60[17], w6012, w6013);
  FullAdder U1180 (w6013, w5902, IN61[16], w6014, w6015);
  FullAdder U1181 (w6015, w5904, IN62[15], w6016, w6017);
  FullAdder U1182 (w6017, w5906, IN63[14], w6018, w6019);
  FullAdder U1183 (w6019, w5908, IN64[13], w6020, w6021);
  FullAdder U1184 (w6021, w5910, IN65[12], w6022, w6023);
  FullAdder U1185 (w6023, w5912, IN66[11], w6024, w6025);
  FullAdder U1186 (w6025, w5914, IN67[10], w6026, w6027);
  FullAdder U1187 (w6027, w5916, IN68[9], w6028, w6029);
  FullAdder U1188 (w6029, w5918, IN69[8], w6030, w6031);
  FullAdder U1189 (w6031, w5920, IN70[7], w6032, w6033);
  FullAdder U1190 (w6033, w5922, IN71[6], w6034, w6035);
  FullAdder U1191 (w6035, w5924, IN72[5], w6036, w6037);
  FullAdder U1192 (w6037, w5926, IN73[4], w6038, w6039);
  FullAdder U1193 (w6039, w5928, IN74[3], w6040, w6041);
  FullAdder U1194 (w6041, w5930, IN75[2], w6042, w6043);
  FullAdder U1195 (w6043, w5932, IN76[1], w6044, w6045);
  FullAdder U1196 (w6045, w5933, IN77[0], w6046, w6047);
  HalfAdder U1197 (w5936, IN22[22], Out1[22], w6049);
  FullAdder U1198 (w6049, w5938, IN23[22], w6050, w6051);
  FullAdder U1199 (w6051, w5940, IN24[22], w6052, w6053);
  FullAdder U1200 (w6053, w5942, IN25[22], w6054, w6055);
  FullAdder U1201 (w6055, w5944, IN26[22], w6056, w6057);
  FullAdder U1202 (w6057, w5946, IN27[22], w6058, w6059);
  FullAdder U1203 (w6059, w5948, IN28[22], w6060, w6061);
  FullAdder U1204 (w6061, w5950, IN29[22], w6062, w6063);
  FullAdder U1205 (w6063, w5952, IN30[22], w6064, w6065);
  FullAdder U1206 (w6065, w5954, IN31[22], w6066, w6067);
  FullAdder U1207 (w6067, w5956, IN32[22], w6068, w6069);
  FullAdder U1208 (w6069, w5958, IN33[22], w6070, w6071);
  FullAdder U1209 (w6071, w5960, IN34[22], w6072, w6073);
  FullAdder U1210 (w6073, w5962, IN35[22], w6074, w6075);
  FullAdder U1211 (w6075, w5964, IN36[22], w6076, w6077);
  FullAdder U1212 (w6077, w5966, IN37[22], w6078, w6079);
  FullAdder U1213 (w6079, w5968, IN38[22], w6080, w6081);
  FullAdder U1214 (w6081, w5970, IN39[22], w6082, w6083);
  FullAdder U1215 (w6083, w5972, IN40[22], w6084, w6085);
  FullAdder U1216 (w6085, w5974, IN41[22], w6086, w6087);
  FullAdder U1217 (w6087, w5976, IN42[22], w6088, w6089);
  FullAdder U1218 (w6089, w5978, IN43[22], w6090, w6091);
  FullAdder U1219 (w6091, w5980, IN44[22], w6092, w6093);
  FullAdder U1220 (w6093, w5982, IN45[22], w6094, w6095);
  FullAdder U1221 (w6095, w5984, IN46[22], w6096, w6097);
  FullAdder U1222 (w6097, w5986, IN47[22], w6098, w6099);
  FullAdder U1223 (w6099, w5988, IN48[22], w6100, w6101);
  FullAdder U1224 (w6101, w5990, IN49[22], w6102, w6103);
  FullAdder U1225 (w6103, w5992, IN50[22], w6104, w6105);
  FullAdder U1226 (w6105, w5994, IN51[22], w6106, w6107);
  FullAdder U1227 (w6107, w5996, IN52[22], w6108, w6109);
  FullAdder U1228 (w6109, w5998, IN53[22], w6110, w6111);
  FullAdder U1229 (w6111, w6000, IN54[22], w6112, w6113);
  FullAdder U1230 (w6113, w6002, IN55[22], w6114, w6115);
  FullAdder U1231 (w6115, w6004, IN56[22], w6116, w6117);
  FullAdder U1232 (w6117, w6006, IN57[22], w6118, w6119);
  FullAdder U1233 (w6119, w6008, IN58[20], w6120, w6121);
  FullAdder U1234 (w6121, w6010, IN59[19], w6122, w6123);
  FullAdder U1235 (w6123, w6012, IN60[18], w6124, w6125);
  FullAdder U1236 (w6125, w6014, IN61[17], w6126, w6127);
  FullAdder U1237 (w6127, w6016, IN62[16], w6128, w6129);
  FullAdder U1238 (w6129, w6018, IN63[15], w6130, w6131);
  FullAdder U1239 (w6131, w6020, IN64[14], w6132, w6133);
  FullAdder U1240 (w6133, w6022, IN65[13], w6134, w6135);
  FullAdder U1241 (w6135, w6024, IN66[12], w6136, w6137);
  FullAdder U1242 (w6137, w6026, IN67[11], w6138, w6139);
  FullAdder U1243 (w6139, w6028, IN68[10], w6140, w6141);
  FullAdder U1244 (w6141, w6030, IN69[9], w6142, w6143);
  FullAdder U1245 (w6143, w6032, IN70[8], w6144, w6145);
  FullAdder U1246 (w6145, w6034, IN71[7], w6146, w6147);
  FullAdder U1247 (w6147, w6036, IN72[6], w6148, w6149);
  FullAdder U1248 (w6149, w6038, IN73[5], w6150, w6151);
  FullAdder U1249 (w6151, w6040, IN74[4], w6152, w6153);
  FullAdder U1250 (w6153, w6042, IN75[3], w6154, w6155);
  FullAdder U1251 (w6155, w6044, IN76[2], w6156, w6157);
  FullAdder U1252 (w6157, w6046, IN77[1], w6158, w6159);
  FullAdder U1253 (w6159, w6047, IN78[0], w6160, w6161);
  HalfAdder U1254 (w6050, IN23[23], Out1[23], w6163);
  FullAdder U1255 (w6163, w6052, IN24[23], w6164, w6165);
  FullAdder U1256 (w6165, w6054, IN25[23], w6166, w6167);
  FullAdder U1257 (w6167, w6056, IN26[23], w6168, w6169);
  FullAdder U1258 (w6169, w6058, IN27[23], w6170, w6171);
  FullAdder U1259 (w6171, w6060, IN28[23], w6172, w6173);
  FullAdder U1260 (w6173, w6062, IN29[23], w6174, w6175);
  FullAdder U1261 (w6175, w6064, IN30[23], w6176, w6177);
  FullAdder U1262 (w6177, w6066, IN31[23], w6178, w6179);
  FullAdder U1263 (w6179, w6068, IN32[23], w6180, w6181);
  FullAdder U1264 (w6181, w6070, IN33[23], w6182, w6183);
  FullAdder U1265 (w6183, w6072, IN34[23], w6184, w6185);
  FullAdder U1266 (w6185, w6074, IN35[23], w6186, w6187);
  FullAdder U1267 (w6187, w6076, IN36[23], w6188, w6189);
  FullAdder U1268 (w6189, w6078, IN37[23], w6190, w6191);
  FullAdder U1269 (w6191, w6080, IN38[23], w6192, w6193);
  FullAdder U1270 (w6193, w6082, IN39[23], w6194, w6195);
  FullAdder U1271 (w6195, w6084, IN40[23], w6196, w6197);
  FullAdder U1272 (w6197, w6086, IN41[23], w6198, w6199);
  FullAdder U1273 (w6199, w6088, IN42[23], w6200, w6201);
  FullAdder U1274 (w6201, w6090, IN43[23], w6202, w6203);
  FullAdder U1275 (w6203, w6092, IN44[23], w6204, w6205);
  FullAdder U1276 (w6205, w6094, IN45[23], w6206, w6207);
  FullAdder U1277 (w6207, w6096, IN46[23], w6208, w6209);
  FullAdder U1278 (w6209, w6098, IN47[23], w6210, w6211);
  FullAdder U1279 (w6211, w6100, IN48[23], w6212, w6213);
  FullAdder U1280 (w6213, w6102, IN49[23], w6214, w6215);
  FullAdder U1281 (w6215, w6104, IN50[23], w6216, w6217);
  FullAdder U1282 (w6217, w6106, IN51[23], w6218, w6219);
  FullAdder U1283 (w6219, w6108, IN52[23], w6220, w6221);
  FullAdder U1284 (w6221, w6110, IN53[23], w6222, w6223);
  FullAdder U1285 (w6223, w6112, IN54[23], w6224, w6225);
  FullAdder U1286 (w6225, w6114, IN55[23], w6226, w6227);
  FullAdder U1287 (w6227, w6116, IN56[23], w6228, w6229);
  FullAdder U1288 (w6229, w6118, IN57[23], w6230, w6231);
  FullAdder U1289 (w6231, w6120, IN58[21], w6232, w6233);
  FullAdder U1290 (w6233, w6122, IN59[20], w6234, w6235);
  FullAdder U1291 (w6235, w6124, IN60[19], w6236, w6237);
  FullAdder U1292 (w6237, w6126, IN61[18], w6238, w6239);
  FullAdder U1293 (w6239, w6128, IN62[17], w6240, w6241);
  FullAdder U1294 (w6241, w6130, IN63[16], w6242, w6243);
  FullAdder U1295 (w6243, w6132, IN64[15], w6244, w6245);
  FullAdder U1296 (w6245, w6134, IN65[14], w6246, w6247);
  FullAdder U1297 (w6247, w6136, IN66[13], w6248, w6249);
  FullAdder U1298 (w6249, w6138, IN67[12], w6250, w6251);
  FullAdder U1299 (w6251, w6140, IN68[11], w6252, w6253);
  FullAdder U1300 (w6253, w6142, IN69[10], w6254, w6255);
  FullAdder U1301 (w6255, w6144, IN70[9], w6256, w6257);
  FullAdder U1302 (w6257, w6146, IN71[8], w6258, w6259);
  FullAdder U1303 (w6259, w6148, IN72[7], w6260, w6261);
  FullAdder U1304 (w6261, w6150, IN73[6], w6262, w6263);
  FullAdder U1305 (w6263, w6152, IN74[5], w6264, w6265);
  FullAdder U1306 (w6265, w6154, IN75[4], w6266, w6267);
  FullAdder U1307 (w6267, w6156, IN76[3], w6268, w6269);
  FullAdder U1308 (w6269, w6158, IN77[2], w6270, w6271);
  FullAdder U1309 (w6271, w6160, IN78[1], w6272, w6273);
  FullAdder U1310 (w6273, w6161, IN79[0], w6274, w6275);
  HalfAdder U1311 (w6164, IN24[24], Out1[24], w6277);
  FullAdder U1312 (w6277, w6166, IN25[24], w6278, w6279);
  FullAdder U1313 (w6279, w6168, IN26[24], w6280, w6281);
  FullAdder U1314 (w6281, w6170, IN27[24], w6282, w6283);
  FullAdder U1315 (w6283, w6172, IN28[24], w6284, w6285);
  FullAdder U1316 (w6285, w6174, IN29[24], w6286, w6287);
  FullAdder U1317 (w6287, w6176, IN30[24], w6288, w6289);
  FullAdder U1318 (w6289, w6178, IN31[24], w6290, w6291);
  FullAdder U1319 (w6291, w6180, IN32[24], w6292, w6293);
  FullAdder U1320 (w6293, w6182, IN33[24], w6294, w6295);
  FullAdder U1321 (w6295, w6184, IN34[24], w6296, w6297);
  FullAdder U1322 (w6297, w6186, IN35[24], w6298, w6299);
  FullAdder U1323 (w6299, w6188, IN36[24], w6300, w6301);
  FullAdder U1324 (w6301, w6190, IN37[24], w6302, w6303);
  FullAdder U1325 (w6303, w6192, IN38[24], w6304, w6305);
  FullAdder U1326 (w6305, w6194, IN39[24], w6306, w6307);
  FullAdder U1327 (w6307, w6196, IN40[24], w6308, w6309);
  FullAdder U1328 (w6309, w6198, IN41[24], w6310, w6311);
  FullAdder U1329 (w6311, w6200, IN42[24], w6312, w6313);
  FullAdder U1330 (w6313, w6202, IN43[24], w6314, w6315);
  FullAdder U1331 (w6315, w6204, IN44[24], w6316, w6317);
  FullAdder U1332 (w6317, w6206, IN45[24], w6318, w6319);
  FullAdder U1333 (w6319, w6208, IN46[24], w6320, w6321);
  FullAdder U1334 (w6321, w6210, IN47[24], w6322, w6323);
  FullAdder U1335 (w6323, w6212, IN48[24], w6324, w6325);
  FullAdder U1336 (w6325, w6214, IN49[24], w6326, w6327);
  FullAdder U1337 (w6327, w6216, IN50[24], w6328, w6329);
  FullAdder U1338 (w6329, w6218, IN51[24], w6330, w6331);
  FullAdder U1339 (w6331, w6220, IN52[24], w6332, w6333);
  FullAdder U1340 (w6333, w6222, IN53[24], w6334, w6335);
  FullAdder U1341 (w6335, w6224, IN54[24], w6336, w6337);
  FullAdder U1342 (w6337, w6226, IN55[24], w6338, w6339);
  FullAdder U1343 (w6339, w6228, IN56[24], w6340, w6341);
  FullAdder U1344 (w6341, w6230, IN57[24], w6342, w6343);
  FullAdder U1345 (w6343, w6232, IN58[22], w6344, w6345);
  FullAdder U1346 (w6345, w6234, IN59[21], w6346, w6347);
  FullAdder U1347 (w6347, w6236, IN60[20], w6348, w6349);
  FullAdder U1348 (w6349, w6238, IN61[19], w6350, w6351);
  FullAdder U1349 (w6351, w6240, IN62[18], w6352, w6353);
  FullAdder U1350 (w6353, w6242, IN63[17], w6354, w6355);
  FullAdder U1351 (w6355, w6244, IN64[16], w6356, w6357);
  FullAdder U1352 (w6357, w6246, IN65[15], w6358, w6359);
  FullAdder U1353 (w6359, w6248, IN66[14], w6360, w6361);
  FullAdder U1354 (w6361, w6250, IN67[13], w6362, w6363);
  FullAdder U1355 (w6363, w6252, IN68[12], w6364, w6365);
  FullAdder U1356 (w6365, w6254, IN69[11], w6366, w6367);
  FullAdder U1357 (w6367, w6256, IN70[10], w6368, w6369);
  FullAdder U1358 (w6369, w6258, IN71[9], w6370, w6371);
  FullAdder U1359 (w6371, w6260, IN72[8], w6372, w6373);
  FullAdder U1360 (w6373, w6262, IN73[7], w6374, w6375);
  FullAdder U1361 (w6375, w6264, IN74[6], w6376, w6377);
  FullAdder U1362 (w6377, w6266, IN75[5], w6378, w6379);
  FullAdder U1363 (w6379, w6268, IN76[4], w6380, w6381);
  FullAdder U1364 (w6381, w6270, IN77[3], w6382, w6383);
  FullAdder U1365 (w6383, w6272, IN78[2], w6384, w6385);
  FullAdder U1366 (w6385, w6274, IN79[1], w6386, w6387);
  FullAdder U1367 (w6387, w6275, IN80[0], w6388, w6389);
  HalfAdder U1368 (w6278, IN25[25], Out1[25], w6391);
  FullAdder U1369 (w6391, w6280, IN26[25], w6392, w6393);
  FullAdder U1370 (w6393, w6282, IN27[25], w6394, w6395);
  FullAdder U1371 (w6395, w6284, IN28[25], w6396, w6397);
  FullAdder U1372 (w6397, w6286, IN29[25], w6398, w6399);
  FullAdder U1373 (w6399, w6288, IN30[25], w6400, w6401);
  FullAdder U1374 (w6401, w6290, IN31[25], w6402, w6403);
  FullAdder U1375 (w6403, w6292, IN32[25], w6404, w6405);
  FullAdder U1376 (w6405, w6294, IN33[25], w6406, w6407);
  FullAdder U1377 (w6407, w6296, IN34[25], w6408, w6409);
  FullAdder U1378 (w6409, w6298, IN35[25], w6410, w6411);
  FullAdder U1379 (w6411, w6300, IN36[25], w6412, w6413);
  FullAdder U1380 (w6413, w6302, IN37[25], w6414, w6415);
  FullAdder U1381 (w6415, w6304, IN38[25], w6416, w6417);
  FullAdder U1382 (w6417, w6306, IN39[25], w6418, w6419);
  FullAdder U1383 (w6419, w6308, IN40[25], w6420, w6421);
  FullAdder U1384 (w6421, w6310, IN41[25], w6422, w6423);
  FullAdder U1385 (w6423, w6312, IN42[25], w6424, w6425);
  FullAdder U1386 (w6425, w6314, IN43[25], w6426, w6427);
  FullAdder U1387 (w6427, w6316, IN44[25], w6428, w6429);
  FullAdder U1388 (w6429, w6318, IN45[25], w6430, w6431);
  FullAdder U1389 (w6431, w6320, IN46[25], w6432, w6433);
  FullAdder U1390 (w6433, w6322, IN47[25], w6434, w6435);
  FullAdder U1391 (w6435, w6324, IN48[25], w6436, w6437);
  FullAdder U1392 (w6437, w6326, IN49[25], w6438, w6439);
  FullAdder U1393 (w6439, w6328, IN50[25], w6440, w6441);
  FullAdder U1394 (w6441, w6330, IN51[25], w6442, w6443);
  FullAdder U1395 (w6443, w6332, IN52[25], w6444, w6445);
  FullAdder U1396 (w6445, w6334, IN53[25], w6446, w6447);
  FullAdder U1397 (w6447, w6336, IN54[25], w6448, w6449);
  FullAdder U1398 (w6449, w6338, IN55[25], w6450, w6451);
  FullAdder U1399 (w6451, w6340, IN56[25], w6452, w6453);
  FullAdder U1400 (w6453, w6342, IN57[25], w6454, w6455);
  FullAdder U1401 (w6455, w6344, IN58[23], w6456, w6457);
  FullAdder U1402 (w6457, w6346, IN59[22], w6458, w6459);
  FullAdder U1403 (w6459, w6348, IN60[21], w6460, w6461);
  FullAdder U1404 (w6461, w6350, IN61[20], w6462, w6463);
  FullAdder U1405 (w6463, w6352, IN62[19], w6464, w6465);
  FullAdder U1406 (w6465, w6354, IN63[18], w6466, w6467);
  FullAdder U1407 (w6467, w6356, IN64[17], w6468, w6469);
  FullAdder U1408 (w6469, w6358, IN65[16], w6470, w6471);
  FullAdder U1409 (w6471, w6360, IN66[15], w6472, w6473);
  FullAdder U1410 (w6473, w6362, IN67[14], w6474, w6475);
  FullAdder U1411 (w6475, w6364, IN68[13], w6476, w6477);
  FullAdder U1412 (w6477, w6366, IN69[12], w6478, w6479);
  FullAdder U1413 (w6479, w6368, IN70[11], w6480, w6481);
  FullAdder U1414 (w6481, w6370, IN71[10], w6482, w6483);
  FullAdder U1415 (w6483, w6372, IN72[9], w6484, w6485);
  FullAdder U1416 (w6485, w6374, IN73[8], w6486, w6487);
  FullAdder U1417 (w6487, w6376, IN74[7], w6488, w6489);
  FullAdder U1418 (w6489, w6378, IN75[6], w6490, w6491);
  FullAdder U1419 (w6491, w6380, IN76[5], w6492, w6493);
  FullAdder U1420 (w6493, w6382, IN77[4], w6494, w6495);
  FullAdder U1421 (w6495, w6384, IN78[3], w6496, w6497);
  FullAdder U1422 (w6497, w6386, IN79[2], w6498, w6499);
  FullAdder U1423 (w6499, w6388, IN80[1], w6500, w6501);
  FullAdder U1424 (w6501, w6389, IN81[0], w6502, w6503);
  HalfAdder U1425 (w6392, IN26[26], Out1[26], w6505);
  FullAdder U1426 (w6505, w6394, IN27[26], w6506, w6507);
  FullAdder U1427 (w6507, w6396, IN28[26], w6508, w6509);
  FullAdder U1428 (w6509, w6398, IN29[26], w6510, w6511);
  FullAdder U1429 (w6511, w6400, IN30[26], w6512, w6513);
  FullAdder U1430 (w6513, w6402, IN31[26], w6514, w6515);
  FullAdder U1431 (w6515, w6404, IN32[26], w6516, w6517);
  FullAdder U1432 (w6517, w6406, IN33[26], w6518, w6519);
  FullAdder U1433 (w6519, w6408, IN34[26], w6520, w6521);
  FullAdder U1434 (w6521, w6410, IN35[26], w6522, w6523);
  FullAdder U1435 (w6523, w6412, IN36[26], w6524, w6525);
  FullAdder U1436 (w6525, w6414, IN37[26], w6526, w6527);
  FullAdder U1437 (w6527, w6416, IN38[26], w6528, w6529);
  FullAdder U1438 (w6529, w6418, IN39[26], w6530, w6531);
  FullAdder U1439 (w6531, w6420, IN40[26], w6532, w6533);
  FullAdder U1440 (w6533, w6422, IN41[26], w6534, w6535);
  FullAdder U1441 (w6535, w6424, IN42[26], w6536, w6537);
  FullAdder U1442 (w6537, w6426, IN43[26], w6538, w6539);
  FullAdder U1443 (w6539, w6428, IN44[26], w6540, w6541);
  FullAdder U1444 (w6541, w6430, IN45[26], w6542, w6543);
  FullAdder U1445 (w6543, w6432, IN46[26], w6544, w6545);
  FullAdder U1446 (w6545, w6434, IN47[26], w6546, w6547);
  FullAdder U1447 (w6547, w6436, IN48[26], w6548, w6549);
  FullAdder U1448 (w6549, w6438, IN49[26], w6550, w6551);
  FullAdder U1449 (w6551, w6440, IN50[26], w6552, w6553);
  FullAdder U1450 (w6553, w6442, IN51[26], w6554, w6555);
  FullAdder U1451 (w6555, w6444, IN52[26], w6556, w6557);
  FullAdder U1452 (w6557, w6446, IN53[26], w6558, w6559);
  FullAdder U1453 (w6559, w6448, IN54[26], w6560, w6561);
  FullAdder U1454 (w6561, w6450, IN55[26], w6562, w6563);
  FullAdder U1455 (w6563, w6452, IN56[26], w6564, w6565);
  FullAdder U1456 (w6565, w6454, IN57[26], w6566, w6567);
  FullAdder U1457 (w6567, w6456, IN58[24], w6568, w6569);
  FullAdder U1458 (w6569, w6458, IN59[23], w6570, w6571);
  FullAdder U1459 (w6571, w6460, IN60[22], w6572, w6573);
  FullAdder U1460 (w6573, w6462, IN61[21], w6574, w6575);
  FullAdder U1461 (w6575, w6464, IN62[20], w6576, w6577);
  FullAdder U1462 (w6577, w6466, IN63[19], w6578, w6579);
  FullAdder U1463 (w6579, w6468, IN64[18], w6580, w6581);
  FullAdder U1464 (w6581, w6470, IN65[17], w6582, w6583);
  FullAdder U1465 (w6583, w6472, IN66[16], w6584, w6585);
  FullAdder U1466 (w6585, w6474, IN67[15], w6586, w6587);
  FullAdder U1467 (w6587, w6476, IN68[14], w6588, w6589);
  FullAdder U1468 (w6589, w6478, IN69[13], w6590, w6591);
  FullAdder U1469 (w6591, w6480, IN70[12], w6592, w6593);
  FullAdder U1470 (w6593, w6482, IN71[11], w6594, w6595);
  FullAdder U1471 (w6595, w6484, IN72[10], w6596, w6597);
  FullAdder U1472 (w6597, w6486, IN73[9], w6598, w6599);
  FullAdder U1473 (w6599, w6488, IN74[8], w6600, w6601);
  FullAdder U1474 (w6601, w6490, IN75[7], w6602, w6603);
  FullAdder U1475 (w6603, w6492, IN76[6], w6604, w6605);
  FullAdder U1476 (w6605, w6494, IN77[5], w6606, w6607);
  FullAdder U1477 (w6607, w6496, IN78[4], w6608, w6609);
  FullAdder U1478 (w6609, w6498, IN79[3], w6610, w6611);
  FullAdder U1479 (w6611, w6500, IN80[2], w6612, w6613);
  FullAdder U1480 (w6613, w6502, IN81[1], w6614, w6615);
  FullAdder U1481 (w6615, w6503, IN82[0], w6616, w6617);
  HalfAdder U1482 (w6506, IN27[27], Out1[27], w6619);
  FullAdder U1483 (w6619, w6508, IN28[27], w6620, w6621);
  FullAdder U1484 (w6621, w6510, IN29[27], w6622, w6623);
  FullAdder U1485 (w6623, w6512, IN30[27], w6624, w6625);
  FullAdder U1486 (w6625, w6514, IN31[27], w6626, w6627);
  FullAdder U1487 (w6627, w6516, IN32[27], w6628, w6629);
  FullAdder U1488 (w6629, w6518, IN33[27], w6630, w6631);
  FullAdder U1489 (w6631, w6520, IN34[27], w6632, w6633);
  FullAdder U1490 (w6633, w6522, IN35[27], w6634, w6635);
  FullAdder U1491 (w6635, w6524, IN36[27], w6636, w6637);
  FullAdder U1492 (w6637, w6526, IN37[27], w6638, w6639);
  FullAdder U1493 (w6639, w6528, IN38[27], w6640, w6641);
  FullAdder U1494 (w6641, w6530, IN39[27], w6642, w6643);
  FullAdder U1495 (w6643, w6532, IN40[27], w6644, w6645);
  FullAdder U1496 (w6645, w6534, IN41[27], w6646, w6647);
  FullAdder U1497 (w6647, w6536, IN42[27], w6648, w6649);
  FullAdder U1498 (w6649, w6538, IN43[27], w6650, w6651);
  FullAdder U1499 (w6651, w6540, IN44[27], w6652, w6653);
  FullAdder U1500 (w6653, w6542, IN45[27], w6654, w6655);
  FullAdder U1501 (w6655, w6544, IN46[27], w6656, w6657);
  FullAdder U1502 (w6657, w6546, IN47[27], w6658, w6659);
  FullAdder U1503 (w6659, w6548, IN48[27], w6660, w6661);
  FullAdder U1504 (w6661, w6550, IN49[27], w6662, w6663);
  FullAdder U1505 (w6663, w6552, IN50[27], w6664, w6665);
  FullAdder U1506 (w6665, w6554, IN51[27], w6666, w6667);
  FullAdder U1507 (w6667, w6556, IN52[27], w6668, w6669);
  FullAdder U1508 (w6669, w6558, IN53[27], w6670, w6671);
  FullAdder U1509 (w6671, w6560, IN54[27], w6672, w6673);
  FullAdder U1510 (w6673, w6562, IN55[27], w6674, w6675);
  FullAdder U1511 (w6675, w6564, IN56[27], w6676, w6677);
  FullAdder U1512 (w6677, w6566, IN57[27], w6678, w6679);
  FullAdder U1513 (w6679, w6568, IN58[25], w6680, w6681);
  FullAdder U1514 (w6681, w6570, IN59[24], w6682, w6683);
  FullAdder U1515 (w6683, w6572, IN60[23], w6684, w6685);
  FullAdder U1516 (w6685, w6574, IN61[22], w6686, w6687);
  FullAdder U1517 (w6687, w6576, IN62[21], w6688, w6689);
  FullAdder U1518 (w6689, w6578, IN63[20], w6690, w6691);
  FullAdder U1519 (w6691, w6580, IN64[19], w6692, w6693);
  FullAdder U1520 (w6693, w6582, IN65[18], w6694, w6695);
  FullAdder U1521 (w6695, w6584, IN66[17], w6696, w6697);
  FullAdder U1522 (w6697, w6586, IN67[16], w6698, w6699);
  FullAdder U1523 (w6699, w6588, IN68[15], w6700, w6701);
  FullAdder U1524 (w6701, w6590, IN69[14], w6702, w6703);
  FullAdder U1525 (w6703, w6592, IN70[13], w6704, w6705);
  FullAdder U1526 (w6705, w6594, IN71[12], w6706, w6707);
  FullAdder U1527 (w6707, w6596, IN72[11], w6708, w6709);
  FullAdder U1528 (w6709, w6598, IN73[10], w6710, w6711);
  FullAdder U1529 (w6711, w6600, IN74[9], w6712, w6713);
  FullAdder U1530 (w6713, w6602, IN75[8], w6714, w6715);
  FullAdder U1531 (w6715, w6604, IN76[7], w6716, w6717);
  FullAdder U1532 (w6717, w6606, IN77[6], w6718, w6719);
  FullAdder U1533 (w6719, w6608, IN78[5], w6720, w6721);
  FullAdder U1534 (w6721, w6610, IN79[4], w6722, w6723);
  FullAdder U1535 (w6723, w6612, IN80[3], w6724, w6725);
  FullAdder U1536 (w6725, w6614, IN81[2], w6726, w6727);
  FullAdder U1537 (w6727, w6616, IN82[1], w6728, w6729);
  FullAdder U1538 (w6729, w6617, IN83[0], w6730, w6731);
  HalfAdder U1539 (w6620, IN28[28], Out1[28], w6733);
  FullAdder U1540 (w6733, w6622, IN29[28], w6734, w6735);
  FullAdder U1541 (w6735, w6624, IN30[28], w6736, w6737);
  FullAdder U1542 (w6737, w6626, IN31[28], w6738, w6739);
  FullAdder U1543 (w6739, w6628, IN32[28], w6740, w6741);
  FullAdder U1544 (w6741, w6630, IN33[28], w6742, w6743);
  FullAdder U1545 (w6743, w6632, IN34[28], w6744, w6745);
  FullAdder U1546 (w6745, w6634, IN35[28], w6746, w6747);
  FullAdder U1547 (w6747, w6636, IN36[28], w6748, w6749);
  FullAdder U1548 (w6749, w6638, IN37[28], w6750, w6751);
  FullAdder U1549 (w6751, w6640, IN38[28], w6752, w6753);
  FullAdder U1550 (w6753, w6642, IN39[28], w6754, w6755);
  FullAdder U1551 (w6755, w6644, IN40[28], w6756, w6757);
  FullAdder U1552 (w6757, w6646, IN41[28], w6758, w6759);
  FullAdder U1553 (w6759, w6648, IN42[28], w6760, w6761);
  FullAdder U1554 (w6761, w6650, IN43[28], w6762, w6763);
  FullAdder U1555 (w6763, w6652, IN44[28], w6764, w6765);
  FullAdder U1556 (w6765, w6654, IN45[28], w6766, w6767);
  FullAdder U1557 (w6767, w6656, IN46[28], w6768, w6769);
  FullAdder U1558 (w6769, w6658, IN47[28], w6770, w6771);
  FullAdder U1559 (w6771, w6660, IN48[28], w6772, w6773);
  FullAdder U1560 (w6773, w6662, IN49[28], w6774, w6775);
  FullAdder U1561 (w6775, w6664, IN50[28], w6776, w6777);
  FullAdder U1562 (w6777, w6666, IN51[28], w6778, w6779);
  FullAdder U1563 (w6779, w6668, IN52[28], w6780, w6781);
  FullAdder U1564 (w6781, w6670, IN53[28], w6782, w6783);
  FullAdder U1565 (w6783, w6672, IN54[28], w6784, w6785);
  FullAdder U1566 (w6785, w6674, IN55[28], w6786, w6787);
  FullAdder U1567 (w6787, w6676, IN56[28], w6788, w6789);
  FullAdder U1568 (w6789, w6678, IN57[28], w6790, w6791);
  FullAdder U1569 (w6791, w6680, IN58[26], w6792, w6793);
  FullAdder U1570 (w6793, w6682, IN59[25], w6794, w6795);
  FullAdder U1571 (w6795, w6684, IN60[24], w6796, w6797);
  FullAdder U1572 (w6797, w6686, IN61[23], w6798, w6799);
  FullAdder U1573 (w6799, w6688, IN62[22], w6800, w6801);
  FullAdder U1574 (w6801, w6690, IN63[21], w6802, w6803);
  FullAdder U1575 (w6803, w6692, IN64[20], w6804, w6805);
  FullAdder U1576 (w6805, w6694, IN65[19], w6806, w6807);
  FullAdder U1577 (w6807, w6696, IN66[18], w6808, w6809);
  FullAdder U1578 (w6809, w6698, IN67[17], w6810, w6811);
  FullAdder U1579 (w6811, w6700, IN68[16], w6812, w6813);
  FullAdder U1580 (w6813, w6702, IN69[15], w6814, w6815);
  FullAdder U1581 (w6815, w6704, IN70[14], w6816, w6817);
  FullAdder U1582 (w6817, w6706, IN71[13], w6818, w6819);
  FullAdder U1583 (w6819, w6708, IN72[12], w6820, w6821);
  FullAdder U1584 (w6821, w6710, IN73[11], w6822, w6823);
  FullAdder U1585 (w6823, w6712, IN74[10], w6824, w6825);
  FullAdder U1586 (w6825, w6714, IN75[9], w6826, w6827);
  FullAdder U1587 (w6827, w6716, IN76[8], w6828, w6829);
  FullAdder U1588 (w6829, w6718, IN77[7], w6830, w6831);
  FullAdder U1589 (w6831, w6720, IN78[6], w6832, w6833);
  FullAdder U1590 (w6833, w6722, IN79[5], w6834, w6835);
  FullAdder U1591 (w6835, w6724, IN80[4], w6836, w6837);
  FullAdder U1592 (w6837, w6726, IN81[3], w6838, w6839);
  FullAdder U1593 (w6839, w6728, IN82[2], w6840, w6841);
  FullAdder U1594 (w6841, w6730, IN83[1], w6842, w6843);
  FullAdder U1595 (w6843, w6731, IN84[0], w6844, w6845);
  HalfAdder U1596 (w6734, IN29[29], Out1[29], w6847);
  FullAdder U1597 (w6847, w6736, IN30[29], w6848, w6849);
  FullAdder U1598 (w6849, w6738, IN31[29], w6850, w6851);
  FullAdder U1599 (w6851, w6740, IN32[29], w6852, w6853);
  FullAdder U1600 (w6853, w6742, IN33[29], w6854, w6855);
  FullAdder U1601 (w6855, w6744, IN34[29], w6856, w6857);
  FullAdder U1602 (w6857, w6746, IN35[29], w6858, w6859);
  FullAdder U1603 (w6859, w6748, IN36[29], w6860, w6861);
  FullAdder U1604 (w6861, w6750, IN37[29], w6862, w6863);
  FullAdder U1605 (w6863, w6752, IN38[29], w6864, w6865);
  FullAdder U1606 (w6865, w6754, IN39[29], w6866, w6867);
  FullAdder U1607 (w6867, w6756, IN40[29], w6868, w6869);
  FullAdder U1608 (w6869, w6758, IN41[29], w6870, w6871);
  FullAdder U1609 (w6871, w6760, IN42[29], w6872, w6873);
  FullAdder U1610 (w6873, w6762, IN43[29], w6874, w6875);
  FullAdder U1611 (w6875, w6764, IN44[29], w6876, w6877);
  FullAdder U1612 (w6877, w6766, IN45[29], w6878, w6879);
  FullAdder U1613 (w6879, w6768, IN46[29], w6880, w6881);
  FullAdder U1614 (w6881, w6770, IN47[29], w6882, w6883);
  FullAdder U1615 (w6883, w6772, IN48[29], w6884, w6885);
  FullAdder U1616 (w6885, w6774, IN49[29], w6886, w6887);
  FullAdder U1617 (w6887, w6776, IN50[29], w6888, w6889);
  FullAdder U1618 (w6889, w6778, IN51[29], w6890, w6891);
  FullAdder U1619 (w6891, w6780, IN52[29], w6892, w6893);
  FullAdder U1620 (w6893, w6782, IN53[29], w6894, w6895);
  FullAdder U1621 (w6895, w6784, IN54[29], w6896, w6897);
  FullAdder U1622 (w6897, w6786, IN55[29], w6898, w6899);
  FullAdder U1623 (w6899, w6788, IN56[29], w6900, w6901);
  FullAdder U1624 (w6901, w6790, IN57[29], w6902, w6903);
  FullAdder U1625 (w6903, w6792, IN58[27], w6904, w6905);
  FullAdder U1626 (w6905, w6794, IN59[26], w6906, w6907);
  FullAdder U1627 (w6907, w6796, IN60[25], w6908, w6909);
  FullAdder U1628 (w6909, w6798, IN61[24], w6910, w6911);
  FullAdder U1629 (w6911, w6800, IN62[23], w6912, w6913);
  FullAdder U1630 (w6913, w6802, IN63[22], w6914, w6915);
  FullAdder U1631 (w6915, w6804, IN64[21], w6916, w6917);
  FullAdder U1632 (w6917, w6806, IN65[20], w6918, w6919);
  FullAdder U1633 (w6919, w6808, IN66[19], w6920, w6921);
  FullAdder U1634 (w6921, w6810, IN67[18], w6922, w6923);
  FullAdder U1635 (w6923, w6812, IN68[17], w6924, w6925);
  FullAdder U1636 (w6925, w6814, IN69[16], w6926, w6927);
  FullAdder U1637 (w6927, w6816, IN70[15], w6928, w6929);
  FullAdder U1638 (w6929, w6818, IN71[14], w6930, w6931);
  FullAdder U1639 (w6931, w6820, IN72[13], w6932, w6933);
  FullAdder U1640 (w6933, w6822, IN73[12], w6934, w6935);
  FullAdder U1641 (w6935, w6824, IN74[11], w6936, w6937);
  FullAdder U1642 (w6937, w6826, IN75[10], w6938, w6939);
  FullAdder U1643 (w6939, w6828, IN76[9], w6940, w6941);
  FullAdder U1644 (w6941, w6830, IN77[8], w6942, w6943);
  FullAdder U1645 (w6943, w6832, IN78[7], w6944, w6945);
  FullAdder U1646 (w6945, w6834, IN79[6], w6946, w6947);
  FullAdder U1647 (w6947, w6836, IN80[5], w6948, w6949);
  FullAdder U1648 (w6949, w6838, IN81[4], w6950, w6951);
  FullAdder U1649 (w6951, w6840, IN82[3], w6952, w6953);
  FullAdder U1650 (w6953, w6842, IN83[2], w6954, w6955);
  FullAdder U1651 (w6955, w6844, IN84[1], w6956, w6957);
  FullAdder U1652 (w6957, w6845, IN85[0], w6958, w6959);
  HalfAdder U1653 (w6848, IN30[30], Out1[30], w6961);
  FullAdder U1654 (w6961, w6850, IN31[30], w6962, w6963);
  FullAdder U1655 (w6963, w6852, IN32[30], w6964, w6965);
  FullAdder U1656 (w6965, w6854, IN33[30], w6966, w6967);
  FullAdder U1657 (w6967, w6856, IN34[30], w6968, w6969);
  FullAdder U1658 (w6969, w6858, IN35[30], w6970, w6971);
  FullAdder U1659 (w6971, w6860, IN36[30], w6972, w6973);
  FullAdder U1660 (w6973, w6862, IN37[30], w6974, w6975);
  FullAdder U1661 (w6975, w6864, IN38[30], w6976, w6977);
  FullAdder U1662 (w6977, w6866, IN39[30], w6978, w6979);
  FullAdder U1663 (w6979, w6868, IN40[30], w6980, w6981);
  FullAdder U1664 (w6981, w6870, IN41[30], w6982, w6983);
  FullAdder U1665 (w6983, w6872, IN42[30], w6984, w6985);
  FullAdder U1666 (w6985, w6874, IN43[30], w6986, w6987);
  FullAdder U1667 (w6987, w6876, IN44[30], w6988, w6989);
  FullAdder U1668 (w6989, w6878, IN45[30], w6990, w6991);
  FullAdder U1669 (w6991, w6880, IN46[30], w6992, w6993);
  FullAdder U1670 (w6993, w6882, IN47[30], w6994, w6995);
  FullAdder U1671 (w6995, w6884, IN48[30], w6996, w6997);
  FullAdder U1672 (w6997, w6886, IN49[30], w6998, w6999);
  FullAdder U1673 (w6999, w6888, IN50[30], w7000, w7001);
  FullAdder U1674 (w7001, w6890, IN51[30], w7002, w7003);
  FullAdder U1675 (w7003, w6892, IN52[30], w7004, w7005);
  FullAdder U1676 (w7005, w6894, IN53[30], w7006, w7007);
  FullAdder U1677 (w7007, w6896, IN54[30], w7008, w7009);
  FullAdder U1678 (w7009, w6898, IN55[30], w7010, w7011);
  FullAdder U1679 (w7011, w6900, IN56[30], w7012, w7013);
  FullAdder U1680 (w7013, w6902, IN57[30], w7014, w7015);
  FullAdder U1681 (w7015, w6904, IN58[28], w7016, w7017);
  FullAdder U1682 (w7017, w6906, IN59[27], w7018, w7019);
  FullAdder U1683 (w7019, w6908, IN60[26], w7020, w7021);
  FullAdder U1684 (w7021, w6910, IN61[25], w7022, w7023);
  FullAdder U1685 (w7023, w6912, IN62[24], w7024, w7025);
  FullAdder U1686 (w7025, w6914, IN63[23], w7026, w7027);
  FullAdder U1687 (w7027, w6916, IN64[22], w7028, w7029);
  FullAdder U1688 (w7029, w6918, IN65[21], w7030, w7031);
  FullAdder U1689 (w7031, w6920, IN66[20], w7032, w7033);
  FullAdder U1690 (w7033, w6922, IN67[19], w7034, w7035);
  FullAdder U1691 (w7035, w6924, IN68[18], w7036, w7037);
  FullAdder U1692 (w7037, w6926, IN69[17], w7038, w7039);
  FullAdder U1693 (w7039, w6928, IN70[16], w7040, w7041);
  FullAdder U1694 (w7041, w6930, IN71[15], w7042, w7043);
  FullAdder U1695 (w7043, w6932, IN72[14], w7044, w7045);
  FullAdder U1696 (w7045, w6934, IN73[13], w7046, w7047);
  FullAdder U1697 (w7047, w6936, IN74[12], w7048, w7049);
  FullAdder U1698 (w7049, w6938, IN75[11], w7050, w7051);
  FullAdder U1699 (w7051, w6940, IN76[10], w7052, w7053);
  FullAdder U1700 (w7053, w6942, IN77[9], w7054, w7055);
  FullAdder U1701 (w7055, w6944, IN78[8], w7056, w7057);
  FullAdder U1702 (w7057, w6946, IN79[7], w7058, w7059);
  FullAdder U1703 (w7059, w6948, IN80[6], w7060, w7061);
  FullAdder U1704 (w7061, w6950, IN81[5], w7062, w7063);
  FullAdder U1705 (w7063, w6952, IN82[4], w7064, w7065);
  FullAdder U1706 (w7065, w6954, IN83[3], w7066, w7067);
  FullAdder U1707 (w7067, w6956, IN84[2], w7068, w7069);
  FullAdder U1708 (w7069, w6958, IN85[1], w7070, w7071);
  FullAdder U1709 (w7071, w6959, IN86[0], w7072, w7073);
  HalfAdder U1710 (w6962, IN31[31], Out1[31], w7075);
  FullAdder U1711 (w7075, w6964, IN32[31], w7076, w7077);
  FullAdder U1712 (w7077, w6966, IN33[31], w7078, w7079);
  FullAdder U1713 (w7079, w6968, IN34[31], w7080, w7081);
  FullAdder U1714 (w7081, w6970, IN35[31], w7082, w7083);
  FullAdder U1715 (w7083, w6972, IN36[31], w7084, w7085);
  FullAdder U1716 (w7085, w6974, IN37[31], w7086, w7087);
  FullAdder U1717 (w7087, w6976, IN38[31], w7088, w7089);
  FullAdder U1718 (w7089, w6978, IN39[31], w7090, w7091);
  FullAdder U1719 (w7091, w6980, IN40[31], w7092, w7093);
  FullAdder U1720 (w7093, w6982, IN41[31], w7094, w7095);
  FullAdder U1721 (w7095, w6984, IN42[31], w7096, w7097);
  FullAdder U1722 (w7097, w6986, IN43[31], w7098, w7099);
  FullAdder U1723 (w7099, w6988, IN44[31], w7100, w7101);
  FullAdder U1724 (w7101, w6990, IN45[31], w7102, w7103);
  FullAdder U1725 (w7103, w6992, IN46[31], w7104, w7105);
  FullAdder U1726 (w7105, w6994, IN47[31], w7106, w7107);
  FullAdder U1727 (w7107, w6996, IN48[31], w7108, w7109);
  FullAdder U1728 (w7109, w6998, IN49[31], w7110, w7111);
  FullAdder U1729 (w7111, w7000, IN50[31], w7112, w7113);
  FullAdder U1730 (w7113, w7002, IN51[31], w7114, w7115);
  FullAdder U1731 (w7115, w7004, IN52[31], w7116, w7117);
  FullAdder U1732 (w7117, w7006, IN53[31], w7118, w7119);
  FullAdder U1733 (w7119, w7008, IN54[31], w7120, w7121);
  FullAdder U1734 (w7121, w7010, IN55[31], w7122, w7123);
  FullAdder U1735 (w7123, w7012, IN56[31], w7124, w7125);
  FullAdder U1736 (w7125, w7014, IN57[31], w7126, w7127);
  FullAdder U1737 (w7127, w7016, IN58[29], w7128, w7129);
  FullAdder U1738 (w7129, w7018, IN59[28], w7130, w7131);
  FullAdder U1739 (w7131, w7020, IN60[27], w7132, w7133);
  FullAdder U1740 (w7133, w7022, IN61[26], w7134, w7135);
  FullAdder U1741 (w7135, w7024, IN62[25], w7136, w7137);
  FullAdder U1742 (w7137, w7026, IN63[24], w7138, w7139);
  FullAdder U1743 (w7139, w7028, IN64[23], w7140, w7141);
  FullAdder U1744 (w7141, w7030, IN65[22], w7142, w7143);
  FullAdder U1745 (w7143, w7032, IN66[21], w7144, w7145);
  FullAdder U1746 (w7145, w7034, IN67[20], w7146, w7147);
  FullAdder U1747 (w7147, w7036, IN68[19], w7148, w7149);
  FullAdder U1748 (w7149, w7038, IN69[18], w7150, w7151);
  FullAdder U1749 (w7151, w7040, IN70[17], w7152, w7153);
  FullAdder U1750 (w7153, w7042, IN71[16], w7154, w7155);
  FullAdder U1751 (w7155, w7044, IN72[15], w7156, w7157);
  FullAdder U1752 (w7157, w7046, IN73[14], w7158, w7159);
  FullAdder U1753 (w7159, w7048, IN74[13], w7160, w7161);
  FullAdder U1754 (w7161, w7050, IN75[12], w7162, w7163);
  FullAdder U1755 (w7163, w7052, IN76[11], w7164, w7165);
  FullAdder U1756 (w7165, w7054, IN77[10], w7166, w7167);
  FullAdder U1757 (w7167, w7056, IN78[9], w7168, w7169);
  FullAdder U1758 (w7169, w7058, IN79[8], w7170, w7171);
  FullAdder U1759 (w7171, w7060, IN80[7], w7172, w7173);
  FullAdder U1760 (w7173, w7062, IN81[6], w7174, w7175);
  FullAdder U1761 (w7175, w7064, IN82[5], w7176, w7177);
  FullAdder U1762 (w7177, w7066, IN83[4], w7178, w7179);
  FullAdder U1763 (w7179, w7068, IN84[3], w7180, w7181);
  FullAdder U1764 (w7181, w7070, IN85[2], w7182, w7183);
  FullAdder U1765 (w7183, w7072, IN86[1], w7184, w7185);
  FullAdder U1766 (w7185, w7073, IN87[0], w7186, w7187);
  HalfAdder U1767 (w7076, IN32[32], Out1[32], w7189);
  FullAdder U1768 (w7189, w7078, IN33[32], w7190, w7191);
  FullAdder U1769 (w7191, w7080, IN34[32], w7192, w7193);
  FullAdder U1770 (w7193, w7082, IN35[32], w7194, w7195);
  FullAdder U1771 (w7195, w7084, IN36[32], w7196, w7197);
  FullAdder U1772 (w7197, w7086, IN37[32], w7198, w7199);
  FullAdder U1773 (w7199, w7088, IN38[32], w7200, w7201);
  FullAdder U1774 (w7201, w7090, IN39[32], w7202, w7203);
  FullAdder U1775 (w7203, w7092, IN40[32], w7204, w7205);
  FullAdder U1776 (w7205, w7094, IN41[32], w7206, w7207);
  FullAdder U1777 (w7207, w7096, IN42[32], w7208, w7209);
  FullAdder U1778 (w7209, w7098, IN43[32], w7210, w7211);
  FullAdder U1779 (w7211, w7100, IN44[32], w7212, w7213);
  FullAdder U1780 (w7213, w7102, IN45[32], w7214, w7215);
  FullAdder U1781 (w7215, w7104, IN46[32], w7216, w7217);
  FullAdder U1782 (w7217, w7106, IN47[32], w7218, w7219);
  FullAdder U1783 (w7219, w7108, IN48[32], w7220, w7221);
  FullAdder U1784 (w7221, w7110, IN49[32], w7222, w7223);
  FullAdder U1785 (w7223, w7112, IN50[32], w7224, w7225);
  FullAdder U1786 (w7225, w7114, IN51[32], w7226, w7227);
  FullAdder U1787 (w7227, w7116, IN52[32], w7228, w7229);
  FullAdder U1788 (w7229, w7118, IN53[32], w7230, w7231);
  FullAdder U1789 (w7231, w7120, IN54[32], w7232, w7233);
  FullAdder U1790 (w7233, w7122, IN55[32], w7234, w7235);
  FullAdder U1791 (w7235, w7124, IN56[32], w7236, w7237);
  FullAdder U1792 (w7237, w7126, IN57[32], w7238, w7239);
  FullAdder U1793 (w7239, w7128, IN58[30], w7240, w7241);
  FullAdder U1794 (w7241, w7130, IN59[29], w7242, w7243);
  FullAdder U1795 (w7243, w7132, IN60[28], w7244, w7245);
  FullAdder U1796 (w7245, w7134, IN61[27], w7246, w7247);
  FullAdder U1797 (w7247, w7136, IN62[26], w7248, w7249);
  FullAdder U1798 (w7249, w7138, IN63[25], w7250, w7251);
  FullAdder U1799 (w7251, w7140, IN64[24], w7252, w7253);
  FullAdder U1800 (w7253, w7142, IN65[23], w7254, w7255);
  FullAdder U1801 (w7255, w7144, IN66[22], w7256, w7257);
  FullAdder U1802 (w7257, w7146, IN67[21], w7258, w7259);
  FullAdder U1803 (w7259, w7148, IN68[20], w7260, w7261);
  FullAdder U1804 (w7261, w7150, IN69[19], w7262, w7263);
  FullAdder U1805 (w7263, w7152, IN70[18], w7264, w7265);
  FullAdder U1806 (w7265, w7154, IN71[17], w7266, w7267);
  FullAdder U1807 (w7267, w7156, IN72[16], w7268, w7269);
  FullAdder U1808 (w7269, w7158, IN73[15], w7270, w7271);
  FullAdder U1809 (w7271, w7160, IN74[14], w7272, w7273);
  FullAdder U1810 (w7273, w7162, IN75[13], w7274, w7275);
  FullAdder U1811 (w7275, w7164, IN76[12], w7276, w7277);
  FullAdder U1812 (w7277, w7166, IN77[11], w7278, w7279);
  FullAdder U1813 (w7279, w7168, IN78[10], w7280, w7281);
  FullAdder U1814 (w7281, w7170, IN79[9], w7282, w7283);
  FullAdder U1815 (w7283, w7172, IN80[8], w7284, w7285);
  FullAdder U1816 (w7285, w7174, IN81[7], w7286, w7287);
  FullAdder U1817 (w7287, w7176, IN82[6], w7288, w7289);
  FullAdder U1818 (w7289, w7178, IN83[5], w7290, w7291);
  FullAdder U1819 (w7291, w7180, IN84[4], w7292, w7293);
  FullAdder U1820 (w7293, w7182, IN85[3], w7294, w7295);
  FullAdder U1821 (w7295, w7184, IN86[2], w7296, w7297);
  FullAdder U1822 (w7297, w7186, IN87[1], w7298, w7299);
  FullAdder U1823 (w7299, w7187, IN88[0], w7300, w7301);
  HalfAdder U1824 (w7190, IN33[33], Out1[33], w7303);
  FullAdder U1825 (w7303, w7192, IN34[33], w7304, w7305);
  FullAdder U1826 (w7305, w7194, IN35[33], w7306, w7307);
  FullAdder U1827 (w7307, w7196, IN36[33], w7308, w7309);
  FullAdder U1828 (w7309, w7198, IN37[33], w7310, w7311);
  FullAdder U1829 (w7311, w7200, IN38[33], w7312, w7313);
  FullAdder U1830 (w7313, w7202, IN39[33], w7314, w7315);
  FullAdder U1831 (w7315, w7204, IN40[33], w7316, w7317);
  FullAdder U1832 (w7317, w7206, IN41[33], w7318, w7319);
  FullAdder U1833 (w7319, w7208, IN42[33], w7320, w7321);
  FullAdder U1834 (w7321, w7210, IN43[33], w7322, w7323);
  FullAdder U1835 (w7323, w7212, IN44[33], w7324, w7325);
  FullAdder U1836 (w7325, w7214, IN45[33], w7326, w7327);
  FullAdder U1837 (w7327, w7216, IN46[33], w7328, w7329);
  FullAdder U1838 (w7329, w7218, IN47[33], w7330, w7331);
  FullAdder U1839 (w7331, w7220, IN48[33], w7332, w7333);
  FullAdder U1840 (w7333, w7222, IN49[33], w7334, w7335);
  FullAdder U1841 (w7335, w7224, IN50[33], w7336, w7337);
  FullAdder U1842 (w7337, w7226, IN51[33], w7338, w7339);
  FullAdder U1843 (w7339, w7228, IN52[33], w7340, w7341);
  FullAdder U1844 (w7341, w7230, IN53[33], w7342, w7343);
  FullAdder U1845 (w7343, w7232, IN54[33], w7344, w7345);
  FullAdder U1846 (w7345, w7234, IN55[33], w7346, w7347);
  FullAdder U1847 (w7347, w7236, IN56[33], w7348, w7349);
  FullAdder U1848 (w7349, w7238, IN57[33], w7350, w7351);
  FullAdder U1849 (w7351, w7240, IN58[31], w7352, w7353);
  FullAdder U1850 (w7353, w7242, IN59[30], w7354, w7355);
  FullAdder U1851 (w7355, w7244, IN60[29], w7356, w7357);
  FullAdder U1852 (w7357, w7246, IN61[28], w7358, w7359);
  FullAdder U1853 (w7359, w7248, IN62[27], w7360, w7361);
  FullAdder U1854 (w7361, w7250, IN63[26], w7362, w7363);
  FullAdder U1855 (w7363, w7252, IN64[25], w7364, w7365);
  FullAdder U1856 (w7365, w7254, IN65[24], w7366, w7367);
  FullAdder U1857 (w7367, w7256, IN66[23], w7368, w7369);
  FullAdder U1858 (w7369, w7258, IN67[22], w7370, w7371);
  FullAdder U1859 (w7371, w7260, IN68[21], w7372, w7373);
  FullAdder U1860 (w7373, w7262, IN69[20], w7374, w7375);
  FullAdder U1861 (w7375, w7264, IN70[19], w7376, w7377);
  FullAdder U1862 (w7377, w7266, IN71[18], w7378, w7379);
  FullAdder U1863 (w7379, w7268, IN72[17], w7380, w7381);
  FullAdder U1864 (w7381, w7270, IN73[16], w7382, w7383);
  FullAdder U1865 (w7383, w7272, IN74[15], w7384, w7385);
  FullAdder U1866 (w7385, w7274, IN75[14], w7386, w7387);
  FullAdder U1867 (w7387, w7276, IN76[13], w7388, w7389);
  FullAdder U1868 (w7389, w7278, IN77[12], w7390, w7391);
  FullAdder U1869 (w7391, w7280, IN78[11], w7392, w7393);
  FullAdder U1870 (w7393, w7282, IN79[10], w7394, w7395);
  FullAdder U1871 (w7395, w7284, IN80[9], w7396, w7397);
  FullAdder U1872 (w7397, w7286, IN81[8], w7398, w7399);
  FullAdder U1873 (w7399, w7288, IN82[7], w7400, w7401);
  FullAdder U1874 (w7401, w7290, IN83[6], w7402, w7403);
  FullAdder U1875 (w7403, w7292, IN84[5], w7404, w7405);
  FullAdder U1876 (w7405, w7294, IN85[4], w7406, w7407);
  FullAdder U1877 (w7407, w7296, IN86[3], w7408, w7409);
  FullAdder U1878 (w7409, w7298, IN87[2], w7410, w7411);
  FullAdder U1879 (w7411, w7300, IN88[1], w7412, w7413);
  FullAdder U1880 (w7413, w7301, IN89[0], w7414, w7415);
  HalfAdder U1881 (w7304, IN34[34], Out1[34], w7417);
  FullAdder U1882 (w7417, w7306, IN35[34], w7418, w7419);
  FullAdder U1883 (w7419, w7308, IN36[34], w7420, w7421);
  FullAdder U1884 (w7421, w7310, IN37[34], w7422, w7423);
  FullAdder U1885 (w7423, w7312, IN38[34], w7424, w7425);
  FullAdder U1886 (w7425, w7314, IN39[34], w7426, w7427);
  FullAdder U1887 (w7427, w7316, IN40[34], w7428, w7429);
  FullAdder U1888 (w7429, w7318, IN41[34], w7430, w7431);
  FullAdder U1889 (w7431, w7320, IN42[34], w7432, w7433);
  FullAdder U1890 (w7433, w7322, IN43[34], w7434, w7435);
  FullAdder U1891 (w7435, w7324, IN44[34], w7436, w7437);
  FullAdder U1892 (w7437, w7326, IN45[34], w7438, w7439);
  FullAdder U1893 (w7439, w7328, IN46[34], w7440, w7441);
  FullAdder U1894 (w7441, w7330, IN47[34], w7442, w7443);
  FullAdder U1895 (w7443, w7332, IN48[34], w7444, w7445);
  FullAdder U1896 (w7445, w7334, IN49[34], w7446, w7447);
  FullAdder U1897 (w7447, w7336, IN50[34], w7448, w7449);
  FullAdder U1898 (w7449, w7338, IN51[34], w7450, w7451);
  FullAdder U1899 (w7451, w7340, IN52[34], w7452, w7453);
  FullAdder U1900 (w7453, w7342, IN53[34], w7454, w7455);
  FullAdder U1901 (w7455, w7344, IN54[34], w7456, w7457);
  FullAdder U1902 (w7457, w7346, IN55[34], w7458, w7459);
  FullAdder U1903 (w7459, w7348, IN56[34], w7460, w7461);
  FullAdder U1904 (w7461, w7350, IN57[34], w7462, w7463);
  FullAdder U1905 (w7463, w7352, IN58[32], w7464, w7465);
  FullAdder U1906 (w7465, w7354, IN59[31], w7466, w7467);
  FullAdder U1907 (w7467, w7356, IN60[30], w7468, w7469);
  FullAdder U1908 (w7469, w7358, IN61[29], w7470, w7471);
  FullAdder U1909 (w7471, w7360, IN62[28], w7472, w7473);
  FullAdder U1910 (w7473, w7362, IN63[27], w7474, w7475);
  FullAdder U1911 (w7475, w7364, IN64[26], w7476, w7477);
  FullAdder U1912 (w7477, w7366, IN65[25], w7478, w7479);
  FullAdder U1913 (w7479, w7368, IN66[24], w7480, w7481);
  FullAdder U1914 (w7481, w7370, IN67[23], w7482, w7483);
  FullAdder U1915 (w7483, w7372, IN68[22], w7484, w7485);
  FullAdder U1916 (w7485, w7374, IN69[21], w7486, w7487);
  FullAdder U1917 (w7487, w7376, IN70[20], w7488, w7489);
  FullAdder U1918 (w7489, w7378, IN71[19], w7490, w7491);
  FullAdder U1919 (w7491, w7380, IN72[18], w7492, w7493);
  FullAdder U1920 (w7493, w7382, IN73[17], w7494, w7495);
  FullAdder U1921 (w7495, w7384, IN74[16], w7496, w7497);
  FullAdder U1922 (w7497, w7386, IN75[15], w7498, w7499);
  FullAdder U1923 (w7499, w7388, IN76[14], w7500, w7501);
  FullAdder U1924 (w7501, w7390, IN77[13], w7502, w7503);
  FullAdder U1925 (w7503, w7392, IN78[12], w7504, w7505);
  FullAdder U1926 (w7505, w7394, IN79[11], w7506, w7507);
  FullAdder U1927 (w7507, w7396, IN80[10], w7508, w7509);
  FullAdder U1928 (w7509, w7398, IN81[9], w7510, w7511);
  FullAdder U1929 (w7511, w7400, IN82[8], w7512, w7513);
  FullAdder U1930 (w7513, w7402, IN83[7], w7514, w7515);
  FullAdder U1931 (w7515, w7404, IN84[6], w7516, w7517);
  FullAdder U1932 (w7517, w7406, IN85[5], w7518, w7519);
  FullAdder U1933 (w7519, w7408, IN86[4], w7520, w7521);
  FullAdder U1934 (w7521, w7410, IN87[3], w7522, w7523);
  FullAdder U1935 (w7523, w7412, IN88[2], w7524, w7525);
  FullAdder U1936 (w7525, w7414, IN89[1], w7526, w7527);
  FullAdder U1937 (w7527, w7415, IN90[0], w7528, w7529);
  HalfAdder U1938 (w7418, IN35[35], Out1[35], w7531);
  FullAdder U1939 (w7531, w7420, IN36[35], w7532, w7533);
  FullAdder U1940 (w7533, w7422, IN37[35], w7534, w7535);
  FullAdder U1941 (w7535, w7424, IN38[35], w7536, w7537);
  FullAdder U1942 (w7537, w7426, IN39[35], w7538, w7539);
  FullAdder U1943 (w7539, w7428, IN40[35], w7540, w7541);
  FullAdder U1944 (w7541, w7430, IN41[35], w7542, w7543);
  FullAdder U1945 (w7543, w7432, IN42[35], w7544, w7545);
  FullAdder U1946 (w7545, w7434, IN43[35], w7546, w7547);
  FullAdder U1947 (w7547, w7436, IN44[35], w7548, w7549);
  FullAdder U1948 (w7549, w7438, IN45[35], w7550, w7551);
  FullAdder U1949 (w7551, w7440, IN46[35], w7552, w7553);
  FullAdder U1950 (w7553, w7442, IN47[35], w7554, w7555);
  FullAdder U1951 (w7555, w7444, IN48[35], w7556, w7557);
  FullAdder U1952 (w7557, w7446, IN49[35], w7558, w7559);
  FullAdder U1953 (w7559, w7448, IN50[35], w7560, w7561);
  FullAdder U1954 (w7561, w7450, IN51[35], w7562, w7563);
  FullAdder U1955 (w7563, w7452, IN52[35], w7564, w7565);
  FullAdder U1956 (w7565, w7454, IN53[35], w7566, w7567);
  FullAdder U1957 (w7567, w7456, IN54[35], w7568, w7569);
  FullAdder U1958 (w7569, w7458, IN55[35], w7570, w7571);
  FullAdder U1959 (w7571, w7460, IN56[35], w7572, w7573);
  FullAdder U1960 (w7573, w7462, IN57[35], w7574, w7575);
  FullAdder U1961 (w7575, w7464, IN58[33], w7576, w7577);
  FullAdder U1962 (w7577, w7466, IN59[32], w7578, w7579);
  FullAdder U1963 (w7579, w7468, IN60[31], w7580, w7581);
  FullAdder U1964 (w7581, w7470, IN61[30], w7582, w7583);
  FullAdder U1965 (w7583, w7472, IN62[29], w7584, w7585);
  FullAdder U1966 (w7585, w7474, IN63[28], w7586, w7587);
  FullAdder U1967 (w7587, w7476, IN64[27], w7588, w7589);
  FullAdder U1968 (w7589, w7478, IN65[26], w7590, w7591);
  FullAdder U1969 (w7591, w7480, IN66[25], w7592, w7593);
  FullAdder U1970 (w7593, w7482, IN67[24], w7594, w7595);
  FullAdder U1971 (w7595, w7484, IN68[23], w7596, w7597);
  FullAdder U1972 (w7597, w7486, IN69[22], w7598, w7599);
  FullAdder U1973 (w7599, w7488, IN70[21], w7600, w7601);
  FullAdder U1974 (w7601, w7490, IN71[20], w7602, w7603);
  FullAdder U1975 (w7603, w7492, IN72[19], w7604, w7605);
  FullAdder U1976 (w7605, w7494, IN73[18], w7606, w7607);
  FullAdder U1977 (w7607, w7496, IN74[17], w7608, w7609);
  FullAdder U1978 (w7609, w7498, IN75[16], w7610, w7611);
  FullAdder U1979 (w7611, w7500, IN76[15], w7612, w7613);
  FullAdder U1980 (w7613, w7502, IN77[14], w7614, w7615);
  FullAdder U1981 (w7615, w7504, IN78[13], w7616, w7617);
  FullAdder U1982 (w7617, w7506, IN79[12], w7618, w7619);
  FullAdder U1983 (w7619, w7508, IN80[11], w7620, w7621);
  FullAdder U1984 (w7621, w7510, IN81[10], w7622, w7623);
  FullAdder U1985 (w7623, w7512, IN82[9], w7624, w7625);
  FullAdder U1986 (w7625, w7514, IN83[8], w7626, w7627);
  FullAdder U1987 (w7627, w7516, IN84[7], w7628, w7629);
  FullAdder U1988 (w7629, w7518, IN85[6], w7630, w7631);
  FullAdder U1989 (w7631, w7520, IN86[5], w7632, w7633);
  FullAdder U1990 (w7633, w7522, IN87[4], w7634, w7635);
  FullAdder U1991 (w7635, w7524, IN88[3], w7636, w7637);
  FullAdder U1992 (w7637, w7526, IN89[2], w7638, w7639);
  FullAdder U1993 (w7639, w7528, IN90[1], w7640, w7641);
  FullAdder U1994 (w7641, w7529, IN91[0], w7642, w7643);
  HalfAdder U1995 (w7532, IN36[36], Out1[36], w7645);
  FullAdder U1996 (w7645, w7534, IN37[36], w7646, w7647);
  FullAdder U1997 (w7647, w7536, IN38[36], w7648, w7649);
  FullAdder U1998 (w7649, w7538, IN39[36], w7650, w7651);
  FullAdder U1999 (w7651, w7540, IN40[36], w7652, w7653);
  FullAdder U2000 (w7653, w7542, IN41[36], w7654, w7655);
  FullAdder U2001 (w7655, w7544, IN42[36], w7656, w7657);
  FullAdder U2002 (w7657, w7546, IN43[36], w7658, w7659);
  FullAdder U2003 (w7659, w7548, IN44[36], w7660, w7661);
  FullAdder U2004 (w7661, w7550, IN45[36], w7662, w7663);
  FullAdder U2005 (w7663, w7552, IN46[36], w7664, w7665);
  FullAdder U2006 (w7665, w7554, IN47[36], w7666, w7667);
  FullAdder U2007 (w7667, w7556, IN48[36], w7668, w7669);
  FullAdder U2008 (w7669, w7558, IN49[36], w7670, w7671);
  FullAdder U2009 (w7671, w7560, IN50[36], w7672, w7673);
  FullAdder U2010 (w7673, w7562, IN51[36], w7674, w7675);
  FullAdder U2011 (w7675, w7564, IN52[36], w7676, w7677);
  FullAdder U2012 (w7677, w7566, IN53[36], w7678, w7679);
  FullAdder U2013 (w7679, w7568, IN54[36], w7680, w7681);
  FullAdder U2014 (w7681, w7570, IN55[36], w7682, w7683);
  FullAdder U2015 (w7683, w7572, IN56[36], w7684, w7685);
  FullAdder U2016 (w7685, w7574, IN57[36], w7686, w7687);
  FullAdder U2017 (w7687, w7576, IN58[34], w7688, w7689);
  FullAdder U2018 (w7689, w7578, IN59[33], w7690, w7691);
  FullAdder U2019 (w7691, w7580, IN60[32], w7692, w7693);
  FullAdder U2020 (w7693, w7582, IN61[31], w7694, w7695);
  FullAdder U2021 (w7695, w7584, IN62[30], w7696, w7697);
  FullAdder U2022 (w7697, w7586, IN63[29], w7698, w7699);
  FullAdder U2023 (w7699, w7588, IN64[28], w7700, w7701);
  FullAdder U2024 (w7701, w7590, IN65[27], w7702, w7703);
  FullAdder U2025 (w7703, w7592, IN66[26], w7704, w7705);
  FullAdder U2026 (w7705, w7594, IN67[25], w7706, w7707);
  FullAdder U2027 (w7707, w7596, IN68[24], w7708, w7709);
  FullAdder U2028 (w7709, w7598, IN69[23], w7710, w7711);
  FullAdder U2029 (w7711, w7600, IN70[22], w7712, w7713);
  FullAdder U2030 (w7713, w7602, IN71[21], w7714, w7715);
  FullAdder U2031 (w7715, w7604, IN72[20], w7716, w7717);
  FullAdder U2032 (w7717, w7606, IN73[19], w7718, w7719);
  FullAdder U2033 (w7719, w7608, IN74[18], w7720, w7721);
  FullAdder U2034 (w7721, w7610, IN75[17], w7722, w7723);
  FullAdder U2035 (w7723, w7612, IN76[16], w7724, w7725);
  FullAdder U2036 (w7725, w7614, IN77[15], w7726, w7727);
  FullAdder U2037 (w7727, w7616, IN78[14], w7728, w7729);
  FullAdder U2038 (w7729, w7618, IN79[13], w7730, w7731);
  FullAdder U2039 (w7731, w7620, IN80[12], w7732, w7733);
  FullAdder U2040 (w7733, w7622, IN81[11], w7734, w7735);
  FullAdder U2041 (w7735, w7624, IN82[10], w7736, w7737);
  FullAdder U2042 (w7737, w7626, IN83[9], w7738, w7739);
  FullAdder U2043 (w7739, w7628, IN84[8], w7740, w7741);
  FullAdder U2044 (w7741, w7630, IN85[7], w7742, w7743);
  FullAdder U2045 (w7743, w7632, IN86[6], w7744, w7745);
  FullAdder U2046 (w7745, w7634, IN87[5], w7746, w7747);
  FullAdder U2047 (w7747, w7636, IN88[4], w7748, w7749);
  FullAdder U2048 (w7749, w7638, IN89[3], w7750, w7751);
  FullAdder U2049 (w7751, w7640, IN90[2], w7752, w7753);
  FullAdder U2050 (w7753, w7642, IN91[1], w7754, w7755);
  FullAdder U2051 (w7755, w7643, IN92[0], w7756, w7757);
  HalfAdder U2052 (w7646, IN37[37], Out1[37], w7759);
  FullAdder U2053 (w7759, w7648, IN38[37], w7760, w7761);
  FullAdder U2054 (w7761, w7650, IN39[37], w7762, w7763);
  FullAdder U2055 (w7763, w7652, IN40[37], w7764, w7765);
  FullAdder U2056 (w7765, w7654, IN41[37], w7766, w7767);
  FullAdder U2057 (w7767, w7656, IN42[37], w7768, w7769);
  FullAdder U2058 (w7769, w7658, IN43[37], w7770, w7771);
  FullAdder U2059 (w7771, w7660, IN44[37], w7772, w7773);
  FullAdder U2060 (w7773, w7662, IN45[37], w7774, w7775);
  FullAdder U2061 (w7775, w7664, IN46[37], w7776, w7777);
  FullAdder U2062 (w7777, w7666, IN47[37], w7778, w7779);
  FullAdder U2063 (w7779, w7668, IN48[37], w7780, w7781);
  FullAdder U2064 (w7781, w7670, IN49[37], w7782, w7783);
  FullAdder U2065 (w7783, w7672, IN50[37], w7784, w7785);
  FullAdder U2066 (w7785, w7674, IN51[37], w7786, w7787);
  FullAdder U2067 (w7787, w7676, IN52[37], w7788, w7789);
  FullAdder U2068 (w7789, w7678, IN53[37], w7790, w7791);
  FullAdder U2069 (w7791, w7680, IN54[37], w7792, w7793);
  FullAdder U2070 (w7793, w7682, IN55[37], w7794, w7795);
  FullAdder U2071 (w7795, w7684, IN56[37], w7796, w7797);
  FullAdder U2072 (w7797, w7686, IN57[37], w7798, w7799);
  FullAdder U2073 (w7799, w7688, IN58[35], w7800, w7801);
  FullAdder U2074 (w7801, w7690, IN59[34], w7802, w7803);
  FullAdder U2075 (w7803, w7692, IN60[33], w7804, w7805);
  FullAdder U2076 (w7805, w7694, IN61[32], w7806, w7807);
  FullAdder U2077 (w7807, w7696, IN62[31], w7808, w7809);
  FullAdder U2078 (w7809, w7698, IN63[30], w7810, w7811);
  FullAdder U2079 (w7811, w7700, IN64[29], w7812, w7813);
  FullAdder U2080 (w7813, w7702, IN65[28], w7814, w7815);
  FullAdder U2081 (w7815, w7704, IN66[27], w7816, w7817);
  FullAdder U2082 (w7817, w7706, IN67[26], w7818, w7819);
  FullAdder U2083 (w7819, w7708, IN68[25], w7820, w7821);
  FullAdder U2084 (w7821, w7710, IN69[24], w7822, w7823);
  FullAdder U2085 (w7823, w7712, IN70[23], w7824, w7825);
  FullAdder U2086 (w7825, w7714, IN71[22], w7826, w7827);
  FullAdder U2087 (w7827, w7716, IN72[21], w7828, w7829);
  FullAdder U2088 (w7829, w7718, IN73[20], w7830, w7831);
  FullAdder U2089 (w7831, w7720, IN74[19], w7832, w7833);
  FullAdder U2090 (w7833, w7722, IN75[18], w7834, w7835);
  FullAdder U2091 (w7835, w7724, IN76[17], w7836, w7837);
  FullAdder U2092 (w7837, w7726, IN77[16], w7838, w7839);
  FullAdder U2093 (w7839, w7728, IN78[15], w7840, w7841);
  FullAdder U2094 (w7841, w7730, IN79[14], w7842, w7843);
  FullAdder U2095 (w7843, w7732, IN80[13], w7844, w7845);
  FullAdder U2096 (w7845, w7734, IN81[12], w7846, w7847);
  FullAdder U2097 (w7847, w7736, IN82[11], w7848, w7849);
  FullAdder U2098 (w7849, w7738, IN83[10], w7850, w7851);
  FullAdder U2099 (w7851, w7740, IN84[9], w7852, w7853);
  FullAdder U2100 (w7853, w7742, IN85[8], w7854, w7855);
  FullAdder U2101 (w7855, w7744, IN86[7], w7856, w7857);
  FullAdder U2102 (w7857, w7746, IN87[6], w7858, w7859);
  FullAdder U2103 (w7859, w7748, IN88[5], w7860, w7861);
  FullAdder U2104 (w7861, w7750, IN89[4], w7862, w7863);
  FullAdder U2105 (w7863, w7752, IN90[3], w7864, w7865);
  FullAdder U2106 (w7865, w7754, IN91[2], w7866, w7867);
  FullAdder U2107 (w7867, w7756, IN92[1], w7868, w7869);
  FullAdder U2108 (w7869, w7757, IN93[0], w7870, w7871);
  HalfAdder U2109 (w7760, IN38[38], Out1[38], w7873);
  FullAdder U2110 (w7873, w7762, IN39[38], w7874, w7875);
  FullAdder U2111 (w7875, w7764, IN40[38], w7876, w7877);
  FullAdder U2112 (w7877, w7766, IN41[38], w7878, w7879);
  FullAdder U2113 (w7879, w7768, IN42[38], w7880, w7881);
  FullAdder U2114 (w7881, w7770, IN43[38], w7882, w7883);
  FullAdder U2115 (w7883, w7772, IN44[38], w7884, w7885);
  FullAdder U2116 (w7885, w7774, IN45[38], w7886, w7887);
  FullAdder U2117 (w7887, w7776, IN46[38], w7888, w7889);
  FullAdder U2118 (w7889, w7778, IN47[38], w7890, w7891);
  FullAdder U2119 (w7891, w7780, IN48[38], w7892, w7893);
  FullAdder U2120 (w7893, w7782, IN49[38], w7894, w7895);
  FullAdder U2121 (w7895, w7784, IN50[38], w7896, w7897);
  FullAdder U2122 (w7897, w7786, IN51[38], w7898, w7899);
  FullAdder U2123 (w7899, w7788, IN52[38], w7900, w7901);
  FullAdder U2124 (w7901, w7790, IN53[38], w7902, w7903);
  FullAdder U2125 (w7903, w7792, IN54[38], w7904, w7905);
  FullAdder U2126 (w7905, w7794, IN55[38], w7906, w7907);
  FullAdder U2127 (w7907, w7796, IN56[38], w7908, w7909);
  FullAdder U2128 (w7909, w7798, IN57[38], w7910, w7911);
  FullAdder U2129 (w7911, w7800, IN58[36], w7912, w7913);
  FullAdder U2130 (w7913, w7802, IN59[35], w7914, w7915);
  FullAdder U2131 (w7915, w7804, IN60[34], w7916, w7917);
  FullAdder U2132 (w7917, w7806, IN61[33], w7918, w7919);
  FullAdder U2133 (w7919, w7808, IN62[32], w7920, w7921);
  FullAdder U2134 (w7921, w7810, IN63[31], w7922, w7923);
  FullAdder U2135 (w7923, w7812, IN64[30], w7924, w7925);
  FullAdder U2136 (w7925, w7814, IN65[29], w7926, w7927);
  FullAdder U2137 (w7927, w7816, IN66[28], w7928, w7929);
  FullAdder U2138 (w7929, w7818, IN67[27], w7930, w7931);
  FullAdder U2139 (w7931, w7820, IN68[26], w7932, w7933);
  FullAdder U2140 (w7933, w7822, IN69[25], w7934, w7935);
  FullAdder U2141 (w7935, w7824, IN70[24], w7936, w7937);
  FullAdder U2142 (w7937, w7826, IN71[23], w7938, w7939);
  FullAdder U2143 (w7939, w7828, IN72[22], w7940, w7941);
  FullAdder U2144 (w7941, w7830, IN73[21], w7942, w7943);
  FullAdder U2145 (w7943, w7832, IN74[20], w7944, w7945);
  FullAdder U2146 (w7945, w7834, IN75[19], w7946, w7947);
  FullAdder U2147 (w7947, w7836, IN76[18], w7948, w7949);
  FullAdder U2148 (w7949, w7838, IN77[17], w7950, w7951);
  FullAdder U2149 (w7951, w7840, IN78[16], w7952, w7953);
  FullAdder U2150 (w7953, w7842, IN79[15], w7954, w7955);
  FullAdder U2151 (w7955, w7844, IN80[14], w7956, w7957);
  FullAdder U2152 (w7957, w7846, IN81[13], w7958, w7959);
  FullAdder U2153 (w7959, w7848, IN82[12], w7960, w7961);
  FullAdder U2154 (w7961, w7850, IN83[11], w7962, w7963);
  FullAdder U2155 (w7963, w7852, IN84[10], w7964, w7965);
  FullAdder U2156 (w7965, w7854, IN85[9], w7966, w7967);
  FullAdder U2157 (w7967, w7856, IN86[8], w7968, w7969);
  FullAdder U2158 (w7969, w7858, IN87[7], w7970, w7971);
  FullAdder U2159 (w7971, w7860, IN88[6], w7972, w7973);
  FullAdder U2160 (w7973, w7862, IN89[5], w7974, w7975);
  FullAdder U2161 (w7975, w7864, IN90[4], w7976, w7977);
  FullAdder U2162 (w7977, w7866, IN91[3], w7978, w7979);
  FullAdder U2163 (w7979, w7868, IN92[2], w7980, w7981);
  FullAdder U2164 (w7981, w7870, IN93[1], w7982, w7983);
  FullAdder U2165 (w7983, w7871, IN94[0], w7984, w7985);
  HalfAdder U2166 (w7874, IN39[39], Out1[39], w7987);
  FullAdder U2167 (w7987, w7876, IN40[39], w7988, w7989);
  FullAdder U2168 (w7989, w7878, IN41[39], w7990, w7991);
  FullAdder U2169 (w7991, w7880, IN42[39], w7992, w7993);
  FullAdder U2170 (w7993, w7882, IN43[39], w7994, w7995);
  FullAdder U2171 (w7995, w7884, IN44[39], w7996, w7997);
  FullAdder U2172 (w7997, w7886, IN45[39], w7998, w7999);
  FullAdder U2173 (w7999, w7888, IN46[39], w8000, w8001);
  FullAdder U2174 (w8001, w7890, IN47[39], w8002, w8003);
  FullAdder U2175 (w8003, w7892, IN48[39], w8004, w8005);
  FullAdder U2176 (w8005, w7894, IN49[39], w8006, w8007);
  FullAdder U2177 (w8007, w7896, IN50[39], w8008, w8009);
  FullAdder U2178 (w8009, w7898, IN51[39], w8010, w8011);
  FullAdder U2179 (w8011, w7900, IN52[39], w8012, w8013);
  FullAdder U2180 (w8013, w7902, IN53[39], w8014, w8015);
  FullAdder U2181 (w8015, w7904, IN54[39], w8016, w8017);
  FullAdder U2182 (w8017, w7906, IN55[39], w8018, w8019);
  FullAdder U2183 (w8019, w7908, IN56[39], w8020, w8021);
  FullAdder U2184 (w8021, w7910, IN57[39], w8022, w8023);
  FullAdder U2185 (w8023, w7912, IN58[37], w8024, w8025);
  FullAdder U2186 (w8025, w7914, IN59[36], w8026, w8027);
  FullAdder U2187 (w8027, w7916, IN60[35], w8028, w8029);
  FullAdder U2188 (w8029, w7918, IN61[34], w8030, w8031);
  FullAdder U2189 (w8031, w7920, IN62[33], w8032, w8033);
  FullAdder U2190 (w8033, w7922, IN63[32], w8034, w8035);
  FullAdder U2191 (w8035, w7924, IN64[31], w8036, w8037);
  FullAdder U2192 (w8037, w7926, IN65[30], w8038, w8039);
  FullAdder U2193 (w8039, w7928, IN66[29], w8040, w8041);
  FullAdder U2194 (w8041, w7930, IN67[28], w8042, w8043);
  FullAdder U2195 (w8043, w7932, IN68[27], w8044, w8045);
  FullAdder U2196 (w8045, w7934, IN69[26], w8046, w8047);
  FullAdder U2197 (w8047, w7936, IN70[25], w8048, w8049);
  FullAdder U2198 (w8049, w7938, IN71[24], w8050, w8051);
  FullAdder U2199 (w8051, w7940, IN72[23], w8052, w8053);
  FullAdder U2200 (w8053, w7942, IN73[22], w8054, w8055);
  FullAdder U2201 (w8055, w7944, IN74[21], w8056, w8057);
  FullAdder U2202 (w8057, w7946, IN75[20], w8058, w8059);
  FullAdder U2203 (w8059, w7948, IN76[19], w8060, w8061);
  FullAdder U2204 (w8061, w7950, IN77[18], w8062, w8063);
  FullAdder U2205 (w8063, w7952, IN78[17], w8064, w8065);
  FullAdder U2206 (w8065, w7954, IN79[16], w8066, w8067);
  FullAdder U2207 (w8067, w7956, IN80[15], w8068, w8069);
  FullAdder U2208 (w8069, w7958, IN81[14], w8070, w8071);
  FullAdder U2209 (w8071, w7960, IN82[13], w8072, w8073);
  FullAdder U2210 (w8073, w7962, IN83[12], w8074, w8075);
  FullAdder U2211 (w8075, w7964, IN84[11], w8076, w8077);
  FullAdder U2212 (w8077, w7966, IN85[10], w8078, w8079);
  FullAdder U2213 (w8079, w7968, IN86[9], w8080, w8081);
  FullAdder U2214 (w8081, w7970, IN87[8], w8082, w8083);
  FullAdder U2215 (w8083, w7972, IN88[7], w8084, w8085);
  FullAdder U2216 (w8085, w7974, IN89[6], w8086, w8087);
  FullAdder U2217 (w8087, w7976, IN90[5], w8088, w8089);
  FullAdder U2218 (w8089, w7978, IN91[4], w8090, w8091);
  FullAdder U2219 (w8091, w7980, IN92[3], w8092, w8093);
  FullAdder U2220 (w8093, w7982, IN93[2], w8094, w8095);
  FullAdder U2221 (w8095, w7984, IN94[1], w8096, w8097);
  FullAdder U2222 (w8097, w7985, IN95[0], w8098, w8099);
  HalfAdder U2223 (w7988, IN40[40], Out1[40], w8101);
  FullAdder U2224 (w8101, w7990, IN41[40], w8102, w8103);
  FullAdder U2225 (w8103, w7992, IN42[40], w8104, w8105);
  FullAdder U2226 (w8105, w7994, IN43[40], w8106, w8107);
  FullAdder U2227 (w8107, w7996, IN44[40], w8108, w8109);
  FullAdder U2228 (w8109, w7998, IN45[40], w8110, w8111);
  FullAdder U2229 (w8111, w8000, IN46[40], w8112, w8113);
  FullAdder U2230 (w8113, w8002, IN47[40], w8114, w8115);
  FullAdder U2231 (w8115, w8004, IN48[40], w8116, w8117);
  FullAdder U2232 (w8117, w8006, IN49[40], w8118, w8119);
  FullAdder U2233 (w8119, w8008, IN50[40], w8120, w8121);
  FullAdder U2234 (w8121, w8010, IN51[40], w8122, w8123);
  FullAdder U2235 (w8123, w8012, IN52[40], w8124, w8125);
  FullAdder U2236 (w8125, w8014, IN53[40], w8126, w8127);
  FullAdder U2237 (w8127, w8016, IN54[40], w8128, w8129);
  FullAdder U2238 (w8129, w8018, IN55[40], w8130, w8131);
  FullAdder U2239 (w8131, w8020, IN56[40], w8132, w8133);
  FullAdder U2240 (w8133, w8022, IN57[40], w8134, w8135);
  FullAdder U2241 (w8135, w8024, IN58[38], w8136, w8137);
  FullAdder U2242 (w8137, w8026, IN59[37], w8138, w8139);
  FullAdder U2243 (w8139, w8028, IN60[36], w8140, w8141);
  FullAdder U2244 (w8141, w8030, IN61[35], w8142, w8143);
  FullAdder U2245 (w8143, w8032, IN62[34], w8144, w8145);
  FullAdder U2246 (w8145, w8034, IN63[33], w8146, w8147);
  FullAdder U2247 (w8147, w8036, IN64[32], w8148, w8149);
  FullAdder U2248 (w8149, w8038, IN65[31], w8150, w8151);
  FullAdder U2249 (w8151, w8040, IN66[30], w8152, w8153);
  FullAdder U2250 (w8153, w8042, IN67[29], w8154, w8155);
  FullAdder U2251 (w8155, w8044, IN68[28], w8156, w8157);
  FullAdder U2252 (w8157, w8046, IN69[27], w8158, w8159);
  FullAdder U2253 (w8159, w8048, IN70[26], w8160, w8161);
  FullAdder U2254 (w8161, w8050, IN71[25], w8162, w8163);
  FullAdder U2255 (w8163, w8052, IN72[24], w8164, w8165);
  FullAdder U2256 (w8165, w8054, IN73[23], w8166, w8167);
  FullAdder U2257 (w8167, w8056, IN74[22], w8168, w8169);
  FullAdder U2258 (w8169, w8058, IN75[21], w8170, w8171);
  FullAdder U2259 (w8171, w8060, IN76[20], w8172, w8173);
  FullAdder U2260 (w8173, w8062, IN77[19], w8174, w8175);
  FullAdder U2261 (w8175, w8064, IN78[18], w8176, w8177);
  FullAdder U2262 (w8177, w8066, IN79[17], w8178, w8179);
  FullAdder U2263 (w8179, w8068, IN80[16], w8180, w8181);
  FullAdder U2264 (w8181, w8070, IN81[15], w8182, w8183);
  FullAdder U2265 (w8183, w8072, IN82[14], w8184, w8185);
  FullAdder U2266 (w8185, w8074, IN83[13], w8186, w8187);
  FullAdder U2267 (w8187, w8076, IN84[12], w8188, w8189);
  FullAdder U2268 (w8189, w8078, IN85[11], w8190, w8191);
  FullAdder U2269 (w8191, w8080, IN86[10], w8192, w8193);
  FullAdder U2270 (w8193, w8082, IN87[9], w8194, w8195);
  FullAdder U2271 (w8195, w8084, IN88[8], w8196, w8197);
  FullAdder U2272 (w8197, w8086, IN89[7], w8198, w8199);
  FullAdder U2273 (w8199, w8088, IN90[6], w8200, w8201);
  FullAdder U2274 (w8201, w8090, IN91[5], w8202, w8203);
  FullAdder U2275 (w8203, w8092, IN92[4], w8204, w8205);
  FullAdder U2276 (w8205, w8094, IN93[3], w8206, w8207);
  FullAdder U2277 (w8207, w8096, IN94[2], w8208, w8209);
  FullAdder U2278 (w8209, w8098, IN95[1], w8210, w8211);
  FullAdder U2279 (w8211, w8099, IN96[0], w8212, w8213);
  HalfAdder U2280 (w8102, IN41[41], Out1[41], w8215);
  FullAdder U2281 (w8215, w8104, IN42[41], w8216, w8217);
  FullAdder U2282 (w8217, w8106, IN43[41], w8218, w8219);
  FullAdder U2283 (w8219, w8108, IN44[41], w8220, w8221);
  FullAdder U2284 (w8221, w8110, IN45[41], w8222, w8223);
  FullAdder U2285 (w8223, w8112, IN46[41], w8224, w8225);
  FullAdder U2286 (w8225, w8114, IN47[41], w8226, w8227);
  FullAdder U2287 (w8227, w8116, IN48[41], w8228, w8229);
  FullAdder U2288 (w8229, w8118, IN49[41], w8230, w8231);
  FullAdder U2289 (w8231, w8120, IN50[41], w8232, w8233);
  FullAdder U2290 (w8233, w8122, IN51[41], w8234, w8235);
  FullAdder U2291 (w8235, w8124, IN52[41], w8236, w8237);
  FullAdder U2292 (w8237, w8126, IN53[41], w8238, w8239);
  FullAdder U2293 (w8239, w8128, IN54[41], w8240, w8241);
  FullAdder U2294 (w8241, w8130, IN55[41], w8242, w8243);
  FullAdder U2295 (w8243, w8132, IN56[41], w8244, w8245);
  FullAdder U2296 (w8245, w8134, IN57[41], w8246, w8247);
  FullAdder U2297 (w8247, w8136, IN58[39], w8248, w8249);
  FullAdder U2298 (w8249, w8138, IN59[38], w8250, w8251);
  FullAdder U2299 (w8251, w8140, IN60[37], w8252, w8253);
  FullAdder U2300 (w8253, w8142, IN61[36], w8254, w8255);
  FullAdder U2301 (w8255, w8144, IN62[35], w8256, w8257);
  FullAdder U2302 (w8257, w8146, IN63[34], w8258, w8259);
  FullAdder U2303 (w8259, w8148, IN64[33], w8260, w8261);
  FullAdder U2304 (w8261, w8150, IN65[32], w8262, w8263);
  FullAdder U2305 (w8263, w8152, IN66[31], w8264, w8265);
  FullAdder U2306 (w8265, w8154, IN67[30], w8266, w8267);
  FullAdder U2307 (w8267, w8156, IN68[29], w8268, w8269);
  FullAdder U2308 (w8269, w8158, IN69[28], w8270, w8271);
  FullAdder U2309 (w8271, w8160, IN70[27], w8272, w8273);
  FullAdder U2310 (w8273, w8162, IN71[26], w8274, w8275);
  FullAdder U2311 (w8275, w8164, IN72[25], w8276, w8277);
  FullAdder U2312 (w8277, w8166, IN73[24], w8278, w8279);
  FullAdder U2313 (w8279, w8168, IN74[23], w8280, w8281);
  FullAdder U2314 (w8281, w8170, IN75[22], w8282, w8283);
  FullAdder U2315 (w8283, w8172, IN76[21], w8284, w8285);
  FullAdder U2316 (w8285, w8174, IN77[20], w8286, w8287);
  FullAdder U2317 (w8287, w8176, IN78[19], w8288, w8289);
  FullAdder U2318 (w8289, w8178, IN79[18], w8290, w8291);
  FullAdder U2319 (w8291, w8180, IN80[17], w8292, w8293);
  FullAdder U2320 (w8293, w8182, IN81[16], w8294, w8295);
  FullAdder U2321 (w8295, w8184, IN82[15], w8296, w8297);
  FullAdder U2322 (w8297, w8186, IN83[14], w8298, w8299);
  FullAdder U2323 (w8299, w8188, IN84[13], w8300, w8301);
  FullAdder U2324 (w8301, w8190, IN85[12], w8302, w8303);
  FullAdder U2325 (w8303, w8192, IN86[11], w8304, w8305);
  FullAdder U2326 (w8305, w8194, IN87[10], w8306, w8307);
  FullAdder U2327 (w8307, w8196, IN88[9], w8308, w8309);
  FullAdder U2328 (w8309, w8198, IN89[8], w8310, w8311);
  FullAdder U2329 (w8311, w8200, IN90[7], w8312, w8313);
  FullAdder U2330 (w8313, w8202, IN91[6], w8314, w8315);
  FullAdder U2331 (w8315, w8204, IN92[5], w8316, w8317);
  FullAdder U2332 (w8317, w8206, IN93[4], w8318, w8319);
  FullAdder U2333 (w8319, w8208, IN94[3], w8320, w8321);
  FullAdder U2334 (w8321, w8210, IN95[2], w8322, w8323);
  FullAdder U2335 (w8323, w8212, IN96[1], w8324, w8325);
  FullAdder U2336 (w8325, w8213, IN97[0], w8326, w8327);
  HalfAdder U2337 (w8216, IN42[42], Out1[42], w8329);
  FullAdder U2338 (w8329, w8218, IN43[42], w8330, w8331);
  FullAdder U2339 (w8331, w8220, IN44[42], w8332, w8333);
  FullAdder U2340 (w8333, w8222, IN45[42], w8334, w8335);
  FullAdder U2341 (w8335, w8224, IN46[42], w8336, w8337);
  FullAdder U2342 (w8337, w8226, IN47[42], w8338, w8339);
  FullAdder U2343 (w8339, w8228, IN48[42], w8340, w8341);
  FullAdder U2344 (w8341, w8230, IN49[42], w8342, w8343);
  FullAdder U2345 (w8343, w8232, IN50[42], w8344, w8345);
  FullAdder U2346 (w8345, w8234, IN51[42], w8346, w8347);
  FullAdder U2347 (w8347, w8236, IN52[42], w8348, w8349);
  FullAdder U2348 (w8349, w8238, IN53[42], w8350, w8351);
  FullAdder U2349 (w8351, w8240, IN54[42], w8352, w8353);
  FullAdder U2350 (w8353, w8242, IN55[42], w8354, w8355);
  FullAdder U2351 (w8355, w8244, IN56[42], w8356, w8357);
  FullAdder U2352 (w8357, w8246, IN57[42], w8358, w8359);
  FullAdder U2353 (w8359, w8248, IN58[40], w8360, w8361);
  FullAdder U2354 (w8361, w8250, IN59[39], w8362, w8363);
  FullAdder U2355 (w8363, w8252, IN60[38], w8364, w8365);
  FullAdder U2356 (w8365, w8254, IN61[37], w8366, w8367);
  FullAdder U2357 (w8367, w8256, IN62[36], w8368, w8369);
  FullAdder U2358 (w8369, w8258, IN63[35], w8370, w8371);
  FullAdder U2359 (w8371, w8260, IN64[34], w8372, w8373);
  FullAdder U2360 (w8373, w8262, IN65[33], w8374, w8375);
  FullAdder U2361 (w8375, w8264, IN66[32], w8376, w8377);
  FullAdder U2362 (w8377, w8266, IN67[31], w8378, w8379);
  FullAdder U2363 (w8379, w8268, IN68[30], w8380, w8381);
  FullAdder U2364 (w8381, w8270, IN69[29], w8382, w8383);
  FullAdder U2365 (w8383, w8272, IN70[28], w8384, w8385);
  FullAdder U2366 (w8385, w8274, IN71[27], w8386, w8387);
  FullAdder U2367 (w8387, w8276, IN72[26], w8388, w8389);
  FullAdder U2368 (w8389, w8278, IN73[25], w8390, w8391);
  FullAdder U2369 (w8391, w8280, IN74[24], w8392, w8393);
  FullAdder U2370 (w8393, w8282, IN75[23], w8394, w8395);
  FullAdder U2371 (w8395, w8284, IN76[22], w8396, w8397);
  FullAdder U2372 (w8397, w8286, IN77[21], w8398, w8399);
  FullAdder U2373 (w8399, w8288, IN78[20], w8400, w8401);
  FullAdder U2374 (w8401, w8290, IN79[19], w8402, w8403);
  FullAdder U2375 (w8403, w8292, IN80[18], w8404, w8405);
  FullAdder U2376 (w8405, w8294, IN81[17], w8406, w8407);
  FullAdder U2377 (w8407, w8296, IN82[16], w8408, w8409);
  FullAdder U2378 (w8409, w8298, IN83[15], w8410, w8411);
  FullAdder U2379 (w8411, w8300, IN84[14], w8412, w8413);
  FullAdder U2380 (w8413, w8302, IN85[13], w8414, w8415);
  FullAdder U2381 (w8415, w8304, IN86[12], w8416, w8417);
  FullAdder U2382 (w8417, w8306, IN87[11], w8418, w8419);
  FullAdder U2383 (w8419, w8308, IN88[10], w8420, w8421);
  FullAdder U2384 (w8421, w8310, IN89[9], w8422, w8423);
  FullAdder U2385 (w8423, w8312, IN90[8], w8424, w8425);
  FullAdder U2386 (w8425, w8314, IN91[7], w8426, w8427);
  FullAdder U2387 (w8427, w8316, IN92[6], w8428, w8429);
  FullAdder U2388 (w8429, w8318, IN93[5], w8430, w8431);
  FullAdder U2389 (w8431, w8320, IN94[4], w8432, w8433);
  FullAdder U2390 (w8433, w8322, IN95[3], w8434, w8435);
  FullAdder U2391 (w8435, w8324, IN96[2], w8436, w8437);
  FullAdder U2392 (w8437, w8326, IN97[1], w8438, w8439);
  FullAdder U2393 (w8439, w8327, IN98[0], w8440, w8441);
  HalfAdder U2394 (w8330, IN43[43], Out1[43], w8443);
  FullAdder U2395 (w8443, w8332, IN44[43], w8444, w8445);
  FullAdder U2396 (w8445, w8334, IN45[43], w8446, w8447);
  FullAdder U2397 (w8447, w8336, IN46[43], w8448, w8449);
  FullAdder U2398 (w8449, w8338, IN47[43], w8450, w8451);
  FullAdder U2399 (w8451, w8340, IN48[43], w8452, w8453);
  FullAdder U2400 (w8453, w8342, IN49[43], w8454, w8455);
  FullAdder U2401 (w8455, w8344, IN50[43], w8456, w8457);
  FullAdder U2402 (w8457, w8346, IN51[43], w8458, w8459);
  FullAdder U2403 (w8459, w8348, IN52[43], w8460, w8461);
  FullAdder U2404 (w8461, w8350, IN53[43], w8462, w8463);
  FullAdder U2405 (w8463, w8352, IN54[43], w8464, w8465);
  FullAdder U2406 (w8465, w8354, IN55[43], w8466, w8467);
  FullAdder U2407 (w8467, w8356, IN56[43], w8468, w8469);
  FullAdder U2408 (w8469, w8358, IN57[43], w8470, w8471);
  FullAdder U2409 (w8471, w8360, IN58[41], w8472, w8473);
  FullAdder U2410 (w8473, w8362, IN59[40], w8474, w8475);
  FullAdder U2411 (w8475, w8364, IN60[39], w8476, w8477);
  FullAdder U2412 (w8477, w8366, IN61[38], w8478, w8479);
  FullAdder U2413 (w8479, w8368, IN62[37], w8480, w8481);
  FullAdder U2414 (w8481, w8370, IN63[36], w8482, w8483);
  FullAdder U2415 (w8483, w8372, IN64[35], w8484, w8485);
  FullAdder U2416 (w8485, w8374, IN65[34], w8486, w8487);
  FullAdder U2417 (w8487, w8376, IN66[33], w8488, w8489);
  FullAdder U2418 (w8489, w8378, IN67[32], w8490, w8491);
  FullAdder U2419 (w8491, w8380, IN68[31], w8492, w8493);
  FullAdder U2420 (w8493, w8382, IN69[30], w8494, w8495);
  FullAdder U2421 (w8495, w8384, IN70[29], w8496, w8497);
  FullAdder U2422 (w8497, w8386, IN71[28], w8498, w8499);
  FullAdder U2423 (w8499, w8388, IN72[27], w8500, w8501);
  FullAdder U2424 (w8501, w8390, IN73[26], w8502, w8503);
  FullAdder U2425 (w8503, w8392, IN74[25], w8504, w8505);
  FullAdder U2426 (w8505, w8394, IN75[24], w8506, w8507);
  FullAdder U2427 (w8507, w8396, IN76[23], w8508, w8509);
  FullAdder U2428 (w8509, w8398, IN77[22], w8510, w8511);
  FullAdder U2429 (w8511, w8400, IN78[21], w8512, w8513);
  FullAdder U2430 (w8513, w8402, IN79[20], w8514, w8515);
  FullAdder U2431 (w8515, w8404, IN80[19], w8516, w8517);
  FullAdder U2432 (w8517, w8406, IN81[18], w8518, w8519);
  FullAdder U2433 (w8519, w8408, IN82[17], w8520, w8521);
  FullAdder U2434 (w8521, w8410, IN83[16], w8522, w8523);
  FullAdder U2435 (w8523, w8412, IN84[15], w8524, w8525);
  FullAdder U2436 (w8525, w8414, IN85[14], w8526, w8527);
  FullAdder U2437 (w8527, w8416, IN86[13], w8528, w8529);
  FullAdder U2438 (w8529, w8418, IN87[12], w8530, w8531);
  FullAdder U2439 (w8531, w8420, IN88[11], w8532, w8533);
  FullAdder U2440 (w8533, w8422, IN89[10], w8534, w8535);
  FullAdder U2441 (w8535, w8424, IN90[9], w8536, w8537);
  FullAdder U2442 (w8537, w8426, IN91[8], w8538, w8539);
  FullAdder U2443 (w8539, w8428, IN92[7], w8540, w8541);
  FullAdder U2444 (w8541, w8430, IN93[6], w8542, w8543);
  FullAdder U2445 (w8543, w8432, IN94[5], w8544, w8545);
  FullAdder U2446 (w8545, w8434, IN95[4], w8546, w8547);
  FullAdder U2447 (w8547, w8436, IN96[3], w8548, w8549);
  FullAdder U2448 (w8549, w8438, IN97[2], w8550, w8551);
  FullAdder U2449 (w8551, w8440, IN98[1], w8552, w8553);
  FullAdder U2450 (w8553, w8441, IN99[0], w8554, w8555);
  HalfAdder U2451 (w8444, IN44[44], Out1[44], w8557);
  FullAdder U2452 (w8557, w8446, IN45[44], w8558, w8559);
  FullAdder U2453 (w8559, w8448, IN46[44], w8560, w8561);
  FullAdder U2454 (w8561, w8450, IN47[44], w8562, w8563);
  FullAdder U2455 (w8563, w8452, IN48[44], w8564, w8565);
  FullAdder U2456 (w8565, w8454, IN49[44], w8566, w8567);
  FullAdder U2457 (w8567, w8456, IN50[44], w8568, w8569);
  FullAdder U2458 (w8569, w8458, IN51[44], w8570, w8571);
  FullAdder U2459 (w8571, w8460, IN52[44], w8572, w8573);
  FullAdder U2460 (w8573, w8462, IN53[44], w8574, w8575);
  FullAdder U2461 (w8575, w8464, IN54[44], w8576, w8577);
  FullAdder U2462 (w8577, w8466, IN55[44], w8578, w8579);
  FullAdder U2463 (w8579, w8468, IN56[44], w8580, w8581);
  FullAdder U2464 (w8581, w8470, IN57[44], w8582, w8583);
  FullAdder U2465 (w8583, w8472, IN58[42], w8584, w8585);
  FullAdder U2466 (w8585, w8474, IN59[41], w8586, w8587);
  FullAdder U2467 (w8587, w8476, IN60[40], w8588, w8589);
  FullAdder U2468 (w8589, w8478, IN61[39], w8590, w8591);
  FullAdder U2469 (w8591, w8480, IN62[38], w8592, w8593);
  FullAdder U2470 (w8593, w8482, IN63[37], w8594, w8595);
  FullAdder U2471 (w8595, w8484, IN64[36], w8596, w8597);
  FullAdder U2472 (w8597, w8486, IN65[35], w8598, w8599);
  FullAdder U2473 (w8599, w8488, IN66[34], w8600, w8601);
  FullAdder U2474 (w8601, w8490, IN67[33], w8602, w8603);
  FullAdder U2475 (w8603, w8492, IN68[32], w8604, w8605);
  FullAdder U2476 (w8605, w8494, IN69[31], w8606, w8607);
  FullAdder U2477 (w8607, w8496, IN70[30], w8608, w8609);
  FullAdder U2478 (w8609, w8498, IN71[29], w8610, w8611);
  FullAdder U2479 (w8611, w8500, IN72[28], w8612, w8613);
  FullAdder U2480 (w8613, w8502, IN73[27], w8614, w8615);
  FullAdder U2481 (w8615, w8504, IN74[26], w8616, w8617);
  FullAdder U2482 (w8617, w8506, IN75[25], w8618, w8619);
  FullAdder U2483 (w8619, w8508, IN76[24], w8620, w8621);
  FullAdder U2484 (w8621, w8510, IN77[23], w8622, w8623);
  FullAdder U2485 (w8623, w8512, IN78[22], w8624, w8625);
  FullAdder U2486 (w8625, w8514, IN79[21], w8626, w8627);
  FullAdder U2487 (w8627, w8516, IN80[20], w8628, w8629);
  FullAdder U2488 (w8629, w8518, IN81[19], w8630, w8631);
  FullAdder U2489 (w8631, w8520, IN82[18], w8632, w8633);
  FullAdder U2490 (w8633, w8522, IN83[17], w8634, w8635);
  FullAdder U2491 (w8635, w8524, IN84[16], w8636, w8637);
  FullAdder U2492 (w8637, w8526, IN85[15], w8638, w8639);
  FullAdder U2493 (w8639, w8528, IN86[14], w8640, w8641);
  FullAdder U2494 (w8641, w8530, IN87[13], w8642, w8643);
  FullAdder U2495 (w8643, w8532, IN88[12], w8644, w8645);
  FullAdder U2496 (w8645, w8534, IN89[11], w8646, w8647);
  FullAdder U2497 (w8647, w8536, IN90[10], w8648, w8649);
  FullAdder U2498 (w8649, w8538, IN91[9], w8650, w8651);
  FullAdder U2499 (w8651, w8540, IN92[8], w8652, w8653);
  FullAdder U2500 (w8653, w8542, IN93[7], w8654, w8655);
  FullAdder U2501 (w8655, w8544, IN94[6], w8656, w8657);
  FullAdder U2502 (w8657, w8546, IN95[5], w8658, w8659);
  FullAdder U2503 (w8659, w8548, IN96[4], w8660, w8661);
  FullAdder U2504 (w8661, w8550, IN97[3], w8662, w8663);
  FullAdder U2505 (w8663, w8552, IN98[2], w8664, w8665);
  FullAdder U2506 (w8665, w8554, IN99[1], w8666, w8667);
  FullAdder U2507 (w8667, w8555, IN100[0], w8668, w8669);
  HalfAdder U2508 (w8558, IN45[45], Out1[45], w8671);
  FullAdder U2509 (w8671, w8560, IN46[45], w8672, w8673);
  FullAdder U2510 (w8673, w8562, IN47[45], w8674, w8675);
  FullAdder U2511 (w8675, w8564, IN48[45], w8676, w8677);
  FullAdder U2512 (w8677, w8566, IN49[45], w8678, w8679);
  FullAdder U2513 (w8679, w8568, IN50[45], w8680, w8681);
  FullAdder U2514 (w8681, w8570, IN51[45], w8682, w8683);
  FullAdder U2515 (w8683, w8572, IN52[45], w8684, w8685);
  FullAdder U2516 (w8685, w8574, IN53[45], w8686, w8687);
  FullAdder U2517 (w8687, w8576, IN54[45], w8688, w8689);
  FullAdder U2518 (w8689, w8578, IN55[45], w8690, w8691);
  FullAdder U2519 (w8691, w8580, IN56[45], w8692, w8693);
  FullAdder U2520 (w8693, w8582, IN57[45], w8694, w8695);
  FullAdder U2521 (w8695, w8584, IN58[43], w8696, w8697);
  FullAdder U2522 (w8697, w8586, IN59[42], w8698, w8699);
  FullAdder U2523 (w8699, w8588, IN60[41], w8700, w8701);
  FullAdder U2524 (w8701, w8590, IN61[40], w8702, w8703);
  FullAdder U2525 (w8703, w8592, IN62[39], w8704, w8705);
  FullAdder U2526 (w8705, w8594, IN63[38], w8706, w8707);
  FullAdder U2527 (w8707, w8596, IN64[37], w8708, w8709);
  FullAdder U2528 (w8709, w8598, IN65[36], w8710, w8711);
  FullAdder U2529 (w8711, w8600, IN66[35], w8712, w8713);
  FullAdder U2530 (w8713, w8602, IN67[34], w8714, w8715);
  FullAdder U2531 (w8715, w8604, IN68[33], w8716, w8717);
  FullAdder U2532 (w8717, w8606, IN69[32], w8718, w8719);
  FullAdder U2533 (w8719, w8608, IN70[31], w8720, w8721);
  FullAdder U2534 (w8721, w8610, IN71[30], w8722, w8723);
  FullAdder U2535 (w8723, w8612, IN72[29], w8724, w8725);
  FullAdder U2536 (w8725, w8614, IN73[28], w8726, w8727);
  FullAdder U2537 (w8727, w8616, IN74[27], w8728, w8729);
  FullAdder U2538 (w8729, w8618, IN75[26], w8730, w8731);
  FullAdder U2539 (w8731, w8620, IN76[25], w8732, w8733);
  FullAdder U2540 (w8733, w8622, IN77[24], w8734, w8735);
  FullAdder U2541 (w8735, w8624, IN78[23], w8736, w8737);
  FullAdder U2542 (w8737, w8626, IN79[22], w8738, w8739);
  FullAdder U2543 (w8739, w8628, IN80[21], w8740, w8741);
  FullAdder U2544 (w8741, w8630, IN81[20], w8742, w8743);
  FullAdder U2545 (w8743, w8632, IN82[19], w8744, w8745);
  FullAdder U2546 (w8745, w8634, IN83[18], w8746, w8747);
  FullAdder U2547 (w8747, w8636, IN84[17], w8748, w8749);
  FullAdder U2548 (w8749, w8638, IN85[16], w8750, w8751);
  FullAdder U2549 (w8751, w8640, IN86[15], w8752, w8753);
  FullAdder U2550 (w8753, w8642, IN87[14], w8754, w8755);
  FullAdder U2551 (w8755, w8644, IN88[13], w8756, w8757);
  FullAdder U2552 (w8757, w8646, IN89[12], w8758, w8759);
  FullAdder U2553 (w8759, w8648, IN90[11], w8760, w8761);
  FullAdder U2554 (w8761, w8650, IN91[10], w8762, w8763);
  FullAdder U2555 (w8763, w8652, IN92[9], w8764, w8765);
  FullAdder U2556 (w8765, w8654, IN93[8], w8766, w8767);
  FullAdder U2557 (w8767, w8656, IN94[7], w8768, w8769);
  FullAdder U2558 (w8769, w8658, IN95[6], w8770, w8771);
  FullAdder U2559 (w8771, w8660, IN96[5], w8772, w8773);
  FullAdder U2560 (w8773, w8662, IN97[4], w8774, w8775);
  FullAdder U2561 (w8775, w8664, IN98[3], w8776, w8777);
  FullAdder U2562 (w8777, w8666, IN99[2], w8778, w8779);
  FullAdder U2563 (w8779, w8668, IN100[1], w8780, w8781);
  FullAdder U2564 (w8781, w8669, IN101[0], w8782, w8783);
  HalfAdder U2565 (w8672, IN46[46], Out1[46], w8785);
  FullAdder U2566 (w8785, w8674, IN47[46], w8786, w8787);
  FullAdder U2567 (w8787, w8676, IN48[46], w8788, w8789);
  FullAdder U2568 (w8789, w8678, IN49[46], w8790, w8791);
  FullAdder U2569 (w8791, w8680, IN50[46], w8792, w8793);
  FullAdder U2570 (w8793, w8682, IN51[46], w8794, w8795);
  FullAdder U2571 (w8795, w8684, IN52[46], w8796, w8797);
  FullAdder U2572 (w8797, w8686, IN53[46], w8798, w8799);
  FullAdder U2573 (w8799, w8688, IN54[46], w8800, w8801);
  FullAdder U2574 (w8801, w8690, IN55[46], w8802, w8803);
  FullAdder U2575 (w8803, w8692, IN56[46], w8804, w8805);
  FullAdder U2576 (w8805, w8694, IN57[46], w8806, w8807);
  FullAdder U2577 (w8807, w8696, IN58[44], w8808, w8809);
  FullAdder U2578 (w8809, w8698, IN59[43], w8810, w8811);
  FullAdder U2579 (w8811, w8700, IN60[42], w8812, w8813);
  FullAdder U2580 (w8813, w8702, IN61[41], w8814, w8815);
  FullAdder U2581 (w8815, w8704, IN62[40], w8816, w8817);
  FullAdder U2582 (w8817, w8706, IN63[39], w8818, w8819);
  FullAdder U2583 (w8819, w8708, IN64[38], w8820, w8821);
  FullAdder U2584 (w8821, w8710, IN65[37], w8822, w8823);
  FullAdder U2585 (w8823, w8712, IN66[36], w8824, w8825);
  FullAdder U2586 (w8825, w8714, IN67[35], w8826, w8827);
  FullAdder U2587 (w8827, w8716, IN68[34], w8828, w8829);
  FullAdder U2588 (w8829, w8718, IN69[33], w8830, w8831);
  FullAdder U2589 (w8831, w8720, IN70[32], w8832, w8833);
  FullAdder U2590 (w8833, w8722, IN71[31], w8834, w8835);
  FullAdder U2591 (w8835, w8724, IN72[30], w8836, w8837);
  FullAdder U2592 (w8837, w8726, IN73[29], w8838, w8839);
  FullAdder U2593 (w8839, w8728, IN74[28], w8840, w8841);
  FullAdder U2594 (w8841, w8730, IN75[27], w8842, w8843);
  FullAdder U2595 (w8843, w8732, IN76[26], w8844, w8845);
  FullAdder U2596 (w8845, w8734, IN77[25], w8846, w8847);
  FullAdder U2597 (w8847, w8736, IN78[24], w8848, w8849);
  FullAdder U2598 (w8849, w8738, IN79[23], w8850, w8851);
  FullAdder U2599 (w8851, w8740, IN80[22], w8852, w8853);
  FullAdder U2600 (w8853, w8742, IN81[21], w8854, w8855);
  FullAdder U2601 (w8855, w8744, IN82[20], w8856, w8857);
  FullAdder U2602 (w8857, w8746, IN83[19], w8858, w8859);
  FullAdder U2603 (w8859, w8748, IN84[18], w8860, w8861);
  FullAdder U2604 (w8861, w8750, IN85[17], w8862, w8863);
  FullAdder U2605 (w8863, w8752, IN86[16], w8864, w8865);
  FullAdder U2606 (w8865, w8754, IN87[15], w8866, w8867);
  FullAdder U2607 (w8867, w8756, IN88[14], w8868, w8869);
  FullAdder U2608 (w8869, w8758, IN89[13], w8870, w8871);
  FullAdder U2609 (w8871, w8760, IN90[12], w8872, w8873);
  FullAdder U2610 (w8873, w8762, IN91[11], w8874, w8875);
  FullAdder U2611 (w8875, w8764, IN92[10], w8876, w8877);
  FullAdder U2612 (w8877, w8766, IN93[9], w8878, w8879);
  FullAdder U2613 (w8879, w8768, IN94[8], w8880, w8881);
  FullAdder U2614 (w8881, w8770, IN95[7], w8882, w8883);
  FullAdder U2615 (w8883, w8772, IN96[6], w8884, w8885);
  FullAdder U2616 (w8885, w8774, IN97[5], w8886, w8887);
  FullAdder U2617 (w8887, w8776, IN98[4], w8888, w8889);
  FullAdder U2618 (w8889, w8778, IN99[3], w8890, w8891);
  FullAdder U2619 (w8891, w8780, IN100[2], w8892, w8893);
  FullAdder U2620 (w8893, w8782, IN101[1], w8894, w8895);
  FullAdder U2621 (w8895, w8783, IN102[0], w8896, w8897);
  HalfAdder U2622 (w8786, IN47[47], Out1[47], w8899);
  FullAdder U2623 (w8899, w8788, IN48[47], w8900, w8901);
  FullAdder U2624 (w8901, w8790, IN49[47], w8902, w8903);
  FullAdder U2625 (w8903, w8792, IN50[47], w8904, w8905);
  FullAdder U2626 (w8905, w8794, IN51[47], w8906, w8907);
  FullAdder U2627 (w8907, w8796, IN52[47], w8908, w8909);
  FullAdder U2628 (w8909, w8798, IN53[47], w8910, w8911);
  FullAdder U2629 (w8911, w8800, IN54[47], w8912, w8913);
  FullAdder U2630 (w8913, w8802, IN55[47], w8914, w8915);
  FullAdder U2631 (w8915, w8804, IN56[47], w8916, w8917);
  FullAdder U2632 (w8917, w8806, IN57[47], w8918, w8919);
  FullAdder U2633 (w8919, w8808, IN58[45], w8920, w8921);
  FullAdder U2634 (w8921, w8810, IN59[44], w8922, w8923);
  FullAdder U2635 (w8923, w8812, IN60[43], w8924, w8925);
  FullAdder U2636 (w8925, w8814, IN61[42], w8926, w8927);
  FullAdder U2637 (w8927, w8816, IN62[41], w8928, w8929);
  FullAdder U2638 (w8929, w8818, IN63[40], w8930, w8931);
  FullAdder U2639 (w8931, w8820, IN64[39], w8932, w8933);
  FullAdder U2640 (w8933, w8822, IN65[38], w8934, w8935);
  FullAdder U2641 (w8935, w8824, IN66[37], w8936, w8937);
  FullAdder U2642 (w8937, w8826, IN67[36], w8938, w8939);
  FullAdder U2643 (w8939, w8828, IN68[35], w8940, w8941);
  FullAdder U2644 (w8941, w8830, IN69[34], w8942, w8943);
  FullAdder U2645 (w8943, w8832, IN70[33], w8944, w8945);
  FullAdder U2646 (w8945, w8834, IN71[32], w8946, w8947);
  FullAdder U2647 (w8947, w8836, IN72[31], w8948, w8949);
  FullAdder U2648 (w8949, w8838, IN73[30], w8950, w8951);
  FullAdder U2649 (w8951, w8840, IN74[29], w8952, w8953);
  FullAdder U2650 (w8953, w8842, IN75[28], w8954, w8955);
  FullAdder U2651 (w8955, w8844, IN76[27], w8956, w8957);
  FullAdder U2652 (w8957, w8846, IN77[26], w8958, w8959);
  FullAdder U2653 (w8959, w8848, IN78[25], w8960, w8961);
  FullAdder U2654 (w8961, w8850, IN79[24], w8962, w8963);
  FullAdder U2655 (w8963, w8852, IN80[23], w8964, w8965);
  FullAdder U2656 (w8965, w8854, IN81[22], w8966, w8967);
  FullAdder U2657 (w8967, w8856, IN82[21], w8968, w8969);
  FullAdder U2658 (w8969, w8858, IN83[20], w8970, w8971);
  FullAdder U2659 (w8971, w8860, IN84[19], w8972, w8973);
  FullAdder U2660 (w8973, w8862, IN85[18], w8974, w8975);
  FullAdder U2661 (w8975, w8864, IN86[17], w8976, w8977);
  FullAdder U2662 (w8977, w8866, IN87[16], w8978, w8979);
  FullAdder U2663 (w8979, w8868, IN88[15], w8980, w8981);
  FullAdder U2664 (w8981, w8870, IN89[14], w8982, w8983);
  FullAdder U2665 (w8983, w8872, IN90[13], w8984, w8985);
  FullAdder U2666 (w8985, w8874, IN91[12], w8986, w8987);
  FullAdder U2667 (w8987, w8876, IN92[11], w8988, w8989);
  FullAdder U2668 (w8989, w8878, IN93[10], w8990, w8991);
  FullAdder U2669 (w8991, w8880, IN94[9], w8992, w8993);
  FullAdder U2670 (w8993, w8882, IN95[8], w8994, w8995);
  FullAdder U2671 (w8995, w8884, IN96[7], w8996, w8997);
  FullAdder U2672 (w8997, w8886, IN97[6], w8998, w8999);
  FullAdder U2673 (w8999, w8888, IN98[5], w9000, w9001);
  FullAdder U2674 (w9001, w8890, IN99[4], w9002, w9003);
  FullAdder U2675 (w9003, w8892, IN100[3], w9004, w9005);
  FullAdder U2676 (w9005, w8894, IN101[2], w9006, w9007);
  FullAdder U2677 (w9007, w8896, IN102[1], w9008, w9009);
  FullAdder U2678 (w9009, w8897, IN103[0], w9010, w9011);
  HalfAdder U2679 (w8900, IN48[48], Out1[48], w9013);
  FullAdder U2680 (w9013, w8902, IN49[48], w9014, w9015);
  FullAdder U2681 (w9015, w8904, IN50[48], w9016, w9017);
  FullAdder U2682 (w9017, w8906, IN51[48], w9018, w9019);
  FullAdder U2683 (w9019, w8908, IN52[48], w9020, w9021);
  FullAdder U2684 (w9021, w8910, IN53[48], w9022, w9023);
  FullAdder U2685 (w9023, w8912, IN54[48], w9024, w9025);
  FullAdder U2686 (w9025, w8914, IN55[48], w9026, w9027);
  FullAdder U2687 (w9027, w8916, IN56[48], w9028, w9029);
  FullAdder U2688 (w9029, w8918, IN57[48], w9030, w9031);
  FullAdder U2689 (w9031, w8920, IN58[46], w9032, w9033);
  FullAdder U2690 (w9033, w8922, IN59[45], w9034, w9035);
  FullAdder U2691 (w9035, w8924, IN60[44], w9036, w9037);
  FullAdder U2692 (w9037, w8926, IN61[43], w9038, w9039);
  FullAdder U2693 (w9039, w8928, IN62[42], w9040, w9041);
  FullAdder U2694 (w9041, w8930, IN63[41], w9042, w9043);
  FullAdder U2695 (w9043, w8932, IN64[40], w9044, w9045);
  FullAdder U2696 (w9045, w8934, IN65[39], w9046, w9047);
  FullAdder U2697 (w9047, w8936, IN66[38], w9048, w9049);
  FullAdder U2698 (w9049, w8938, IN67[37], w9050, w9051);
  FullAdder U2699 (w9051, w8940, IN68[36], w9052, w9053);
  FullAdder U2700 (w9053, w8942, IN69[35], w9054, w9055);
  FullAdder U2701 (w9055, w8944, IN70[34], w9056, w9057);
  FullAdder U2702 (w9057, w8946, IN71[33], w9058, w9059);
  FullAdder U2703 (w9059, w8948, IN72[32], w9060, w9061);
  FullAdder U2704 (w9061, w8950, IN73[31], w9062, w9063);
  FullAdder U2705 (w9063, w8952, IN74[30], w9064, w9065);
  FullAdder U2706 (w9065, w8954, IN75[29], w9066, w9067);
  FullAdder U2707 (w9067, w8956, IN76[28], w9068, w9069);
  FullAdder U2708 (w9069, w8958, IN77[27], w9070, w9071);
  FullAdder U2709 (w9071, w8960, IN78[26], w9072, w9073);
  FullAdder U2710 (w9073, w8962, IN79[25], w9074, w9075);
  FullAdder U2711 (w9075, w8964, IN80[24], w9076, w9077);
  FullAdder U2712 (w9077, w8966, IN81[23], w9078, w9079);
  FullAdder U2713 (w9079, w8968, IN82[22], w9080, w9081);
  FullAdder U2714 (w9081, w8970, IN83[21], w9082, w9083);
  FullAdder U2715 (w9083, w8972, IN84[20], w9084, w9085);
  FullAdder U2716 (w9085, w8974, IN85[19], w9086, w9087);
  FullAdder U2717 (w9087, w8976, IN86[18], w9088, w9089);
  FullAdder U2718 (w9089, w8978, IN87[17], w9090, w9091);
  FullAdder U2719 (w9091, w8980, IN88[16], w9092, w9093);
  FullAdder U2720 (w9093, w8982, IN89[15], w9094, w9095);
  FullAdder U2721 (w9095, w8984, IN90[14], w9096, w9097);
  FullAdder U2722 (w9097, w8986, IN91[13], w9098, w9099);
  FullAdder U2723 (w9099, w8988, IN92[12], w9100, w9101);
  FullAdder U2724 (w9101, w8990, IN93[11], w9102, w9103);
  FullAdder U2725 (w9103, w8992, IN94[10], w9104, w9105);
  FullAdder U2726 (w9105, w8994, IN95[9], w9106, w9107);
  FullAdder U2727 (w9107, w8996, IN96[8], w9108, w9109);
  FullAdder U2728 (w9109, w8998, IN97[7], w9110, w9111);
  FullAdder U2729 (w9111, w9000, IN98[6], w9112, w9113);
  FullAdder U2730 (w9113, w9002, IN99[5], w9114, w9115);
  FullAdder U2731 (w9115, w9004, IN100[4], w9116, w9117);
  FullAdder U2732 (w9117, w9006, IN101[3], w9118, w9119);
  FullAdder U2733 (w9119, w9008, IN102[2], w9120, w9121);
  FullAdder U2734 (w9121, w9010, IN103[1], w9122, w9123);
  FullAdder U2735 (w9123, w9011, IN104[0], w9124, w9125);
  HalfAdder U2736 (w9014, IN49[49], Out1[49], w9127);
  FullAdder U2737 (w9127, w9016, IN50[49], w9128, w9129);
  FullAdder U2738 (w9129, w9018, IN51[49], w9130, w9131);
  FullAdder U2739 (w9131, w9020, IN52[49], w9132, w9133);
  FullAdder U2740 (w9133, w9022, IN53[49], w9134, w9135);
  FullAdder U2741 (w9135, w9024, IN54[49], w9136, w9137);
  FullAdder U2742 (w9137, w9026, IN55[49], w9138, w9139);
  FullAdder U2743 (w9139, w9028, IN56[49], w9140, w9141);
  FullAdder U2744 (w9141, w9030, IN57[49], w9142, w9143);
  FullAdder U2745 (w9143, w9032, IN58[47], w9144, w9145);
  FullAdder U2746 (w9145, w9034, IN59[46], w9146, w9147);
  FullAdder U2747 (w9147, w9036, IN60[45], w9148, w9149);
  FullAdder U2748 (w9149, w9038, IN61[44], w9150, w9151);
  FullAdder U2749 (w9151, w9040, IN62[43], w9152, w9153);
  FullAdder U2750 (w9153, w9042, IN63[42], w9154, w9155);
  FullAdder U2751 (w9155, w9044, IN64[41], w9156, w9157);
  FullAdder U2752 (w9157, w9046, IN65[40], w9158, w9159);
  FullAdder U2753 (w9159, w9048, IN66[39], w9160, w9161);
  FullAdder U2754 (w9161, w9050, IN67[38], w9162, w9163);
  FullAdder U2755 (w9163, w9052, IN68[37], w9164, w9165);
  FullAdder U2756 (w9165, w9054, IN69[36], w9166, w9167);
  FullAdder U2757 (w9167, w9056, IN70[35], w9168, w9169);
  FullAdder U2758 (w9169, w9058, IN71[34], w9170, w9171);
  FullAdder U2759 (w9171, w9060, IN72[33], w9172, w9173);
  FullAdder U2760 (w9173, w9062, IN73[32], w9174, w9175);
  FullAdder U2761 (w9175, w9064, IN74[31], w9176, w9177);
  FullAdder U2762 (w9177, w9066, IN75[30], w9178, w9179);
  FullAdder U2763 (w9179, w9068, IN76[29], w9180, w9181);
  FullAdder U2764 (w9181, w9070, IN77[28], w9182, w9183);
  FullAdder U2765 (w9183, w9072, IN78[27], w9184, w9185);
  FullAdder U2766 (w9185, w9074, IN79[26], w9186, w9187);
  FullAdder U2767 (w9187, w9076, IN80[25], w9188, w9189);
  FullAdder U2768 (w9189, w9078, IN81[24], w9190, w9191);
  FullAdder U2769 (w9191, w9080, IN82[23], w9192, w9193);
  FullAdder U2770 (w9193, w9082, IN83[22], w9194, w9195);
  FullAdder U2771 (w9195, w9084, IN84[21], w9196, w9197);
  FullAdder U2772 (w9197, w9086, IN85[20], w9198, w9199);
  FullAdder U2773 (w9199, w9088, IN86[19], w9200, w9201);
  FullAdder U2774 (w9201, w9090, IN87[18], w9202, w9203);
  FullAdder U2775 (w9203, w9092, IN88[17], w9204, w9205);
  FullAdder U2776 (w9205, w9094, IN89[16], w9206, w9207);
  FullAdder U2777 (w9207, w9096, IN90[15], w9208, w9209);
  FullAdder U2778 (w9209, w9098, IN91[14], w9210, w9211);
  FullAdder U2779 (w9211, w9100, IN92[13], w9212, w9213);
  FullAdder U2780 (w9213, w9102, IN93[12], w9214, w9215);
  FullAdder U2781 (w9215, w9104, IN94[11], w9216, w9217);
  FullAdder U2782 (w9217, w9106, IN95[10], w9218, w9219);
  FullAdder U2783 (w9219, w9108, IN96[9], w9220, w9221);
  FullAdder U2784 (w9221, w9110, IN97[8], w9222, w9223);
  FullAdder U2785 (w9223, w9112, IN98[7], w9224, w9225);
  FullAdder U2786 (w9225, w9114, IN99[6], w9226, w9227);
  FullAdder U2787 (w9227, w9116, IN100[5], w9228, w9229);
  FullAdder U2788 (w9229, w9118, IN101[4], w9230, w9231);
  FullAdder U2789 (w9231, w9120, IN102[3], w9232, w9233);
  FullAdder U2790 (w9233, w9122, IN103[2], w9234, w9235);
  FullAdder U2791 (w9235, w9124, IN104[1], w9236, w9237);
  FullAdder U2792 (w9237, w9125, IN105[0], w9238, w9239);
  HalfAdder U2793 (w9128, IN50[50], Out1[50], w9241);
  FullAdder U2794 (w9241, w9130, IN51[50], w9242, w9243);
  FullAdder U2795 (w9243, w9132, IN52[50], w9244, w9245);
  FullAdder U2796 (w9245, w9134, IN53[50], w9246, w9247);
  FullAdder U2797 (w9247, w9136, IN54[50], w9248, w9249);
  FullAdder U2798 (w9249, w9138, IN55[50], w9250, w9251);
  FullAdder U2799 (w9251, w9140, IN56[50], w9252, w9253);
  FullAdder U2800 (w9253, w9142, IN57[50], w9254, w9255);
  FullAdder U2801 (w9255, w9144, IN58[48], w9256, w9257);
  FullAdder U2802 (w9257, w9146, IN59[47], w9258, w9259);
  FullAdder U2803 (w9259, w9148, IN60[46], w9260, w9261);
  FullAdder U2804 (w9261, w9150, IN61[45], w9262, w9263);
  FullAdder U2805 (w9263, w9152, IN62[44], w9264, w9265);
  FullAdder U2806 (w9265, w9154, IN63[43], w9266, w9267);
  FullAdder U2807 (w9267, w9156, IN64[42], w9268, w9269);
  FullAdder U2808 (w9269, w9158, IN65[41], w9270, w9271);
  FullAdder U2809 (w9271, w9160, IN66[40], w9272, w9273);
  FullAdder U2810 (w9273, w9162, IN67[39], w9274, w9275);
  FullAdder U2811 (w9275, w9164, IN68[38], w9276, w9277);
  FullAdder U2812 (w9277, w9166, IN69[37], w9278, w9279);
  FullAdder U2813 (w9279, w9168, IN70[36], w9280, w9281);
  FullAdder U2814 (w9281, w9170, IN71[35], w9282, w9283);
  FullAdder U2815 (w9283, w9172, IN72[34], w9284, w9285);
  FullAdder U2816 (w9285, w9174, IN73[33], w9286, w9287);
  FullAdder U2817 (w9287, w9176, IN74[32], w9288, w9289);
  FullAdder U2818 (w9289, w9178, IN75[31], w9290, w9291);
  FullAdder U2819 (w9291, w9180, IN76[30], w9292, w9293);
  FullAdder U2820 (w9293, w9182, IN77[29], w9294, w9295);
  FullAdder U2821 (w9295, w9184, IN78[28], w9296, w9297);
  FullAdder U2822 (w9297, w9186, IN79[27], w9298, w9299);
  FullAdder U2823 (w9299, w9188, IN80[26], w9300, w9301);
  FullAdder U2824 (w9301, w9190, IN81[25], w9302, w9303);
  FullAdder U2825 (w9303, w9192, IN82[24], w9304, w9305);
  FullAdder U2826 (w9305, w9194, IN83[23], w9306, w9307);
  FullAdder U2827 (w9307, w9196, IN84[22], w9308, w9309);
  FullAdder U2828 (w9309, w9198, IN85[21], w9310, w9311);
  FullAdder U2829 (w9311, w9200, IN86[20], w9312, w9313);
  FullAdder U2830 (w9313, w9202, IN87[19], w9314, w9315);
  FullAdder U2831 (w9315, w9204, IN88[18], w9316, w9317);
  FullAdder U2832 (w9317, w9206, IN89[17], w9318, w9319);
  FullAdder U2833 (w9319, w9208, IN90[16], w9320, w9321);
  FullAdder U2834 (w9321, w9210, IN91[15], w9322, w9323);
  FullAdder U2835 (w9323, w9212, IN92[14], w9324, w9325);
  FullAdder U2836 (w9325, w9214, IN93[13], w9326, w9327);
  FullAdder U2837 (w9327, w9216, IN94[12], w9328, w9329);
  FullAdder U2838 (w9329, w9218, IN95[11], w9330, w9331);
  FullAdder U2839 (w9331, w9220, IN96[10], w9332, w9333);
  FullAdder U2840 (w9333, w9222, IN97[9], w9334, w9335);
  FullAdder U2841 (w9335, w9224, IN98[8], w9336, w9337);
  FullAdder U2842 (w9337, w9226, IN99[7], w9338, w9339);
  FullAdder U2843 (w9339, w9228, IN100[6], w9340, w9341);
  FullAdder U2844 (w9341, w9230, IN101[5], w9342, w9343);
  FullAdder U2845 (w9343, w9232, IN102[4], w9344, w9345);
  FullAdder U2846 (w9345, w9234, IN103[3], w9346, w9347);
  FullAdder U2847 (w9347, w9236, IN104[2], w9348, w9349);
  FullAdder U2848 (w9349, w9238, IN105[1], w9350, w9351);
  FullAdder U2849 (w9351, w9239, IN106[0], w9352, w9353);
  HalfAdder U2850 (w9242, IN51[51], Out1[51], w9355);
  FullAdder U2851 (w9355, w9244, IN52[51], w9356, w9357);
  FullAdder U2852 (w9357, w9246, IN53[51], w9358, w9359);
  FullAdder U2853 (w9359, w9248, IN54[51], w9360, w9361);
  FullAdder U2854 (w9361, w9250, IN55[51], w9362, w9363);
  FullAdder U2855 (w9363, w9252, IN56[51], w9364, w9365);
  FullAdder U2856 (w9365, w9254, IN57[51], w9366, w9367);
  FullAdder U2857 (w9367, w9256, IN58[49], w9368, w9369);
  FullAdder U2858 (w9369, w9258, IN59[48], w9370, w9371);
  FullAdder U2859 (w9371, w9260, IN60[47], w9372, w9373);
  FullAdder U2860 (w9373, w9262, IN61[46], w9374, w9375);
  FullAdder U2861 (w9375, w9264, IN62[45], w9376, w9377);
  FullAdder U2862 (w9377, w9266, IN63[44], w9378, w9379);
  FullAdder U2863 (w9379, w9268, IN64[43], w9380, w9381);
  FullAdder U2864 (w9381, w9270, IN65[42], w9382, w9383);
  FullAdder U2865 (w9383, w9272, IN66[41], w9384, w9385);
  FullAdder U2866 (w9385, w9274, IN67[40], w9386, w9387);
  FullAdder U2867 (w9387, w9276, IN68[39], w9388, w9389);
  FullAdder U2868 (w9389, w9278, IN69[38], w9390, w9391);
  FullAdder U2869 (w9391, w9280, IN70[37], w9392, w9393);
  FullAdder U2870 (w9393, w9282, IN71[36], w9394, w9395);
  FullAdder U2871 (w9395, w9284, IN72[35], w9396, w9397);
  FullAdder U2872 (w9397, w9286, IN73[34], w9398, w9399);
  FullAdder U2873 (w9399, w9288, IN74[33], w9400, w9401);
  FullAdder U2874 (w9401, w9290, IN75[32], w9402, w9403);
  FullAdder U2875 (w9403, w9292, IN76[31], w9404, w9405);
  FullAdder U2876 (w9405, w9294, IN77[30], w9406, w9407);
  FullAdder U2877 (w9407, w9296, IN78[29], w9408, w9409);
  FullAdder U2878 (w9409, w9298, IN79[28], w9410, w9411);
  FullAdder U2879 (w9411, w9300, IN80[27], w9412, w9413);
  FullAdder U2880 (w9413, w9302, IN81[26], w9414, w9415);
  FullAdder U2881 (w9415, w9304, IN82[25], w9416, w9417);
  FullAdder U2882 (w9417, w9306, IN83[24], w9418, w9419);
  FullAdder U2883 (w9419, w9308, IN84[23], w9420, w9421);
  FullAdder U2884 (w9421, w9310, IN85[22], w9422, w9423);
  FullAdder U2885 (w9423, w9312, IN86[21], w9424, w9425);
  FullAdder U2886 (w9425, w9314, IN87[20], w9426, w9427);
  FullAdder U2887 (w9427, w9316, IN88[19], w9428, w9429);
  FullAdder U2888 (w9429, w9318, IN89[18], w9430, w9431);
  FullAdder U2889 (w9431, w9320, IN90[17], w9432, w9433);
  FullAdder U2890 (w9433, w9322, IN91[16], w9434, w9435);
  FullAdder U2891 (w9435, w9324, IN92[15], w9436, w9437);
  FullAdder U2892 (w9437, w9326, IN93[14], w9438, w9439);
  FullAdder U2893 (w9439, w9328, IN94[13], w9440, w9441);
  FullAdder U2894 (w9441, w9330, IN95[12], w9442, w9443);
  FullAdder U2895 (w9443, w9332, IN96[11], w9444, w9445);
  FullAdder U2896 (w9445, w9334, IN97[10], w9446, w9447);
  FullAdder U2897 (w9447, w9336, IN98[9], w9448, w9449);
  FullAdder U2898 (w9449, w9338, IN99[8], w9450, w9451);
  FullAdder U2899 (w9451, w9340, IN100[7], w9452, w9453);
  FullAdder U2900 (w9453, w9342, IN101[6], w9454, w9455);
  FullAdder U2901 (w9455, w9344, IN102[5], w9456, w9457);
  FullAdder U2902 (w9457, w9346, IN103[4], w9458, w9459);
  FullAdder U2903 (w9459, w9348, IN104[3], w9460, w9461);
  FullAdder U2904 (w9461, w9350, IN105[2], w9462, w9463);
  FullAdder U2905 (w9463, w9352, IN106[1], w9464, w9465);
  FullAdder U2906 (w9465, w9353, IN107[0], w9466, w9467);
  HalfAdder U2907 (w9356, IN52[52], Out1[52], w9469);
  FullAdder U2908 (w9469, w9358, IN53[52], w9470, w9471);
  FullAdder U2909 (w9471, w9360, IN54[52], w9472, w9473);
  FullAdder U2910 (w9473, w9362, IN55[52], w9474, w9475);
  FullAdder U2911 (w9475, w9364, IN56[52], w9476, w9477);
  FullAdder U2912 (w9477, w9366, IN57[52], w9478, w9479);
  FullAdder U2913 (w9479, w9368, IN58[50], w9480, w9481);
  FullAdder U2914 (w9481, w9370, IN59[49], w9482, w9483);
  FullAdder U2915 (w9483, w9372, IN60[48], w9484, w9485);
  FullAdder U2916 (w9485, w9374, IN61[47], w9486, w9487);
  FullAdder U2917 (w9487, w9376, IN62[46], w9488, w9489);
  FullAdder U2918 (w9489, w9378, IN63[45], w9490, w9491);
  FullAdder U2919 (w9491, w9380, IN64[44], w9492, w9493);
  FullAdder U2920 (w9493, w9382, IN65[43], w9494, w9495);
  FullAdder U2921 (w9495, w9384, IN66[42], w9496, w9497);
  FullAdder U2922 (w9497, w9386, IN67[41], w9498, w9499);
  FullAdder U2923 (w9499, w9388, IN68[40], w9500, w9501);
  FullAdder U2924 (w9501, w9390, IN69[39], w9502, w9503);
  FullAdder U2925 (w9503, w9392, IN70[38], w9504, w9505);
  FullAdder U2926 (w9505, w9394, IN71[37], w9506, w9507);
  FullAdder U2927 (w9507, w9396, IN72[36], w9508, w9509);
  FullAdder U2928 (w9509, w9398, IN73[35], w9510, w9511);
  FullAdder U2929 (w9511, w9400, IN74[34], w9512, w9513);
  FullAdder U2930 (w9513, w9402, IN75[33], w9514, w9515);
  FullAdder U2931 (w9515, w9404, IN76[32], w9516, w9517);
  FullAdder U2932 (w9517, w9406, IN77[31], w9518, w9519);
  FullAdder U2933 (w9519, w9408, IN78[30], w9520, w9521);
  FullAdder U2934 (w9521, w9410, IN79[29], w9522, w9523);
  FullAdder U2935 (w9523, w9412, IN80[28], w9524, w9525);
  FullAdder U2936 (w9525, w9414, IN81[27], w9526, w9527);
  FullAdder U2937 (w9527, w9416, IN82[26], w9528, w9529);
  FullAdder U2938 (w9529, w9418, IN83[25], w9530, w9531);
  FullAdder U2939 (w9531, w9420, IN84[24], w9532, w9533);
  FullAdder U2940 (w9533, w9422, IN85[23], w9534, w9535);
  FullAdder U2941 (w9535, w9424, IN86[22], w9536, w9537);
  FullAdder U2942 (w9537, w9426, IN87[21], w9538, w9539);
  FullAdder U2943 (w9539, w9428, IN88[20], w9540, w9541);
  FullAdder U2944 (w9541, w9430, IN89[19], w9542, w9543);
  FullAdder U2945 (w9543, w9432, IN90[18], w9544, w9545);
  FullAdder U2946 (w9545, w9434, IN91[17], w9546, w9547);
  FullAdder U2947 (w9547, w9436, IN92[16], w9548, w9549);
  FullAdder U2948 (w9549, w9438, IN93[15], w9550, w9551);
  FullAdder U2949 (w9551, w9440, IN94[14], w9552, w9553);
  FullAdder U2950 (w9553, w9442, IN95[13], w9554, w9555);
  FullAdder U2951 (w9555, w9444, IN96[12], w9556, w9557);
  FullAdder U2952 (w9557, w9446, IN97[11], w9558, w9559);
  FullAdder U2953 (w9559, w9448, IN98[10], w9560, w9561);
  FullAdder U2954 (w9561, w9450, IN99[9], w9562, w9563);
  FullAdder U2955 (w9563, w9452, IN100[8], w9564, w9565);
  FullAdder U2956 (w9565, w9454, IN101[7], w9566, w9567);
  FullAdder U2957 (w9567, w9456, IN102[6], w9568, w9569);
  FullAdder U2958 (w9569, w9458, IN103[5], w9570, w9571);
  FullAdder U2959 (w9571, w9460, IN104[4], w9572, w9573);
  FullAdder U2960 (w9573, w9462, IN105[3], w9574, w9575);
  FullAdder U2961 (w9575, w9464, IN106[2], w9576, w9577);
  FullAdder U2962 (w9577, w9466, IN107[1], w9578, w9579);
  FullAdder U2963 (w9579, w9467, IN108[0], w9580, w9581);
  HalfAdder U2964 (w9470, IN53[53], Out1[53], w9583);
  FullAdder U2965 (w9583, w9472, IN54[53], w9584, w9585);
  FullAdder U2966 (w9585, w9474, IN55[53], w9586, w9587);
  FullAdder U2967 (w9587, w9476, IN56[53], w9588, w9589);
  FullAdder U2968 (w9589, w9478, IN57[53], w9590, w9591);
  FullAdder U2969 (w9591, w9480, IN58[51], w9592, w9593);
  FullAdder U2970 (w9593, w9482, IN59[50], w9594, w9595);
  FullAdder U2971 (w9595, w9484, IN60[49], w9596, w9597);
  FullAdder U2972 (w9597, w9486, IN61[48], w9598, w9599);
  FullAdder U2973 (w9599, w9488, IN62[47], w9600, w9601);
  FullAdder U2974 (w9601, w9490, IN63[46], w9602, w9603);
  FullAdder U2975 (w9603, w9492, IN64[45], w9604, w9605);
  FullAdder U2976 (w9605, w9494, IN65[44], w9606, w9607);
  FullAdder U2977 (w9607, w9496, IN66[43], w9608, w9609);
  FullAdder U2978 (w9609, w9498, IN67[42], w9610, w9611);
  FullAdder U2979 (w9611, w9500, IN68[41], w9612, w9613);
  FullAdder U2980 (w9613, w9502, IN69[40], w9614, w9615);
  FullAdder U2981 (w9615, w9504, IN70[39], w9616, w9617);
  FullAdder U2982 (w9617, w9506, IN71[38], w9618, w9619);
  FullAdder U2983 (w9619, w9508, IN72[37], w9620, w9621);
  FullAdder U2984 (w9621, w9510, IN73[36], w9622, w9623);
  FullAdder U2985 (w9623, w9512, IN74[35], w9624, w9625);
  FullAdder U2986 (w9625, w9514, IN75[34], w9626, w9627);
  FullAdder U2987 (w9627, w9516, IN76[33], w9628, w9629);
  FullAdder U2988 (w9629, w9518, IN77[32], w9630, w9631);
  FullAdder U2989 (w9631, w9520, IN78[31], w9632, w9633);
  FullAdder U2990 (w9633, w9522, IN79[30], w9634, w9635);
  FullAdder U2991 (w9635, w9524, IN80[29], w9636, w9637);
  FullAdder U2992 (w9637, w9526, IN81[28], w9638, w9639);
  FullAdder U2993 (w9639, w9528, IN82[27], w9640, w9641);
  FullAdder U2994 (w9641, w9530, IN83[26], w9642, w9643);
  FullAdder U2995 (w9643, w9532, IN84[25], w9644, w9645);
  FullAdder U2996 (w9645, w9534, IN85[24], w9646, w9647);
  FullAdder U2997 (w9647, w9536, IN86[23], w9648, w9649);
  FullAdder U2998 (w9649, w9538, IN87[22], w9650, w9651);
  FullAdder U2999 (w9651, w9540, IN88[21], w9652, w9653);
  FullAdder U3000 (w9653, w9542, IN89[20], w9654, w9655);
  FullAdder U3001 (w9655, w9544, IN90[19], w9656, w9657);
  FullAdder U3002 (w9657, w9546, IN91[18], w9658, w9659);
  FullAdder U3003 (w9659, w9548, IN92[17], w9660, w9661);
  FullAdder U3004 (w9661, w9550, IN93[16], w9662, w9663);
  FullAdder U3005 (w9663, w9552, IN94[15], w9664, w9665);
  FullAdder U3006 (w9665, w9554, IN95[14], w9666, w9667);
  FullAdder U3007 (w9667, w9556, IN96[13], w9668, w9669);
  FullAdder U3008 (w9669, w9558, IN97[12], w9670, w9671);
  FullAdder U3009 (w9671, w9560, IN98[11], w9672, w9673);
  FullAdder U3010 (w9673, w9562, IN99[10], w9674, w9675);
  FullAdder U3011 (w9675, w9564, IN100[9], w9676, w9677);
  FullAdder U3012 (w9677, w9566, IN101[8], w9678, w9679);
  FullAdder U3013 (w9679, w9568, IN102[7], w9680, w9681);
  FullAdder U3014 (w9681, w9570, IN103[6], w9682, w9683);
  FullAdder U3015 (w9683, w9572, IN104[5], w9684, w9685);
  FullAdder U3016 (w9685, w9574, IN105[4], w9686, w9687);
  FullAdder U3017 (w9687, w9576, IN106[3], w9688, w9689);
  FullAdder U3018 (w9689, w9578, IN107[2], w9690, w9691);
  FullAdder U3019 (w9691, w9580, IN108[1], w9692, w9693);
  FullAdder U3020 (w9693, w9581, IN109[0], w9694, w9695);
  HalfAdder U3021 (w9584, IN54[54], Out1[54], w9697);
  FullAdder U3022 (w9697, w9586, IN55[54], w9698, w9699);
  FullAdder U3023 (w9699, w9588, IN56[54], w9700, w9701);
  FullAdder U3024 (w9701, w9590, IN57[54], w9702, w9703);
  FullAdder U3025 (w9703, w9592, IN58[52], w9704, w9705);
  FullAdder U3026 (w9705, w9594, IN59[51], w9706, w9707);
  FullAdder U3027 (w9707, w9596, IN60[50], w9708, w9709);
  FullAdder U3028 (w9709, w9598, IN61[49], w9710, w9711);
  FullAdder U3029 (w9711, w9600, IN62[48], w9712, w9713);
  FullAdder U3030 (w9713, w9602, IN63[47], w9714, w9715);
  FullAdder U3031 (w9715, w9604, IN64[46], w9716, w9717);
  FullAdder U3032 (w9717, w9606, IN65[45], w9718, w9719);
  FullAdder U3033 (w9719, w9608, IN66[44], w9720, w9721);
  FullAdder U3034 (w9721, w9610, IN67[43], w9722, w9723);
  FullAdder U3035 (w9723, w9612, IN68[42], w9724, w9725);
  FullAdder U3036 (w9725, w9614, IN69[41], w9726, w9727);
  FullAdder U3037 (w9727, w9616, IN70[40], w9728, w9729);
  FullAdder U3038 (w9729, w9618, IN71[39], w9730, w9731);
  FullAdder U3039 (w9731, w9620, IN72[38], w9732, w9733);
  FullAdder U3040 (w9733, w9622, IN73[37], w9734, w9735);
  FullAdder U3041 (w9735, w9624, IN74[36], w9736, w9737);
  FullAdder U3042 (w9737, w9626, IN75[35], w9738, w9739);
  FullAdder U3043 (w9739, w9628, IN76[34], w9740, w9741);
  FullAdder U3044 (w9741, w9630, IN77[33], w9742, w9743);
  FullAdder U3045 (w9743, w9632, IN78[32], w9744, w9745);
  FullAdder U3046 (w9745, w9634, IN79[31], w9746, w9747);
  FullAdder U3047 (w9747, w9636, IN80[30], w9748, w9749);
  FullAdder U3048 (w9749, w9638, IN81[29], w9750, w9751);
  FullAdder U3049 (w9751, w9640, IN82[28], w9752, w9753);
  FullAdder U3050 (w9753, w9642, IN83[27], w9754, w9755);
  FullAdder U3051 (w9755, w9644, IN84[26], w9756, w9757);
  FullAdder U3052 (w9757, w9646, IN85[25], w9758, w9759);
  FullAdder U3053 (w9759, w9648, IN86[24], w9760, w9761);
  FullAdder U3054 (w9761, w9650, IN87[23], w9762, w9763);
  FullAdder U3055 (w9763, w9652, IN88[22], w9764, w9765);
  FullAdder U3056 (w9765, w9654, IN89[21], w9766, w9767);
  FullAdder U3057 (w9767, w9656, IN90[20], w9768, w9769);
  FullAdder U3058 (w9769, w9658, IN91[19], w9770, w9771);
  FullAdder U3059 (w9771, w9660, IN92[18], w9772, w9773);
  FullAdder U3060 (w9773, w9662, IN93[17], w9774, w9775);
  FullAdder U3061 (w9775, w9664, IN94[16], w9776, w9777);
  FullAdder U3062 (w9777, w9666, IN95[15], w9778, w9779);
  FullAdder U3063 (w9779, w9668, IN96[14], w9780, w9781);
  FullAdder U3064 (w9781, w9670, IN97[13], w9782, w9783);
  FullAdder U3065 (w9783, w9672, IN98[12], w9784, w9785);
  FullAdder U3066 (w9785, w9674, IN99[11], w9786, w9787);
  FullAdder U3067 (w9787, w9676, IN100[10], w9788, w9789);
  FullAdder U3068 (w9789, w9678, IN101[9], w9790, w9791);
  FullAdder U3069 (w9791, w9680, IN102[8], w9792, w9793);
  FullAdder U3070 (w9793, w9682, IN103[7], w9794, w9795);
  FullAdder U3071 (w9795, w9684, IN104[6], w9796, w9797);
  FullAdder U3072 (w9797, w9686, IN105[5], w9798, w9799);
  FullAdder U3073 (w9799, w9688, IN106[4], w9800, w9801);
  FullAdder U3074 (w9801, w9690, IN107[3], w9802, w9803);
  FullAdder U3075 (w9803, w9692, IN108[2], w9804, w9805);
  FullAdder U3076 (w9805, w9694, IN109[1], w9806, w9807);
  FullAdder U3077 (w9807, w9695, IN110[0], w9808, w9809);
  HalfAdder U3078 (w9698, IN55[55], Out1[55], w9811);
  FullAdder U3079 (w9811, w9700, IN56[55], w9812, w9813);
  FullAdder U3080 (w9813, w9702, IN57[55], w9814, w9815);
  FullAdder U3081 (w9815, w9704, IN58[53], w9816, w9817);
  FullAdder U3082 (w9817, w9706, IN59[52], w9818, w9819);
  FullAdder U3083 (w9819, w9708, IN60[51], w9820, w9821);
  FullAdder U3084 (w9821, w9710, IN61[50], w9822, w9823);
  FullAdder U3085 (w9823, w9712, IN62[49], w9824, w9825);
  FullAdder U3086 (w9825, w9714, IN63[48], w9826, w9827);
  FullAdder U3087 (w9827, w9716, IN64[47], w9828, w9829);
  FullAdder U3088 (w9829, w9718, IN65[46], w9830, w9831);
  FullAdder U3089 (w9831, w9720, IN66[45], w9832, w9833);
  FullAdder U3090 (w9833, w9722, IN67[44], w9834, w9835);
  FullAdder U3091 (w9835, w9724, IN68[43], w9836, w9837);
  FullAdder U3092 (w9837, w9726, IN69[42], w9838, w9839);
  FullAdder U3093 (w9839, w9728, IN70[41], w9840, w9841);
  FullAdder U3094 (w9841, w9730, IN71[40], w9842, w9843);
  FullAdder U3095 (w9843, w9732, IN72[39], w9844, w9845);
  FullAdder U3096 (w9845, w9734, IN73[38], w9846, w9847);
  FullAdder U3097 (w9847, w9736, IN74[37], w9848, w9849);
  FullAdder U3098 (w9849, w9738, IN75[36], w9850, w9851);
  FullAdder U3099 (w9851, w9740, IN76[35], w9852, w9853);
  FullAdder U3100 (w9853, w9742, IN77[34], w9854, w9855);
  FullAdder U3101 (w9855, w9744, IN78[33], w9856, w9857);
  FullAdder U3102 (w9857, w9746, IN79[32], w9858, w9859);
  FullAdder U3103 (w9859, w9748, IN80[31], w9860, w9861);
  FullAdder U3104 (w9861, w9750, IN81[30], w9862, w9863);
  FullAdder U3105 (w9863, w9752, IN82[29], w9864, w9865);
  FullAdder U3106 (w9865, w9754, IN83[28], w9866, w9867);
  FullAdder U3107 (w9867, w9756, IN84[27], w9868, w9869);
  FullAdder U3108 (w9869, w9758, IN85[26], w9870, w9871);
  FullAdder U3109 (w9871, w9760, IN86[25], w9872, w9873);
  FullAdder U3110 (w9873, w9762, IN87[24], w9874, w9875);
  FullAdder U3111 (w9875, w9764, IN88[23], w9876, w9877);
  FullAdder U3112 (w9877, w9766, IN89[22], w9878, w9879);
  FullAdder U3113 (w9879, w9768, IN90[21], w9880, w9881);
  FullAdder U3114 (w9881, w9770, IN91[20], w9882, w9883);
  FullAdder U3115 (w9883, w9772, IN92[19], w9884, w9885);
  FullAdder U3116 (w9885, w9774, IN93[18], w9886, w9887);
  FullAdder U3117 (w9887, w9776, IN94[17], w9888, w9889);
  FullAdder U3118 (w9889, w9778, IN95[16], w9890, w9891);
  FullAdder U3119 (w9891, w9780, IN96[15], w9892, w9893);
  FullAdder U3120 (w9893, w9782, IN97[14], w9894, w9895);
  FullAdder U3121 (w9895, w9784, IN98[13], w9896, w9897);
  FullAdder U3122 (w9897, w9786, IN99[12], w9898, w9899);
  FullAdder U3123 (w9899, w9788, IN100[11], w9900, w9901);
  FullAdder U3124 (w9901, w9790, IN101[10], w9902, w9903);
  FullAdder U3125 (w9903, w9792, IN102[9], w9904, w9905);
  FullAdder U3126 (w9905, w9794, IN103[8], w9906, w9907);
  FullAdder U3127 (w9907, w9796, IN104[7], w9908, w9909);
  FullAdder U3128 (w9909, w9798, IN105[6], w9910, w9911);
  FullAdder U3129 (w9911, w9800, IN106[5], w9912, w9913);
  FullAdder U3130 (w9913, w9802, IN107[4], w9914, w9915);
  FullAdder U3131 (w9915, w9804, IN108[3], w9916, w9917);
  FullAdder U3132 (w9917, w9806, IN109[2], w9918, w9919);
  FullAdder U3133 (w9919, w9808, IN110[1], w9920, w9921);
  FullAdder U3134 (w9921, w9809, IN111[0], w9922, w9923);
  HalfAdder U3135 (w9812, IN56[56], Out1[56], w9925);
  FullAdder U3136 (w9925, w9814, IN57[56], w9926, w9927);
  FullAdder U3137 (w9927, w9816, IN58[54], w9928, w9929);
  FullAdder U3138 (w9929, w9818, IN59[53], w9930, w9931);
  FullAdder U3139 (w9931, w9820, IN60[52], w9932, w9933);
  FullAdder U3140 (w9933, w9822, IN61[51], w9934, w9935);
  FullAdder U3141 (w9935, w9824, IN62[50], w9936, w9937);
  FullAdder U3142 (w9937, w9826, IN63[49], w9938, w9939);
  FullAdder U3143 (w9939, w9828, IN64[48], w9940, w9941);
  FullAdder U3144 (w9941, w9830, IN65[47], w9942, w9943);
  FullAdder U3145 (w9943, w9832, IN66[46], w9944, w9945);
  FullAdder U3146 (w9945, w9834, IN67[45], w9946, w9947);
  FullAdder U3147 (w9947, w9836, IN68[44], w9948, w9949);
  FullAdder U3148 (w9949, w9838, IN69[43], w9950, w9951);
  FullAdder U3149 (w9951, w9840, IN70[42], w9952, w9953);
  FullAdder U3150 (w9953, w9842, IN71[41], w9954, w9955);
  FullAdder U3151 (w9955, w9844, IN72[40], w9956, w9957);
  FullAdder U3152 (w9957, w9846, IN73[39], w9958, w9959);
  FullAdder U3153 (w9959, w9848, IN74[38], w9960, w9961);
  FullAdder U3154 (w9961, w9850, IN75[37], w9962, w9963);
  FullAdder U3155 (w9963, w9852, IN76[36], w9964, w9965);
  FullAdder U3156 (w9965, w9854, IN77[35], w9966, w9967);
  FullAdder U3157 (w9967, w9856, IN78[34], w9968, w9969);
  FullAdder U3158 (w9969, w9858, IN79[33], w9970, w9971);
  FullAdder U3159 (w9971, w9860, IN80[32], w9972, w9973);
  FullAdder U3160 (w9973, w9862, IN81[31], w9974, w9975);
  FullAdder U3161 (w9975, w9864, IN82[30], w9976, w9977);
  FullAdder U3162 (w9977, w9866, IN83[29], w9978, w9979);
  FullAdder U3163 (w9979, w9868, IN84[28], w9980, w9981);
  FullAdder U3164 (w9981, w9870, IN85[27], w9982, w9983);
  FullAdder U3165 (w9983, w9872, IN86[26], w9984, w9985);
  FullAdder U3166 (w9985, w9874, IN87[25], w9986, w9987);
  FullAdder U3167 (w9987, w9876, IN88[24], w9988, w9989);
  FullAdder U3168 (w9989, w9878, IN89[23], w9990, w9991);
  FullAdder U3169 (w9991, w9880, IN90[22], w9992, w9993);
  FullAdder U3170 (w9993, w9882, IN91[21], w9994, w9995);
  FullAdder U3171 (w9995, w9884, IN92[20], w9996, w9997);
  FullAdder U3172 (w9997, w9886, IN93[19], w9998, w9999);
  FullAdder U3173 (w9999, w9888, IN94[18], w10000, w10001);
  FullAdder U3174 (w10001, w9890, IN95[17], w10002, w10003);
  FullAdder U3175 (w10003, w9892, IN96[16], w10004, w10005);
  FullAdder U3176 (w10005, w9894, IN97[15], w10006, w10007);
  FullAdder U3177 (w10007, w9896, IN98[14], w10008, w10009);
  FullAdder U3178 (w10009, w9898, IN99[13], w10010, w10011);
  FullAdder U3179 (w10011, w9900, IN100[12], w10012, w10013);
  FullAdder U3180 (w10013, w9902, IN101[11], w10014, w10015);
  FullAdder U3181 (w10015, w9904, IN102[10], w10016, w10017);
  FullAdder U3182 (w10017, w9906, IN103[9], w10018, w10019);
  FullAdder U3183 (w10019, w9908, IN104[8], w10020, w10021);
  FullAdder U3184 (w10021, w9910, IN105[7], w10022, w10023);
  FullAdder U3185 (w10023, w9912, IN106[6], w10024, w10025);
  FullAdder U3186 (w10025, w9914, IN107[5], w10026, w10027);
  FullAdder U3187 (w10027, w9916, IN108[4], w10028, w10029);
  FullAdder U3188 (w10029, w9918, IN109[3], w10030, w10031);
  FullAdder U3189 (w10031, w9920, IN110[2], w10032, w10033);
  FullAdder U3190 (w10033, w9922, IN111[1], w10034, w10035);
  FullAdder U3191 (w10035, w9923, IN112[0], w10036, w10037);
  HalfAdder U3192 (w9926, IN57[57], Out1[57], w10039);
  FullAdder U3193 (w10039, w9928, IN58[55], w10040, w10041);
  FullAdder U3194 (w10041, w9930, IN59[54], w10042, w10043);
  FullAdder U3195 (w10043, w9932, IN60[53], w10044, w10045);
  FullAdder U3196 (w10045, w9934, IN61[52], w10046, w10047);
  FullAdder U3197 (w10047, w9936, IN62[51], w10048, w10049);
  FullAdder U3198 (w10049, w9938, IN63[50], w10050, w10051);
  FullAdder U3199 (w10051, w9940, IN64[49], w10052, w10053);
  FullAdder U3200 (w10053, w9942, IN65[48], w10054, w10055);
  FullAdder U3201 (w10055, w9944, IN66[47], w10056, w10057);
  FullAdder U3202 (w10057, w9946, IN67[46], w10058, w10059);
  FullAdder U3203 (w10059, w9948, IN68[45], w10060, w10061);
  FullAdder U3204 (w10061, w9950, IN69[44], w10062, w10063);
  FullAdder U3205 (w10063, w9952, IN70[43], w10064, w10065);
  FullAdder U3206 (w10065, w9954, IN71[42], w10066, w10067);
  FullAdder U3207 (w10067, w9956, IN72[41], w10068, w10069);
  FullAdder U3208 (w10069, w9958, IN73[40], w10070, w10071);
  FullAdder U3209 (w10071, w9960, IN74[39], w10072, w10073);
  FullAdder U3210 (w10073, w9962, IN75[38], w10074, w10075);
  FullAdder U3211 (w10075, w9964, IN76[37], w10076, w10077);
  FullAdder U3212 (w10077, w9966, IN77[36], w10078, w10079);
  FullAdder U3213 (w10079, w9968, IN78[35], w10080, w10081);
  FullAdder U3214 (w10081, w9970, IN79[34], w10082, w10083);
  FullAdder U3215 (w10083, w9972, IN80[33], w10084, w10085);
  FullAdder U3216 (w10085, w9974, IN81[32], w10086, w10087);
  FullAdder U3217 (w10087, w9976, IN82[31], w10088, w10089);
  FullAdder U3218 (w10089, w9978, IN83[30], w10090, w10091);
  FullAdder U3219 (w10091, w9980, IN84[29], w10092, w10093);
  FullAdder U3220 (w10093, w9982, IN85[28], w10094, w10095);
  FullAdder U3221 (w10095, w9984, IN86[27], w10096, w10097);
  FullAdder U3222 (w10097, w9986, IN87[26], w10098, w10099);
  FullAdder U3223 (w10099, w9988, IN88[25], w10100, w10101);
  FullAdder U3224 (w10101, w9990, IN89[24], w10102, w10103);
  FullAdder U3225 (w10103, w9992, IN90[23], w10104, w10105);
  FullAdder U3226 (w10105, w9994, IN91[22], w10106, w10107);
  FullAdder U3227 (w10107, w9996, IN92[21], w10108, w10109);
  FullAdder U3228 (w10109, w9998, IN93[20], w10110, w10111);
  FullAdder U3229 (w10111, w10000, IN94[19], w10112, w10113);
  FullAdder U3230 (w10113, w10002, IN95[18], w10114, w10115);
  FullAdder U3231 (w10115, w10004, IN96[17], w10116, w10117);
  FullAdder U3232 (w10117, w10006, IN97[16], w10118, w10119);
  FullAdder U3233 (w10119, w10008, IN98[15], w10120, w10121);
  FullAdder U3234 (w10121, w10010, IN99[14], w10122, w10123);
  FullAdder U3235 (w10123, w10012, IN100[13], w10124, w10125);
  FullAdder U3236 (w10125, w10014, IN101[12], w10126, w10127);
  FullAdder U3237 (w10127, w10016, IN102[11], w10128, w10129);
  FullAdder U3238 (w10129, w10018, IN103[10], w10130, w10131);
  FullAdder U3239 (w10131, w10020, IN104[9], w10132, w10133);
  FullAdder U3240 (w10133, w10022, IN105[8], w10134, w10135);
  FullAdder U3241 (w10135, w10024, IN106[7], w10136, w10137);
  FullAdder U3242 (w10137, w10026, IN107[6], w10138, w10139);
  FullAdder U3243 (w10139, w10028, IN108[5], w10140, w10141);
  FullAdder U3244 (w10141, w10030, IN109[4], w10142, w10143);
  FullAdder U3245 (w10143, w10032, IN110[3], w10144, w10145);
  FullAdder U3246 (w10145, w10034, IN111[2], w10146, w10147);
  FullAdder U3247 (w10147, w10036, IN112[1], w10148, w10149);
  FullAdder U3248 (w10149, w10037, IN113[0], w10150, w10151);
  HalfAdder U3249 (w10040, IN58[56], Out1[58], w10153);
  FullAdder U3250 (w10153, w10042, IN59[55], w10154, w10155);
  FullAdder U3251 (w10155, w10044, IN60[54], w10156, w10157);
  FullAdder U3252 (w10157, w10046, IN61[53], w10158, w10159);
  FullAdder U3253 (w10159, w10048, IN62[52], w10160, w10161);
  FullAdder U3254 (w10161, w10050, IN63[51], w10162, w10163);
  FullAdder U3255 (w10163, w10052, IN64[50], w10164, w10165);
  FullAdder U3256 (w10165, w10054, IN65[49], w10166, w10167);
  FullAdder U3257 (w10167, w10056, IN66[48], w10168, w10169);
  FullAdder U3258 (w10169, w10058, IN67[47], w10170, w10171);
  FullAdder U3259 (w10171, w10060, IN68[46], w10172, w10173);
  FullAdder U3260 (w10173, w10062, IN69[45], w10174, w10175);
  FullAdder U3261 (w10175, w10064, IN70[44], w10176, w10177);
  FullAdder U3262 (w10177, w10066, IN71[43], w10178, w10179);
  FullAdder U3263 (w10179, w10068, IN72[42], w10180, w10181);
  FullAdder U3264 (w10181, w10070, IN73[41], w10182, w10183);
  FullAdder U3265 (w10183, w10072, IN74[40], w10184, w10185);
  FullAdder U3266 (w10185, w10074, IN75[39], w10186, w10187);
  FullAdder U3267 (w10187, w10076, IN76[38], w10188, w10189);
  FullAdder U3268 (w10189, w10078, IN77[37], w10190, w10191);
  FullAdder U3269 (w10191, w10080, IN78[36], w10192, w10193);
  FullAdder U3270 (w10193, w10082, IN79[35], w10194, w10195);
  FullAdder U3271 (w10195, w10084, IN80[34], w10196, w10197);
  FullAdder U3272 (w10197, w10086, IN81[33], w10198, w10199);
  FullAdder U3273 (w10199, w10088, IN82[32], w10200, w10201);
  FullAdder U3274 (w10201, w10090, IN83[31], w10202, w10203);
  FullAdder U3275 (w10203, w10092, IN84[30], w10204, w10205);
  FullAdder U3276 (w10205, w10094, IN85[29], w10206, w10207);
  FullAdder U3277 (w10207, w10096, IN86[28], w10208, w10209);
  FullAdder U3278 (w10209, w10098, IN87[27], w10210, w10211);
  FullAdder U3279 (w10211, w10100, IN88[26], w10212, w10213);
  FullAdder U3280 (w10213, w10102, IN89[25], w10214, w10215);
  FullAdder U3281 (w10215, w10104, IN90[24], w10216, w10217);
  FullAdder U3282 (w10217, w10106, IN91[23], w10218, w10219);
  FullAdder U3283 (w10219, w10108, IN92[22], w10220, w10221);
  FullAdder U3284 (w10221, w10110, IN93[21], w10222, w10223);
  FullAdder U3285 (w10223, w10112, IN94[20], w10224, w10225);
  FullAdder U3286 (w10225, w10114, IN95[19], w10226, w10227);
  FullAdder U3287 (w10227, w10116, IN96[18], w10228, w10229);
  FullAdder U3288 (w10229, w10118, IN97[17], w10230, w10231);
  FullAdder U3289 (w10231, w10120, IN98[16], w10232, w10233);
  FullAdder U3290 (w10233, w10122, IN99[15], w10234, w10235);
  FullAdder U3291 (w10235, w10124, IN100[14], w10236, w10237);
  FullAdder U3292 (w10237, w10126, IN101[13], w10238, w10239);
  FullAdder U3293 (w10239, w10128, IN102[12], w10240, w10241);
  FullAdder U3294 (w10241, w10130, IN103[11], w10242, w10243);
  FullAdder U3295 (w10243, w10132, IN104[10], w10244, w10245);
  FullAdder U3296 (w10245, w10134, IN105[9], w10246, w10247);
  FullAdder U3297 (w10247, w10136, IN106[8], w10248, w10249);
  FullAdder U3298 (w10249, w10138, IN107[7], w10250, w10251);
  FullAdder U3299 (w10251, w10140, IN108[6], w10252, w10253);
  FullAdder U3300 (w10253, w10142, IN109[5], w10254, w10255);
  FullAdder U3301 (w10255, w10144, IN110[4], w10256, w10257);
  FullAdder U3302 (w10257, w10146, IN111[3], w10258, w10259);
  FullAdder U3303 (w10259, w10148, IN112[2], w10260, w10261);
  FullAdder U3304 (w10261, w10150, IN113[1], w10262, w10263);
  FullAdder U3305 (w10263, w10151, IN114[0], w10264, w10265);
  HalfAdder U3306 (w10154, IN59[56], Out1[59], w10267);
  FullAdder U3307 (w10267, w10156, IN60[55], w10268, w10269);
  FullAdder U3308 (w10269, w10158, IN61[54], w10270, w10271);
  FullAdder U3309 (w10271, w10160, IN62[53], w10272, w10273);
  FullAdder U3310 (w10273, w10162, IN63[52], w10274, w10275);
  FullAdder U3311 (w10275, w10164, IN64[51], w10276, w10277);
  FullAdder U3312 (w10277, w10166, IN65[50], w10278, w10279);
  FullAdder U3313 (w10279, w10168, IN66[49], w10280, w10281);
  FullAdder U3314 (w10281, w10170, IN67[48], w10282, w10283);
  FullAdder U3315 (w10283, w10172, IN68[47], w10284, w10285);
  FullAdder U3316 (w10285, w10174, IN69[46], w10286, w10287);
  FullAdder U3317 (w10287, w10176, IN70[45], w10288, w10289);
  FullAdder U3318 (w10289, w10178, IN71[44], w10290, w10291);
  FullAdder U3319 (w10291, w10180, IN72[43], w10292, w10293);
  FullAdder U3320 (w10293, w10182, IN73[42], w10294, w10295);
  FullAdder U3321 (w10295, w10184, IN74[41], w10296, w10297);
  FullAdder U3322 (w10297, w10186, IN75[40], w10298, w10299);
  FullAdder U3323 (w10299, w10188, IN76[39], w10300, w10301);
  FullAdder U3324 (w10301, w10190, IN77[38], w10302, w10303);
  FullAdder U3325 (w10303, w10192, IN78[37], w10304, w10305);
  FullAdder U3326 (w10305, w10194, IN79[36], w10306, w10307);
  FullAdder U3327 (w10307, w10196, IN80[35], w10308, w10309);
  FullAdder U3328 (w10309, w10198, IN81[34], w10310, w10311);
  FullAdder U3329 (w10311, w10200, IN82[33], w10312, w10313);
  FullAdder U3330 (w10313, w10202, IN83[32], w10314, w10315);
  FullAdder U3331 (w10315, w10204, IN84[31], w10316, w10317);
  FullAdder U3332 (w10317, w10206, IN85[30], w10318, w10319);
  FullAdder U3333 (w10319, w10208, IN86[29], w10320, w10321);
  FullAdder U3334 (w10321, w10210, IN87[28], w10322, w10323);
  FullAdder U3335 (w10323, w10212, IN88[27], w10324, w10325);
  FullAdder U3336 (w10325, w10214, IN89[26], w10326, w10327);
  FullAdder U3337 (w10327, w10216, IN90[25], w10328, w10329);
  FullAdder U3338 (w10329, w10218, IN91[24], w10330, w10331);
  FullAdder U3339 (w10331, w10220, IN92[23], w10332, w10333);
  FullAdder U3340 (w10333, w10222, IN93[22], w10334, w10335);
  FullAdder U3341 (w10335, w10224, IN94[21], w10336, w10337);
  FullAdder U3342 (w10337, w10226, IN95[20], w10338, w10339);
  FullAdder U3343 (w10339, w10228, IN96[19], w10340, w10341);
  FullAdder U3344 (w10341, w10230, IN97[18], w10342, w10343);
  FullAdder U3345 (w10343, w10232, IN98[17], w10344, w10345);
  FullAdder U3346 (w10345, w10234, IN99[16], w10346, w10347);
  FullAdder U3347 (w10347, w10236, IN100[15], w10348, w10349);
  FullAdder U3348 (w10349, w10238, IN101[14], w10350, w10351);
  FullAdder U3349 (w10351, w10240, IN102[13], w10352, w10353);
  FullAdder U3350 (w10353, w10242, IN103[12], w10354, w10355);
  FullAdder U3351 (w10355, w10244, IN104[11], w10356, w10357);
  FullAdder U3352 (w10357, w10246, IN105[10], w10358, w10359);
  FullAdder U3353 (w10359, w10248, IN106[9], w10360, w10361);
  FullAdder U3354 (w10361, w10250, IN107[8], w10362, w10363);
  FullAdder U3355 (w10363, w10252, IN108[7], w10364, w10365);
  FullAdder U3356 (w10365, w10254, IN109[6], w10366, w10367);
  FullAdder U3357 (w10367, w10256, IN110[5], w10368, w10369);
  FullAdder U3358 (w10369, w10258, IN111[4], w10370, w10371);
  FullAdder U3359 (w10371, w10260, IN112[3], w10372, w10373);
  FullAdder U3360 (w10373, w10262, IN113[2], w10374, w10375);
  FullAdder U3361 (w10375, w10264, IN114[1], w10376, w10377);
  FullAdder U3362 (w10377, w10265, IN115[0], w10378, w10379);
  HalfAdder U3363 (w10268, IN60[56], Out1[60], w10381);
  FullAdder U3364 (w10381, w10270, IN61[55], w10382, w10383);
  FullAdder U3365 (w10383, w10272, IN62[54], w10384, w10385);
  FullAdder U3366 (w10385, w10274, IN63[53], w10386, w10387);
  FullAdder U3367 (w10387, w10276, IN64[52], w10388, w10389);
  FullAdder U3368 (w10389, w10278, IN65[51], w10390, w10391);
  FullAdder U3369 (w10391, w10280, IN66[50], w10392, w10393);
  FullAdder U3370 (w10393, w10282, IN67[49], w10394, w10395);
  FullAdder U3371 (w10395, w10284, IN68[48], w10396, w10397);
  FullAdder U3372 (w10397, w10286, IN69[47], w10398, w10399);
  FullAdder U3373 (w10399, w10288, IN70[46], w10400, w10401);
  FullAdder U3374 (w10401, w10290, IN71[45], w10402, w10403);
  FullAdder U3375 (w10403, w10292, IN72[44], w10404, w10405);
  FullAdder U3376 (w10405, w10294, IN73[43], w10406, w10407);
  FullAdder U3377 (w10407, w10296, IN74[42], w10408, w10409);
  FullAdder U3378 (w10409, w10298, IN75[41], w10410, w10411);
  FullAdder U3379 (w10411, w10300, IN76[40], w10412, w10413);
  FullAdder U3380 (w10413, w10302, IN77[39], w10414, w10415);
  FullAdder U3381 (w10415, w10304, IN78[38], w10416, w10417);
  FullAdder U3382 (w10417, w10306, IN79[37], w10418, w10419);
  FullAdder U3383 (w10419, w10308, IN80[36], w10420, w10421);
  FullAdder U3384 (w10421, w10310, IN81[35], w10422, w10423);
  FullAdder U3385 (w10423, w10312, IN82[34], w10424, w10425);
  FullAdder U3386 (w10425, w10314, IN83[33], w10426, w10427);
  FullAdder U3387 (w10427, w10316, IN84[32], w10428, w10429);
  FullAdder U3388 (w10429, w10318, IN85[31], w10430, w10431);
  FullAdder U3389 (w10431, w10320, IN86[30], w10432, w10433);
  FullAdder U3390 (w10433, w10322, IN87[29], w10434, w10435);
  FullAdder U3391 (w10435, w10324, IN88[28], w10436, w10437);
  FullAdder U3392 (w10437, w10326, IN89[27], w10438, w10439);
  FullAdder U3393 (w10439, w10328, IN90[26], w10440, w10441);
  FullAdder U3394 (w10441, w10330, IN91[25], w10442, w10443);
  FullAdder U3395 (w10443, w10332, IN92[24], w10444, w10445);
  FullAdder U3396 (w10445, w10334, IN93[23], w10446, w10447);
  FullAdder U3397 (w10447, w10336, IN94[22], w10448, w10449);
  FullAdder U3398 (w10449, w10338, IN95[21], w10450, w10451);
  FullAdder U3399 (w10451, w10340, IN96[20], w10452, w10453);
  FullAdder U3400 (w10453, w10342, IN97[19], w10454, w10455);
  FullAdder U3401 (w10455, w10344, IN98[18], w10456, w10457);
  FullAdder U3402 (w10457, w10346, IN99[17], w10458, w10459);
  FullAdder U3403 (w10459, w10348, IN100[16], w10460, w10461);
  FullAdder U3404 (w10461, w10350, IN101[15], w10462, w10463);
  FullAdder U3405 (w10463, w10352, IN102[14], w10464, w10465);
  FullAdder U3406 (w10465, w10354, IN103[13], w10466, w10467);
  FullAdder U3407 (w10467, w10356, IN104[12], w10468, w10469);
  FullAdder U3408 (w10469, w10358, IN105[11], w10470, w10471);
  FullAdder U3409 (w10471, w10360, IN106[10], w10472, w10473);
  FullAdder U3410 (w10473, w10362, IN107[9], w10474, w10475);
  FullAdder U3411 (w10475, w10364, IN108[8], w10476, w10477);
  FullAdder U3412 (w10477, w10366, IN109[7], w10478, w10479);
  FullAdder U3413 (w10479, w10368, IN110[6], w10480, w10481);
  FullAdder U3414 (w10481, w10370, IN111[5], w10482, w10483);
  FullAdder U3415 (w10483, w10372, IN112[4], w10484, w10485);
  FullAdder U3416 (w10485, w10374, IN113[3], w10486, w10487);
  FullAdder U3417 (w10487, w10376, IN114[2], w10488, w10489);
  FullAdder U3418 (w10489, w10378, IN115[1], w10490, w10491);
  FullAdder U3419 (w10491, w10379, IN116[0], w10492, w10493);
  HalfAdder U3420 (w10382, IN61[56], Out1[61], w10495);
  FullAdder U3421 (w10495, w10384, IN62[55], w10496, w10497);
  FullAdder U3422 (w10497, w10386, IN63[54], w10498, w10499);
  FullAdder U3423 (w10499, w10388, IN64[53], w10500, w10501);
  FullAdder U3424 (w10501, w10390, IN65[52], w10502, w10503);
  FullAdder U3425 (w10503, w10392, IN66[51], w10504, w10505);
  FullAdder U3426 (w10505, w10394, IN67[50], w10506, w10507);
  FullAdder U3427 (w10507, w10396, IN68[49], w10508, w10509);
  FullAdder U3428 (w10509, w10398, IN69[48], w10510, w10511);
  FullAdder U3429 (w10511, w10400, IN70[47], w10512, w10513);
  FullAdder U3430 (w10513, w10402, IN71[46], w10514, w10515);
  FullAdder U3431 (w10515, w10404, IN72[45], w10516, w10517);
  FullAdder U3432 (w10517, w10406, IN73[44], w10518, w10519);
  FullAdder U3433 (w10519, w10408, IN74[43], w10520, w10521);
  FullAdder U3434 (w10521, w10410, IN75[42], w10522, w10523);
  FullAdder U3435 (w10523, w10412, IN76[41], w10524, w10525);
  FullAdder U3436 (w10525, w10414, IN77[40], w10526, w10527);
  FullAdder U3437 (w10527, w10416, IN78[39], w10528, w10529);
  FullAdder U3438 (w10529, w10418, IN79[38], w10530, w10531);
  FullAdder U3439 (w10531, w10420, IN80[37], w10532, w10533);
  FullAdder U3440 (w10533, w10422, IN81[36], w10534, w10535);
  FullAdder U3441 (w10535, w10424, IN82[35], w10536, w10537);
  FullAdder U3442 (w10537, w10426, IN83[34], w10538, w10539);
  FullAdder U3443 (w10539, w10428, IN84[33], w10540, w10541);
  FullAdder U3444 (w10541, w10430, IN85[32], w10542, w10543);
  FullAdder U3445 (w10543, w10432, IN86[31], w10544, w10545);
  FullAdder U3446 (w10545, w10434, IN87[30], w10546, w10547);
  FullAdder U3447 (w10547, w10436, IN88[29], w10548, w10549);
  FullAdder U3448 (w10549, w10438, IN89[28], w10550, w10551);
  FullAdder U3449 (w10551, w10440, IN90[27], w10552, w10553);
  FullAdder U3450 (w10553, w10442, IN91[26], w10554, w10555);
  FullAdder U3451 (w10555, w10444, IN92[25], w10556, w10557);
  FullAdder U3452 (w10557, w10446, IN93[24], w10558, w10559);
  FullAdder U3453 (w10559, w10448, IN94[23], w10560, w10561);
  FullAdder U3454 (w10561, w10450, IN95[22], w10562, w10563);
  FullAdder U3455 (w10563, w10452, IN96[21], w10564, w10565);
  FullAdder U3456 (w10565, w10454, IN97[20], w10566, w10567);
  FullAdder U3457 (w10567, w10456, IN98[19], w10568, w10569);
  FullAdder U3458 (w10569, w10458, IN99[18], w10570, w10571);
  FullAdder U3459 (w10571, w10460, IN100[17], w10572, w10573);
  FullAdder U3460 (w10573, w10462, IN101[16], w10574, w10575);
  FullAdder U3461 (w10575, w10464, IN102[15], w10576, w10577);
  FullAdder U3462 (w10577, w10466, IN103[14], w10578, w10579);
  FullAdder U3463 (w10579, w10468, IN104[13], w10580, w10581);
  FullAdder U3464 (w10581, w10470, IN105[12], w10582, w10583);
  FullAdder U3465 (w10583, w10472, IN106[11], w10584, w10585);
  FullAdder U3466 (w10585, w10474, IN107[10], w10586, w10587);
  FullAdder U3467 (w10587, w10476, IN108[9], w10588, w10589);
  FullAdder U3468 (w10589, w10478, IN109[8], w10590, w10591);
  FullAdder U3469 (w10591, w10480, IN110[7], w10592, w10593);
  FullAdder U3470 (w10593, w10482, IN111[6], w10594, w10595);
  FullAdder U3471 (w10595, w10484, IN112[5], w10596, w10597);
  FullAdder U3472 (w10597, w10486, IN113[4], w10598, w10599);
  FullAdder U3473 (w10599, w10488, IN114[3], w10600, w10601);
  FullAdder U3474 (w10601, w10490, IN115[2], w10602, w10603);
  FullAdder U3475 (w10603, w10492, IN116[1], w10604, w10605);
  FullAdder U3476 (w10605, w10493, IN117[0], w10606, w10607);
  HalfAdder U3477 (w10496, IN62[56], Out1[62], w10609);
  FullAdder U3478 (w10609, w10498, IN63[55], Out1[63], w10611);
  FullAdder U3479 (w10611, w10500, IN64[54], Out1[64], w10613);
  FullAdder U3480 (w10613, w10502, IN65[53], Out1[65], w10615);
  FullAdder U3481 (w10615, w10504, IN66[52], Out1[66], w10617);
  FullAdder U3482 (w10617, w10506, IN67[51], Out1[67], w10619);
  FullAdder U3483 (w10619, w10508, IN68[50], Out1[68], w10621);
  FullAdder U3484 (w10621, w10510, IN69[49], Out1[69], w10623);
  FullAdder U3485 (w10623, w10512, IN70[48], Out1[70], w10625);
  FullAdder U3486 (w10625, w10514, IN71[47], Out1[71], w10627);
  FullAdder U3487 (w10627, w10516, IN72[46], Out1[72], w10629);
  FullAdder U3488 (w10629, w10518, IN73[45], Out1[73], w10631);
  FullAdder U3489 (w10631, w10520, IN74[44], Out1[74], w10633);
  FullAdder U3490 (w10633, w10522, IN75[43], Out1[75], w10635);
  FullAdder U3491 (w10635, w10524, IN76[42], Out1[76], w10637);
  FullAdder U3492 (w10637, w10526, IN77[41], Out1[77], w10639);
  FullAdder U3493 (w10639, w10528, IN78[40], Out1[78], w10641);
  FullAdder U3494 (w10641, w10530, IN79[39], Out1[79], w10643);
  FullAdder U3495 (w10643, w10532, IN80[38], Out1[80], w10645);
  FullAdder U3496 (w10645, w10534, IN81[37], Out1[81], w10647);
  FullAdder U3497 (w10647, w10536, IN82[36], Out1[82], w10649);
  FullAdder U3498 (w10649, w10538, IN83[35], Out1[83], w10651);
  FullAdder U3499 (w10651, w10540, IN84[34], Out1[84], w10653);
  FullAdder U3500 (w10653, w10542, IN85[33], Out1[85], w10655);
  FullAdder U3501 (w10655, w10544, IN86[32], Out1[86], w10657);
  FullAdder U3502 (w10657, w10546, IN87[31], Out1[87], w10659);
  FullAdder U3503 (w10659, w10548, IN88[30], Out1[88], w10661);
  FullAdder U3504 (w10661, w10550, IN89[29], Out1[89], w10663);
  FullAdder U3505 (w10663, w10552, IN90[28], Out1[90], w10665);
  FullAdder U3506 (w10665, w10554, IN91[27], Out1[91], w10667);
  FullAdder U3507 (w10667, w10556, IN92[26], Out1[92], w10669);
  FullAdder U3508 (w10669, w10558, IN93[25], Out1[93], w10671);
  FullAdder U3509 (w10671, w10560, IN94[24], Out1[94], w10673);
  FullAdder U3510 (w10673, w10562, IN95[23], Out1[95], w10675);
  FullAdder U3511 (w10675, w10564, IN96[22], Out1[96], w10677);
  FullAdder U3512 (w10677, w10566, IN97[21], Out1[97], w10679);
  FullAdder U3513 (w10679, w10568, IN98[20], Out1[98], w10681);
  FullAdder U3514 (w10681, w10570, IN99[19], Out1[99], w10683);
  FullAdder U3515 (w10683, w10572, IN100[18], Out1[100], w10685);
  FullAdder U3516 (w10685, w10574, IN101[17], Out1[101], w10687);
  FullAdder U3517 (w10687, w10576, IN102[16], Out1[102], w10689);
  FullAdder U3518 (w10689, w10578, IN103[15], Out1[103], w10691);
  FullAdder U3519 (w10691, w10580, IN104[14], Out1[104], w10693);
  FullAdder U3520 (w10693, w10582, IN105[13], Out1[105], w10695);
  FullAdder U3521 (w10695, w10584, IN106[12], Out1[106], w10697);
  FullAdder U3522 (w10697, w10586, IN107[11], Out1[107], w10699);
  FullAdder U3523 (w10699, w10588, IN108[10], Out1[108], w10701);
  FullAdder U3524 (w10701, w10590, IN109[9], Out1[109], w10703);
  FullAdder U3525 (w10703, w10592, IN110[8], Out1[110], w10705);
  FullAdder U3526 (w10705, w10594, IN111[7], Out1[111], w10707);
  FullAdder U3527 (w10707, w10596, IN112[6], Out1[112], w10709);
  FullAdder U3528 (w10709, w10598, IN113[5], Out1[113], w10711);
  FullAdder U3529 (w10711, w10600, IN114[4], Out1[114], w10713);
  FullAdder U3530 (w10713, w10602, IN115[3], Out1[115], w10715);
  FullAdder U3531 (w10715, w10604, IN116[2], Out1[116], w10717);
  FullAdder U3532 (w10717, w10606, IN117[1], Out1[117], w10719);
  FullAdder U3533 (w10719, w10607, IN118[0], Out1[118], Out1[119]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN58[57];
  assign Out2[1] = IN59[57];
  assign Out2[2] = IN60[57];
  assign Out2[3] = IN61[57];
  assign Out2[4] = IN62[57];
  assign Out2[5] = IN63[56];
  assign Out2[6] = IN64[55];
  assign Out2[7] = IN65[54];
  assign Out2[8] = IN66[53];
  assign Out2[9] = IN67[52];
  assign Out2[10] = IN68[51];
  assign Out2[11] = IN69[50];
  assign Out2[12] = IN70[49];
  assign Out2[13] = IN71[48];
  assign Out2[14] = IN72[47];
  assign Out2[15] = IN73[46];
  assign Out2[16] = IN74[45];
  assign Out2[17] = IN75[44];
  assign Out2[18] = IN76[43];
  assign Out2[19] = IN77[42];
  assign Out2[20] = IN78[41];
  assign Out2[21] = IN79[40];
  assign Out2[22] = IN80[39];
  assign Out2[23] = IN81[38];
  assign Out2[24] = IN82[37];
  assign Out2[25] = IN83[36];
  assign Out2[26] = IN84[35];
  assign Out2[27] = IN85[34];
  assign Out2[28] = IN86[33];
  assign Out2[29] = IN87[32];
  assign Out2[30] = IN88[31];
  assign Out2[31] = IN89[30];
  assign Out2[32] = IN90[29];
  assign Out2[33] = IN91[28];
  assign Out2[34] = IN92[27];
  assign Out2[35] = IN93[26];
  assign Out2[36] = IN94[25];
  assign Out2[37] = IN95[24];
  assign Out2[38] = IN96[23];
  assign Out2[39] = IN97[22];
  assign Out2[40] = IN98[21];
  assign Out2[41] = IN99[20];
  assign Out2[42] = IN100[19];
  assign Out2[43] = IN101[18];
  assign Out2[44] = IN102[17];
  assign Out2[45] = IN103[16];
  assign Out2[46] = IN104[15];
  assign Out2[47] = IN105[14];
  assign Out2[48] = IN106[13];
  assign Out2[49] = IN107[12];
  assign Out2[50] = IN108[11];
  assign Out2[51] = IN109[10];
  assign Out2[52] = IN110[9];
  assign Out2[53] = IN111[8];
  assign Out2[54] = IN112[7];
  assign Out2[55] = IN113[6];
  assign Out2[56] = IN114[5];
  assign Out2[57] = IN115[4];
  assign Out2[58] = IN116[3];
  assign Out2[59] = IN117[2];
  assign Out2[60] = IN118[1];
  assign Out2[61] = IN119[0];

endmodule
module RC_62_62(IN1, IN2, Out);
  input [61:0] IN1;
  input [61:0] IN2;
  output [62:0] Out;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  wire w211;
  wire w213;
  wire w215;
  wire w217;
  wire w219;
  wire w221;
  wire w223;
  wire w225;
  wire w227;
  wire w229;
  wire w231;
  wire w233;
  wire w235;
  wire w237;
  wire w239;
  wire w241;
  wire w243;
  wire w245;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w125);
  FullAdder U1 (IN1[1], IN2[1], w125, Out[1], w127);
  FullAdder U2 (IN1[2], IN2[2], w127, Out[2], w129);
  FullAdder U3 (IN1[3], IN2[3], w129, Out[3], w131);
  FullAdder U4 (IN1[4], IN2[4], w131, Out[4], w133);
  FullAdder U5 (IN1[5], IN2[5], w133, Out[5], w135);
  FullAdder U6 (IN1[6], IN2[6], w135, Out[6], w137);
  FullAdder U7 (IN1[7], IN2[7], w137, Out[7], w139);
  FullAdder U8 (IN1[8], IN2[8], w139, Out[8], w141);
  FullAdder U9 (IN1[9], IN2[9], w141, Out[9], w143);
  FullAdder U10 (IN1[10], IN2[10], w143, Out[10], w145);
  FullAdder U11 (IN1[11], IN2[11], w145, Out[11], w147);
  FullAdder U12 (IN1[12], IN2[12], w147, Out[12], w149);
  FullAdder U13 (IN1[13], IN2[13], w149, Out[13], w151);
  FullAdder U14 (IN1[14], IN2[14], w151, Out[14], w153);
  FullAdder U15 (IN1[15], IN2[15], w153, Out[15], w155);
  FullAdder U16 (IN1[16], IN2[16], w155, Out[16], w157);
  FullAdder U17 (IN1[17], IN2[17], w157, Out[17], w159);
  FullAdder U18 (IN1[18], IN2[18], w159, Out[18], w161);
  FullAdder U19 (IN1[19], IN2[19], w161, Out[19], w163);
  FullAdder U20 (IN1[20], IN2[20], w163, Out[20], w165);
  FullAdder U21 (IN1[21], IN2[21], w165, Out[21], w167);
  FullAdder U22 (IN1[22], IN2[22], w167, Out[22], w169);
  FullAdder U23 (IN1[23], IN2[23], w169, Out[23], w171);
  FullAdder U24 (IN1[24], IN2[24], w171, Out[24], w173);
  FullAdder U25 (IN1[25], IN2[25], w173, Out[25], w175);
  FullAdder U26 (IN1[26], IN2[26], w175, Out[26], w177);
  FullAdder U27 (IN1[27], IN2[27], w177, Out[27], w179);
  FullAdder U28 (IN1[28], IN2[28], w179, Out[28], w181);
  FullAdder U29 (IN1[29], IN2[29], w181, Out[29], w183);
  FullAdder U30 (IN1[30], IN2[30], w183, Out[30], w185);
  FullAdder U31 (IN1[31], IN2[31], w185, Out[31], w187);
  FullAdder U32 (IN1[32], IN2[32], w187, Out[32], w189);
  FullAdder U33 (IN1[33], IN2[33], w189, Out[33], w191);
  FullAdder U34 (IN1[34], IN2[34], w191, Out[34], w193);
  FullAdder U35 (IN1[35], IN2[35], w193, Out[35], w195);
  FullAdder U36 (IN1[36], IN2[36], w195, Out[36], w197);
  FullAdder U37 (IN1[37], IN2[37], w197, Out[37], w199);
  FullAdder U38 (IN1[38], IN2[38], w199, Out[38], w201);
  FullAdder U39 (IN1[39], IN2[39], w201, Out[39], w203);
  FullAdder U40 (IN1[40], IN2[40], w203, Out[40], w205);
  FullAdder U41 (IN1[41], IN2[41], w205, Out[41], w207);
  FullAdder U42 (IN1[42], IN2[42], w207, Out[42], w209);
  FullAdder U43 (IN1[43], IN2[43], w209, Out[43], w211);
  FullAdder U44 (IN1[44], IN2[44], w211, Out[44], w213);
  FullAdder U45 (IN1[45], IN2[45], w213, Out[45], w215);
  FullAdder U46 (IN1[46], IN2[46], w215, Out[46], w217);
  FullAdder U47 (IN1[47], IN2[47], w217, Out[47], w219);
  FullAdder U48 (IN1[48], IN2[48], w219, Out[48], w221);
  FullAdder U49 (IN1[49], IN2[49], w221, Out[49], w223);
  FullAdder U50 (IN1[50], IN2[50], w223, Out[50], w225);
  FullAdder U51 (IN1[51], IN2[51], w225, Out[51], w227);
  FullAdder U52 (IN1[52], IN2[52], w227, Out[52], w229);
  FullAdder U53 (IN1[53], IN2[53], w229, Out[53], w231);
  FullAdder U54 (IN1[54], IN2[54], w231, Out[54], w233);
  FullAdder U55 (IN1[55], IN2[55], w233, Out[55], w235);
  FullAdder U56 (IN1[56], IN2[56], w235, Out[56], w237);
  FullAdder U57 (IN1[57], IN2[57], w237, Out[57], w239);
  FullAdder U58 (IN1[58], IN2[58], w239, Out[58], w241);
  FullAdder U59 (IN1[59], IN2[59], w241, Out[59], w243);
  FullAdder U60 (IN1[60], IN2[60], w243, Out[60], w245);
  FullAdder U61 (IN1[61], IN2[61], w245, Out[61], Out[62]);

endmodule
module NR_58_63(IN1, IN2, Out);
  input [57:0] IN1;
  input [62:0] IN2;
  output [120:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [29:0] P29;
  wire [30:0] P30;
  wire [31:0] P31;
  wire [32:0] P32;
  wire [33:0] P33;
  wire [34:0] P34;
  wire [35:0] P35;
  wire [36:0] P36;
  wire [37:0] P37;
  wire [38:0] P38;
  wire [39:0] P39;
  wire [40:0] P40;
  wire [41:0] P41;
  wire [42:0] P42;
  wire [43:0] P43;
  wire [44:0] P44;
  wire [45:0] P45;
  wire [46:0] P46;
  wire [47:0] P47;
  wire [48:0] P48;
  wire [49:0] P49;
  wire [50:0] P50;
  wire [51:0] P51;
  wire [52:0] P52;
  wire [53:0] P53;
  wire [54:0] P54;
  wire [55:0] P55;
  wire [56:0] P56;
  wire [57:0] P57;
  wire [57:0] P58;
  wire [57:0] P59;
  wire [57:0] P60;
  wire [57:0] P61;
  wire [57:0] P62;
  wire [56:0] P63;
  wire [55:0] P64;
  wire [54:0] P65;
  wire [53:0] P66;
  wire [52:0] P67;
  wire [51:0] P68;
  wire [50:0] P69;
  wire [49:0] P70;
  wire [48:0] P71;
  wire [47:0] P72;
  wire [46:0] P73;
  wire [45:0] P74;
  wire [44:0] P75;
  wire [43:0] P76;
  wire [42:0] P77;
  wire [41:0] P78;
  wire [40:0] P79;
  wire [39:0] P80;
  wire [38:0] P81;
  wire [37:0] P82;
  wire [36:0] P83;
  wire [35:0] P84;
  wire [34:0] P85;
  wire [33:0] P86;
  wire [32:0] P87;
  wire [31:0] P88;
  wire [30:0] P89;
  wire [29:0] P90;
  wire [28:0] P91;
  wire [27:0] P92;
  wire [26:0] P93;
  wire [25:0] P94;
  wire [24:0] P95;
  wire [23:0] P96;
  wire [22:0] P97;
  wire [21:0] P98;
  wire [20:0] P99;
  wire [19:0] P100;
  wire [18:0] P101;
  wire [17:0] P102;
  wire [16:0] P103;
  wire [15:0] P104;
  wire [14:0] P105;
  wire [13:0] P106;
  wire [12:0] P107;
  wire [11:0] P108;
  wire [10:0] P109;
  wire [9:0] P110;
  wire [8:0] P111;
  wire [7:0] P112;
  wire [6:0] P113;
  wire [5:0] P114;
  wire [4:0] P115;
  wire [3:0] P116;
  wire [2:0] P117;
  wire [1:0] P118;
  wire [0:0] P119;
  wire [119:0] R1;
  wire [61:0] R2;
  wire [120:0] aOut;
  U_SP_58_63 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, P112, P113, P114, P115, P116, P117, P118, P119);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, P112, P113, P114, P115, P116, P117, P118, P119, R1, R2);
  RC_62_62 S2 (R1[119:58], R2, aOut[120:58]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign aOut[41] = R1[41];
  assign aOut[42] = R1[42];
  assign aOut[43] = R1[43];
  assign aOut[44] = R1[44];
  assign aOut[45] = R1[45];
  assign aOut[46] = R1[46];
  assign aOut[47] = R1[47];
  assign aOut[48] = R1[48];
  assign aOut[49] = R1[49];
  assign aOut[50] = R1[50];
  assign aOut[51] = R1[51];
  assign aOut[52] = R1[52];
  assign aOut[53] = R1[53];
  assign aOut[54] = R1[54];
  assign aOut[55] = R1[55];
  assign aOut[56] = R1[56];
  assign aOut[57] = R1[57];
  assign Out = aOut[120:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
