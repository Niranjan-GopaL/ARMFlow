
module customAdder56_0(
    input [55 : 0] A,
    input [55 : 0] B,
    output [56 : 0] Sum
);

    assign Sum = A+B;

endmodule
