//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 37
  second input length: 7
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_37_7(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42);
  input [36:0] IN1;
  input [6:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [6:0] P7;
  output [6:0] P8;
  output [6:0] P9;
  output [6:0] P10;
  output [6:0] P11;
  output [6:0] P12;
  output [6:0] P13;
  output [6:0] P14;
  output [6:0] P15;
  output [6:0] P16;
  output [6:0] P17;
  output [6:0] P18;
  output [6:0] P19;
  output [6:0] P20;
  output [6:0] P21;
  output [6:0] P22;
  output [6:0] P23;
  output [6:0] P24;
  output [6:0] P25;
  output [6:0] P26;
  output [6:0] P27;
  output [6:0] P28;
  output [6:0] P29;
  output [6:0] P30;
  output [6:0] P31;
  output [6:0] P32;
  output [6:0] P33;
  output [6:0] P34;
  output [6:0] P35;
  output [6:0] P36;
  output [5:0] P37;
  output [4:0] P38;
  output [3:0] P39;
  output [2:0] P40;
  output [1:0] P41;
  output [0:0] P42;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[0] = IN1[1]&IN2[6];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[1] = IN1[2]&IN2[5];
  assign P8[0] = IN1[2]&IN2[6];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[2] = IN1[3]&IN2[4];
  assign P8[1] = IN1[3]&IN2[5];
  assign P9[0] = IN1[3]&IN2[6];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[3] = IN1[4]&IN2[3];
  assign P8[2] = IN1[4]&IN2[4];
  assign P9[1] = IN1[4]&IN2[5];
  assign P10[0] = IN1[4]&IN2[6];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[4] = IN1[5]&IN2[2];
  assign P8[3] = IN1[5]&IN2[3];
  assign P9[2] = IN1[5]&IN2[4];
  assign P10[1] = IN1[5]&IN2[5];
  assign P11[0] = IN1[5]&IN2[6];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[5] = IN1[6]&IN2[1];
  assign P8[4] = IN1[6]&IN2[2];
  assign P9[3] = IN1[6]&IN2[3];
  assign P10[2] = IN1[6]&IN2[4];
  assign P11[1] = IN1[6]&IN2[5];
  assign P12[0] = IN1[6]&IN2[6];
  assign P7[6] = IN1[7]&IN2[0];
  assign P8[5] = IN1[7]&IN2[1];
  assign P9[4] = IN1[7]&IN2[2];
  assign P10[3] = IN1[7]&IN2[3];
  assign P11[2] = IN1[7]&IN2[4];
  assign P12[1] = IN1[7]&IN2[5];
  assign P13[0] = IN1[7]&IN2[6];
  assign P8[6] = IN1[8]&IN2[0];
  assign P9[5] = IN1[8]&IN2[1];
  assign P10[4] = IN1[8]&IN2[2];
  assign P11[3] = IN1[8]&IN2[3];
  assign P12[2] = IN1[8]&IN2[4];
  assign P13[1] = IN1[8]&IN2[5];
  assign P14[0] = IN1[8]&IN2[6];
  assign P9[6] = IN1[9]&IN2[0];
  assign P10[5] = IN1[9]&IN2[1];
  assign P11[4] = IN1[9]&IN2[2];
  assign P12[3] = IN1[9]&IN2[3];
  assign P13[2] = IN1[9]&IN2[4];
  assign P14[1] = IN1[9]&IN2[5];
  assign P15[0] = IN1[9]&IN2[6];
  assign P10[6] = IN1[10]&IN2[0];
  assign P11[5] = IN1[10]&IN2[1];
  assign P12[4] = IN1[10]&IN2[2];
  assign P13[3] = IN1[10]&IN2[3];
  assign P14[2] = IN1[10]&IN2[4];
  assign P15[1] = IN1[10]&IN2[5];
  assign P16[0] = IN1[10]&IN2[6];
  assign P11[6] = IN1[11]&IN2[0];
  assign P12[5] = IN1[11]&IN2[1];
  assign P13[4] = IN1[11]&IN2[2];
  assign P14[3] = IN1[11]&IN2[3];
  assign P15[2] = IN1[11]&IN2[4];
  assign P16[1] = IN1[11]&IN2[5];
  assign P17[0] = IN1[11]&IN2[6];
  assign P12[6] = IN1[12]&IN2[0];
  assign P13[5] = IN1[12]&IN2[1];
  assign P14[4] = IN1[12]&IN2[2];
  assign P15[3] = IN1[12]&IN2[3];
  assign P16[2] = IN1[12]&IN2[4];
  assign P17[1] = IN1[12]&IN2[5];
  assign P18[0] = IN1[12]&IN2[6];
  assign P13[6] = IN1[13]&IN2[0];
  assign P14[5] = IN1[13]&IN2[1];
  assign P15[4] = IN1[13]&IN2[2];
  assign P16[3] = IN1[13]&IN2[3];
  assign P17[2] = IN1[13]&IN2[4];
  assign P18[1] = IN1[13]&IN2[5];
  assign P19[0] = IN1[13]&IN2[6];
  assign P14[6] = IN1[14]&IN2[0];
  assign P15[5] = IN1[14]&IN2[1];
  assign P16[4] = IN1[14]&IN2[2];
  assign P17[3] = IN1[14]&IN2[3];
  assign P18[2] = IN1[14]&IN2[4];
  assign P19[1] = IN1[14]&IN2[5];
  assign P20[0] = IN1[14]&IN2[6];
  assign P15[6] = IN1[15]&IN2[0];
  assign P16[5] = IN1[15]&IN2[1];
  assign P17[4] = IN1[15]&IN2[2];
  assign P18[3] = IN1[15]&IN2[3];
  assign P19[2] = IN1[15]&IN2[4];
  assign P20[1] = IN1[15]&IN2[5];
  assign P21[0] = IN1[15]&IN2[6];
  assign P16[6] = IN1[16]&IN2[0];
  assign P17[5] = IN1[16]&IN2[1];
  assign P18[4] = IN1[16]&IN2[2];
  assign P19[3] = IN1[16]&IN2[3];
  assign P20[2] = IN1[16]&IN2[4];
  assign P21[1] = IN1[16]&IN2[5];
  assign P22[0] = IN1[16]&IN2[6];
  assign P17[6] = IN1[17]&IN2[0];
  assign P18[5] = IN1[17]&IN2[1];
  assign P19[4] = IN1[17]&IN2[2];
  assign P20[3] = IN1[17]&IN2[3];
  assign P21[2] = IN1[17]&IN2[4];
  assign P22[1] = IN1[17]&IN2[5];
  assign P23[0] = IN1[17]&IN2[6];
  assign P18[6] = IN1[18]&IN2[0];
  assign P19[5] = IN1[18]&IN2[1];
  assign P20[4] = IN1[18]&IN2[2];
  assign P21[3] = IN1[18]&IN2[3];
  assign P22[2] = IN1[18]&IN2[4];
  assign P23[1] = IN1[18]&IN2[5];
  assign P24[0] = IN1[18]&IN2[6];
  assign P19[6] = IN1[19]&IN2[0];
  assign P20[5] = IN1[19]&IN2[1];
  assign P21[4] = IN1[19]&IN2[2];
  assign P22[3] = IN1[19]&IN2[3];
  assign P23[2] = IN1[19]&IN2[4];
  assign P24[1] = IN1[19]&IN2[5];
  assign P25[0] = IN1[19]&IN2[6];
  assign P20[6] = IN1[20]&IN2[0];
  assign P21[5] = IN1[20]&IN2[1];
  assign P22[4] = IN1[20]&IN2[2];
  assign P23[3] = IN1[20]&IN2[3];
  assign P24[2] = IN1[20]&IN2[4];
  assign P25[1] = IN1[20]&IN2[5];
  assign P26[0] = IN1[20]&IN2[6];
  assign P21[6] = IN1[21]&IN2[0];
  assign P22[5] = IN1[21]&IN2[1];
  assign P23[4] = IN1[21]&IN2[2];
  assign P24[3] = IN1[21]&IN2[3];
  assign P25[2] = IN1[21]&IN2[4];
  assign P26[1] = IN1[21]&IN2[5];
  assign P27[0] = IN1[21]&IN2[6];
  assign P22[6] = IN1[22]&IN2[0];
  assign P23[5] = IN1[22]&IN2[1];
  assign P24[4] = IN1[22]&IN2[2];
  assign P25[3] = IN1[22]&IN2[3];
  assign P26[2] = IN1[22]&IN2[4];
  assign P27[1] = IN1[22]&IN2[5];
  assign P28[0] = IN1[22]&IN2[6];
  assign P23[6] = IN1[23]&IN2[0];
  assign P24[5] = IN1[23]&IN2[1];
  assign P25[4] = IN1[23]&IN2[2];
  assign P26[3] = IN1[23]&IN2[3];
  assign P27[2] = IN1[23]&IN2[4];
  assign P28[1] = IN1[23]&IN2[5];
  assign P29[0] = IN1[23]&IN2[6];
  assign P24[6] = IN1[24]&IN2[0];
  assign P25[5] = IN1[24]&IN2[1];
  assign P26[4] = IN1[24]&IN2[2];
  assign P27[3] = IN1[24]&IN2[3];
  assign P28[2] = IN1[24]&IN2[4];
  assign P29[1] = IN1[24]&IN2[5];
  assign P30[0] = IN1[24]&IN2[6];
  assign P25[6] = IN1[25]&IN2[0];
  assign P26[5] = IN1[25]&IN2[1];
  assign P27[4] = IN1[25]&IN2[2];
  assign P28[3] = IN1[25]&IN2[3];
  assign P29[2] = IN1[25]&IN2[4];
  assign P30[1] = IN1[25]&IN2[5];
  assign P31[0] = IN1[25]&IN2[6];
  assign P26[6] = IN1[26]&IN2[0];
  assign P27[5] = IN1[26]&IN2[1];
  assign P28[4] = IN1[26]&IN2[2];
  assign P29[3] = IN1[26]&IN2[3];
  assign P30[2] = IN1[26]&IN2[4];
  assign P31[1] = IN1[26]&IN2[5];
  assign P32[0] = IN1[26]&IN2[6];
  assign P27[6] = IN1[27]&IN2[0];
  assign P28[5] = IN1[27]&IN2[1];
  assign P29[4] = IN1[27]&IN2[2];
  assign P30[3] = IN1[27]&IN2[3];
  assign P31[2] = IN1[27]&IN2[4];
  assign P32[1] = IN1[27]&IN2[5];
  assign P33[0] = IN1[27]&IN2[6];
  assign P28[6] = IN1[28]&IN2[0];
  assign P29[5] = IN1[28]&IN2[1];
  assign P30[4] = IN1[28]&IN2[2];
  assign P31[3] = IN1[28]&IN2[3];
  assign P32[2] = IN1[28]&IN2[4];
  assign P33[1] = IN1[28]&IN2[5];
  assign P34[0] = IN1[28]&IN2[6];
  assign P29[6] = IN1[29]&IN2[0];
  assign P30[5] = IN1[29]&IN2[1];
  assign P31[4] = IN1[29]&IN2[2];
  assign P32[3] = IN1[29]&IN2[3];
  assign P33[2] = IN1[29]&IN2[4];
  assign P34[1] = IN1[29]&IN2[5];
  assign P35[0] = IN1[29]&IN2[6];
  assign P30[6] = IN1[30]&IN2[0];
  assign P31[5] = IN1[30]&IN2[1];
  assign P32[4] = IN1[30]&IN2[2];
  assign P33[3] = IN1[30]&IN2[3];
  assign P34[2] = IN1[30]&IN2[4];
  assign P35[1] = IN1[30]&IN2[5];
  assign P36[0] = IN1[30]&IN2[6];
  assign P31[6] = IN1[31]&IN2[0];
  assign P32[5] = IN1[31]&IN2[1];
  assign P33[4] = IN1[31]&IN2[2];
  assign P34[3] = IN1[31]&IN2[3];
  assign P35[2] = IN1[31]&IN2[4];
  assign P36[1] = IN1[31]&IN2[5];
  assign P37[0] = IN1[31]&IN2[6];
  assign P32[6] = IN1[32]&IN2[0];
  assign P33[5] = IN1[32]&IN2[1];
  assign P34[4] = IN1[32]&IN2[2];
  assign P35[3] = IN1[32]&IN2[3];
  assign P36[2] = IN1[32]&IN2[4];
  assign P37[1] = IN1[32]&IN2[5];
  assign P38[0] = IN1[32]&IN2[6];
  assign P33[6] = IN1[33]&IN2[0];
  assign P34[5] = IN1[33]&IN2[1];
  assign P35[4] = IN1[33]&IN2[2];
  assign P36[3] = IN1[33]&IN2[3];
  assign P37[2] = IN1[33]&IN2[4];
  assign P38[1] = IN1[33]&IN2[5];
  assign P39[0] = IN1[33]&IN2[6];
  assign P34[6] = IN1[34]&IN2[0];
  assign P35[5] = IN1[34]&IN2[1];
  assign P36[4] = IN1[34]&IN2[2];
  assign P37[3] = IN1[34]&IN2[3];
  assign P38[2] = IN1[34]&IN2[4];
  assign P39[1] = IN1[34]&IN2[5];
  assign P40[0] = IN1[34]&IN2[6];
  assign P35[6] = IN1[35]&IN2[0];
  assign P36[5] = IN1[35]&IN2[1];
  assign P37[4] = IN1[35]&IN2[2];
  assign P38[3] = IN1[35]&IN2[3];
  assign P39[2] = IN1[35]&IN2[4];
  assign P40[1] = IN1[35]&IN2[5];
  assign P41[0] = IN1[35]&IN2[6];
  assign P36[6] = IN1[36]&IN2[0];
  assign P37[5] = IN1[36]&IN2[1];
  assign P38[4] = IN1[36]&IN2[2];
  assign P39[3] = IN1[36]&IN2[3];
  assign P40[2] = IN1[36]&IN2[4];
  assign P41[1] = IN1[36]&IN2[5];
  assign P42[0] = IN1[36]&IN2[6];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [6:0] IN7;
  input [6:0] IN8;
  input [6:0] IN9;
  input [6:0] IN10;
  input [6:0] IN11;
  input [6:0] IN12;
  input [6:0] IN13;
  input [6:0] IN14;
  input [6:0] IN15;
  input [6:0] IN16;
  input [6:0] IN17;
  input [6:0] IN18;
  input [6:0] IN19;
  input [6:0] IN20;
  input [6:0] IN21;
  input [6:0] IN22;
  input [6:0] IN23;
  input [6:0] IN24;
  input [6:0] IN25;
  input [6:0] IN26;
  input [6:0] IN27;
  input [6:0] IN28;
  input [6:0] IN29;
  input [6:0] IN30;
  input [6:0] IN31;
  input [6:0] IN32;
  input [6:0] IN33;
  input [6:0] IN34;
  input [6:0] IN35;
  input [6:0] IN36;
  input [5:0] IN37;
  input [4:0] IN38;
  input [3:0] IN39;
  input [2:0] IN40;
  input [1:0] IN41;
  input [0:0] IN42;
  output [42:0] Out1;
  output [5:0] Out2;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w620;
  wire w622;
  wire w624;
  wire w626;
  wire w628;
  wire w630;
  wire w632;
  wire w634;
  wire w636;
  wire w638;
  wire w640;
  wire w642;
  wire w644;
  wire w646;
  wire w648;
  wire w650;
  wire w652;
  wire w654;
  wire w656;
  wire w658;
  wire w660;
  wire w662;
  wire w664;
  wire w666;
  wire w668;
  wire w670;
  wire w672;
  wire w674;
  wire w676;
  wire w678;
  wire w680;
  wire w682;
  wire w684;
  wire w686;
  wire w688;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w260);
  FullAdder U1 (w260, IN2[0], IN2[1], w261, w262);
  FullAdder U2 (w262, IN3[0], IN3[1], w263, w264);
  FullAdder U3 (w264, IN4[0], IN4[1], w265, w266);
  FullAdder U4 (w266, IN5[0], IN5[1], w267, w268);
  FullAdder U5 (w268, IN6[0], IN6[1], w269, w270);
  FullAdder U6 (w270, IN7[0], IN7[1], w271, w272);
  FullAdder U7 (w272, IN8[0], IN8[1], w273, w274);
  FullAdder U8 (w274, IN9[0], IN9[1], w275, w276);
  FullAdder U9 (w276, IN10[0], IN10[1], w277, w278);
  FullAdder U10 (w278, IN11[0], IN11[1], w279, w280);
  FullAdder U11 (w280, IN12[0], IN12[1], w281, w282);
  FullAdder U12 (w282, IN13[0], IN13[1], w283, w284);
  FullAdder U13 (w284, IN14[0], IN14[1], w285, w286);
  FullAdder U14 (w286, IN15[0], IN15[1], w287, w288);
  FullAdder U15 (w288, IN16[0], IN16[1], w289, w290);
  FullAdder U16 (w290, IN17[0], IN17[1], w291, w292);
  FullAdder U17 (w292, IN18[0], IN18[1], w293, w294);
  FullAdder U18 (w294, IN19[0], IN19[1], w295, w296);
  FullAdder U19 (w296, IN20[0], IN20[1], w297, w298);
  FullAdder U20 (w298, IN21[0], IN21[1], w299, w300);
  FullAdder U21 (w300, IN22[0], IN22[1], w301, w302);
  FullAdder U22 (w302, IN23[0], IN23[1], w303, w304);
  FullAdder U23 (w304, IN24[0], IN24[1], w305, w306);
  FullAdder U24 (w306, IN25[0], IN25[1], w307, w308);
  FullAdder U25 (w308, IN26[0], IN26[1], w309, w310);
  FullAdder U26 (w310, IN27[0], IN27[1], w311, w312);
  FullAdder U27 (w312, IN28[0], IN28[1], w313, w314);
  FullAdder U28 (w314, IN29[0], IN29[1], w315, w316);
  FullAdder U29 (w316, IN30[0], IN30[1], w317, w318);
  FullAdder U30 (w318, IN31[0], IN31[1], w319, w320);
  FullAdder U31 (w320, IN32[0], IN32[1], w321, w322);
  FullAdder U32 (w322, IN33[0], IN33[1], w323, w324);
  FullAdder U33 (w324, IN34[0], IN34[1], w325, w326);
  FullAdder U34 (w326, IN35[0], IN35[1], w327, w328);
  FullAdder U35 (w328, IN36[0], IN36[1], w329, w330);
  HalfAdder U36 (w261, IN2[2], Out1[2], w332);
  FullAdder U37 (w332, w263, IN3[2], w333, w334);
  FullAdder U38 (w334, w265, IN4[2], w335, w336);
  FullAdder U39 (w336, w267, IN5[2], w337, w338);
  FullAdder U40 (w338, w269, IN6[2], w339, w340);
  FullAdder U41 (w340, w271, IN7[2], w341, w342);
  FullAdder U42 (w342, w273, IN8[2], w343, w344);
  FullAdder U43 (w344, w275, IN9[2], w345, w346);
  FullAdder U44 (w346, w277, IN10[2], w347, w348);
  FullAdder U45 (w348, w279, IN11[2], w349, w350);
  FullAdder U46 (w350, w281, IN12[2], w351, w352);
  FullAdder U47 (w352, w283, IN13[2], w353, w354);
  FullAdder U48 (w354, w285, IN14[2], w355, w356);
  FullAdder U49 (w356, w287, IN15[2], w357, w358);
  FullAdder U50 (w358, w289, IN16[2], w359, w360);
  FullAdder U51 (w360, w291, IN17[2], w361, w362);
  FullAdder U52 (w362, w293, IN18[2], w363, w364);
  FullAdder U53 (w364, w295, IN19[2], w365, w366);
  FullAdder U54 (w366, w297, IN20[2], w367, w368);
  FullAdder U55 (w368, w299, IN21[2], w369, w370);
  FullAdder U56 (w370, w301, IN22[2], w371, w372);
  FullAdder U57 (w372, w303, IN23[2], w373, w374);
  FullAdder U58 (w374, w305, IN24[2], w375, w376);
  FullAdder U59 (w376, w307, IN25[2], w377, w378);
  FullAdder U60 (w378, w309, IN26[2], w379, w380);
  FullAdder U61 (w380, w311, IN27[2], w381, w382);
  FullAdder U62 (w382, w313, IN28[2], w383, w384);
  FullAdder U63 (w384, w315, IN29[2], w385, w386);
  FullAdder U64 (w386, w317, IN30[2], w387, w388);
  FullAdder U65 (w388, w319, IN31[2], w389, w390);
  FullAdder U66 (w390, w321, IN32[2], w391, w392);
  FullAdder U67 (w392, w323, IN33[2], w393, w394);
  FullAdder U68 (w394, w325, IN34[2], w395, w396);
  FullAdder U69 (w396, w327, IN35[2], w397, w398);
  FullAdder U70 (w398, w329, IN36[2], w399, w400);
  FullAdder U71 (w400, w330, IN37[0], w401, w402);
  HalfAdder U72 (w333, IN3[3], Out1[3], w404);
  FullAdder U73 (w404, w335, IN4[3], w405, w406);
  FullAdder U74 (w406, w337, IN5[3], w407, w408);
  FullAdder U75 (w408, w339, IN6[3], w409, w410);
  FullAdder U76 (w410, w341, IN7[3], w411, w412);
  FullAdder U77 (w412, w343, IN8[3], w413, w414);
  FullAdder U78 (w414, w345, IN9[3], w415, w416);
  FullAdder U79 (w416, w347, IN10[3], w417, w418);
  FullAdder U80 (w418, w349, IN11[3], w419, w420);
  FullAdder U81 (w420, w351, IN12[3], w421, w422);
  FullAdder U82 (w422, w353, IN13[3], w423, w424);
  FullAdder U83 (w424, w355, IN14[3], w425, w426);
  FullAdder U84 (w426, w357, IN15[3], w427, w428);
  FullAdder U85 (w428, w359, IN16[3], w429, w430);
  FullAdder U86 (w430, w361, IN17[3], w431, w432);
  FullAdder U87 (w432, w363, IN18[3], w433, w434);
  FullAdder U88 (w434, w365, IN19[3], w435, w436);
  FullAdder U89 (w436, w367, IN20[3], w437, w438);
  FullAdder U90 (w438, w369, IN21[3], w439, w440);
  FullAdder U91 (w440, w371, IN22[3], w441, w442);
  FullAdder U92 (w442, w373, IN23[3], w443, w444);
  FullAdder U93 (w444, w375, IN24[3], w445, w446);
  FullAdder U94 (w446, w377, IN25[3], w447, w448);
  FullAdder U95 (w448, w379, IN26[3], w449, w450);
  FullAdder U96 (w450, w381, IN27[3], w451, w452);
  FullAdder U97 (w452, w383, IN28[3], w453, w454);
  FullAdder U98 (w454, w385, IN29[3], w455, w456);
  FullAdder U99 (w456, w387, IN30[3], w457, w458);
  FullAdder U100 (w458, w389, IN31[3], w459, w460);
  FullAdder U101 (w460, w391, IN32[3], w461, w462);
  FullAdder U102 (w462, w393, IN33[3], w463, w464);
  FullAdder U103 (w464, w395, IN34[3], w465, w466);
  FullAdder U104 (w466, w397, IN35[3], w467, w468);
  FullAdder U105 (w468, w399, IN36[3], w469, w470);
  FullAdder U106 (w470, w401, IN37[1], w471, w472);
  FullAdder U107 (w472, w402, IN38[0], w473, w474);
  HalfAdder U108 (w405, IN4[4], Out1[4], w476);
  FullAdder U109 (w476, w407, IN5[4], w477, w478);
  FullAdder U110 (w478, w409, IN6[4], w479, w480);
  FullAdder U111 (w480, w411, IN7[4], w481, w482);
  FullAdder U112 (w482, w413, IN8[4], w483, w484);
  FullAdder U113 (w484, w415, IN9[4], w485, w486);
  FullAdder U114 (w486, w417, IN10[4], w487, w488);
  FullAdder U115 (w488, w419, IN11[4], w489, w490);
  FullAdder U116 (w490, w421, IN12[4], w491, w492);
  FullAdder U117 (w492, w423, IN13[4], w493, w494);
  FullAdder U118 (w494, w425, IN14[4], w495, w496);
  FullAdder U119 (w496, w427, IN15[4], w497, w498);
  FullAdder U120 (w498, w429, IN16[4], w499, w500);
  FullAdder U121 (w500, w431, IN17[4], w501, w502);
  FullAdder U122 (w502, w433, IN18[4], w503, w504);
  FullAdder U123 (w504, w435, IN19[4], w505, w506);
  FullAdder U124 (w506, w437, IN20[4], w507, w508);
  FullAdder U125 (w508, w439, IN21[4], w509, w510);
  FullAdder U126 (w510, w441, IN22[4], w511, w512);
  FullAdder U127 (w512, w443, IN23[4], w513, w514);
  FullAdder U128 (w514, w445, IN24[4], w515, w516);
  FullAdder U129 (w516, w447, IN25[4], w517, w518);
  FullAdder U130 (w518, w449, IN26[4], w519, w520);
  FullAdder U131 (w520, w451, IN27[4], w521, w522);
  FullAdder U132 (w522, w453, IN28[4], w523, w524);
  FullAdder U133 (w524, w455, IN29[4], w525, w526);
  FullAdder U134 (w526, w457, IN30[4], w527, w528);
  FullAdder U135 (w528, w459, IN31[4], w529, w530);
  FullAdder U136 (w530, w461, IN32[4], w531, w532);
  FullAdder U137 (w532, w463, IN33[4], w533, w534);
  FullAdder U138 (w534, w465, IN34[4], w535, w536);
  FullAdder U139 (w536, w467, IN35[4], w537, w538);
  FullAdder U140 (w538, w469, IN36[4], w539, w540);
  FullAdder U141 (w540, w471, IN37[2], w541, w542);
  FullAdder U142 (w542, w473, IN38[1], w543, w544);
  FullAdder U143 (w544, w474, IN39[0], w545, w546);
  HalfAdder U144 (w477, IN5[5], Out1[5], w548);
  FullAdder U145 (w548, w479, IN6[5], w549, w550);
  FullAdder U146 (w550, w481, IN7[5], w551, w552);
  FullAdder U147 (w552, w483, IN8[5], w553, w554);
  FullAdder U148 (w554, w485, IN9[5], w555, w556);
  FullAdder U149 (w556, w487, IN10[5], w557, w558);
  FullAdder U150 (w558, w489, IN11[5], w559, w560);
  FullAdder U151 (w560, w491, IN12[5], w561, w562);
  FullAdder U152 (w562, w493, IN13[5], w563, w564);
  FullAdder U153 (w564, w495, IN14[5], w565, w566);
  FullAdder U154 (w566, w497, IN15[5], w567, w568);
  FullAdder U155 (w568, w499, IN16[5], w569, w570);
  FullAdder U156 (w570, w501, IN17[5], w571, w572);
  FullAdder U157 (w572, w503, IN18[5], w573, w574);
  FullAdder U158 (w574, w505, IN19[5], w575, w576);
  FullAdder U159 (w576, w507, IN20[5], w577, w578);
  FullAdder U160 (w578, w509, IN21[5], w579, w580);
  FullAdder U161 (w580, w511, IN22[5], w581, w582);
  FullAdder U162 (w582, w513, IN23[5], w583, w584);
  FullAdder U163 (w584, w515, IN24[5], w585, w586);
  FullAdder U164 (w586, w517, IN25[5], w587, w588);
  FullAdder U165 (w588, w519, IN26[5], w589, w590);
  FullAdder U166 (w590, w521, IN27[5], w591, w592);
  FullAdder U167 (w592, w523, IN28[5], w593, w594);
  FullAdder U168 (w594, w525, IN29[5], w595, w596);
  FullAdder U169 (w596, w527, IN30[5], w597, w598);
  FullAdder U170 (w598, w529, IN31[5], w599, w600);
  FullAdder U171 (w600, w531, IN32[5], w601, w602);
  FullAdder U172 (w602, w533, IN33[5], w603, w604);
  FullAdder U173 (w604, w535, IN34[5], w605, w606);
  FullAdder U174 (w606, w537, IN35[5], w607, w608);
  FullAdder U175 (w608, w539, IN36[5], w609, w610);
  FullAdder U176 (w610, w541, IN37[3], w611, w612);
  FullAdder U177 (w612, w543, IN38[2], w613, w614);
  FullAdder U178 (w614, w545, IN39[1], w615, w616);
  FullAdder U179 (w616, w546, IN40[0], w617, w618);
  HalfAdder U180 (w549, IN6[6], Out1[6], w620);
  FullAdder U181 (w620, w551, IN7[6], Out1[7], w622);
  FullAdder U182 (w622, w553, IN8[6], Out1[8], w624);
  FullAdder U183 (w624, w555, IN9[6], Out1[9], w626);
  FullAdder U184 (w626, w557, IN10[6], Out1[10], w628);
  FullAdder U185 (w628, w559, IN11[6], Out1[11], w630);
  FullAdder U186 (w630, w561, IN12[6], Out1[12], w632);
  FullAdder U187 (w632, w563, IN13[6], Out1[13], w634);
  FullAdder U188 (w634, w565, IN14[6], Out1[14], w636);
  FullAdder U189 (w636, w567, IN15[6], Out1[15], w638);
  FullAdder U190 (w638, w569, IN16[6], Out1[16], w640);
  FullAdder U191 (w640, w571, IN17[6], Out1[17], w642);
  FullAdder U192 (w642, w573, IN18[6], Out1[18], w644);
  FullAdder U193 (w644, w575, IN19[6], Out1[19], w646);
  FullAdder U194 (w646, w577, IN20[6], Out1[20], w648);
  FullAdder U195 (w648, w579, IN21[6], Out1[21], w650);
  FullAdder U196 (w650, w581, IN22[6], Out1[22], w652);
  FullAdder U197 (w652, w583, IN23[6], Out1[23], w654);
  FullAdder U198 (w654, w585, IN24[6], Out1[24], w656);
  FullAdder U199 (w656, w587, IN25[6], Out1[25], w658);
  FullAdder U200 (w658, w589, IN26[6], Out1[26], w660);
  FullAdder U201 (w660, w591, IN27[6], Out1[27], w662);
  FullAdder U202 (w662, w593, IN28[6], Out1[28], w664);
  FullAdder U203 (w664, w595, IN29[6], Out1[29], w666);
  FullAdder U204 (w666, w597, IN30[6], Out1[30], w668);
  FullAdder U205 (w668, w599, IN31[6], Out1[31], w670);
  FullAdder U206 (w670, w601, IN32[6], Out1[32], w672);
  FullAdder U207 (w672, w603, IN33[6], Out1[33], w674);
  FullAdder U208 (w674, w605, IN34[6], Out1[34], w676);
  FullAdder U209 (w676, w607, IN35[6], Out1[35], w678);
  FullAdder U210 (w678, w609, IN36[6], Out1[36], w680);
  FullAdder U211 (w680, w611, IN37[4], Out1[37], w682);
  FullAdder U212 (w682, w613, IN38[3], Out1[38], w684);
  FullAdder U213 (w684, w615, IN39[2], Out1[39], w686);
  FullAdder U214 (w686, w617, IN40[1], Out1[40], w688);
  FullAdder U215 (w688, w618, IN41[0], Out1[41], Out1[42]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN37[5];
  assign Out2[1] = IN38[4];
  assign Out2[2] = IN39[3];
  assign Out2[3] = IN40[2];
  assign Out2[4] = IN41[1];
  assign Out2[5] = IN42[0];

endmodule
module RC_6_6(IN1, IN2, Out);
  input [5:0] IN1;
  input [5:0] IN2;
  output [6:0] Out;
  wire w13;
  wire w15;
  wire w17;
  wire w19;
  wire w21;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w13);
  FullAdder U1 (IN1[1], IN2[1], w13, Out[1], w15);
  FullAdder U2 (IN1[2], IN2[2], w15, Out[2], w17);
  FullAdder U3 (IN1[3], IN2[3], w17, Out[3], w19);
  FullAdder U4 (IN1[4], IN2[4], w19, Out[4], w21);
  FullAdder U5 (IN1[5], IN2[5], w21, Out[5], Out[6]);

endmodule
module NR_37_7(IN1, IN2, Out);
  input [36:0] IN1;
  input [6:0] IN2;
  output [43:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [6:0] P7;
  wire [6:0] P8;
  wire [6:0] P9;
  wire [6:0] P10;
  wire [6:0] P11;
  wire [6:0] P12;
  wire [6:0] P13;
  wire [6:0] P14;
  wire [6:0] P15;
  wire [6:0] P16;
  wire [6:0] P17;
  wire [6:0] P18;
  wire [6:0] P19;
  wire [6:0] P20;
  wire [6:0] P21;
  wire [6:0] P22;
  wire [6:0] P23;
  wire [6:0] P24;
  wire [6:0] P25;
  wire [6:0] P26;
  wire [6:0] P27;
  wire [6:0] P28;
  wire [6:0] P29;
  wire [6:0] P30;
  wire [6:0] P31;
  wire [6:0] P32;
  wire [6:0] P33;
  wire [6:0] P34;
  wire [6:0] P35;
  wire [6:0] P36;
  wire [5:0] P37;
  wire [4:0] P38;
  wire [3:0] P39;
  wire [2:0] P40;
  wire [1:0] P41;
  wire [0:0] P42;
  wire [42:0] R1;
  wire [5:0] R2;
  wire [43:0] aOut;
  U_SP_37_7 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, R1, R2);
  RC_6_6 S2 (R1[42:37], R2, aOut[43:37]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign Out = aOut[43:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
