//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 11
  second input length: 33
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_11_33(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42);
  input [10:0] IN1;
  input [32:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [10:0] P11;
  output [10:0] P12;
  output [10:0] P13;
  output [10:0] P14;
  output [10:0] P15;
  output [10:0] P16;
  output [10:0] P17;
  output [10:0] P18;
  output [10:0] P19;
  output [10:0] P20;
  output [10:0] P21;
  output [10:0] P22;
  output [10:0] P23;
  output [10:0] P24;
  output [10:0] P25;
  output [10:0] P26;
  output [10:0] P27;
  output [10:0] P28;
  output [10:0] P29;
  output [10:0] P30;
  output [10:0] P31;
  output [10:0] P32;
  output [9:0] P33;
  output [8:0] P34;
  output [7:0] P35;
  output [6:0] P36;
  output [5:0] P37;
  output [4:0] P38;
  output [3:0] P39;
  output [2:0] P40;
  output [1:0] P41;
  output [0:0] P42;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[0] = IN1[1]&IN2[32];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[1] = IN1[2]&IN2[31];
  assign P34[0] = IN1[2]&IN2[32];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[2] = IN1[3]&IN2[30];
  assign P34[1] = IN1[3]&IN2[31];
  assign P35[0] = IN1[3]&IN2[32];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[3] = IN1[4]&IN2[29];
  assign P34[2] = IN1[4]&IN2[30];
  assign P35[1] = IN1[4]&IN2[31];
  assign P36[0] = IN1[4]&IN2[32];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[4] = IN1[5]&IN2[28];
  assign P34[3] = IN1[5]&IN2[29];
  assign P35[2] = IN1[5]&IN2[30];
  assign P36[1] = IN1[5]&IN2[31];
  assign P37[0] = IN1[5]&IN2[32];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[5] = IN1[6]&IN2[27];
  assign P34[4] = IN1[6]&IN2[28];
  assign P35[3] = IN1[6]&IN2[29];
  assign P36[2] = IN1[6]&IN2[30];
  assign P37[1] = IN1[6]&IN2[31];
  assign P38[0] = IN1[6]&IN2[32];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[6] = IN1[7]&IN2[26];
  assign P34[5] = IN1[7]&IN2[27];
  assign P35[4] = IN1[7]&IN2[28];
  assign P36[3] = IN1[7]&IN2[29];
  assign P37[2] = IN1[7]&IN2[30];
  assign P38[1] = IN1[7]&IN2[31];
  assign P39[0] = IN1[7]&IN2[32];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[7] = IN1[8]&IN2[25];
  assign P34[6] = IN1[8]&IN2[26];
  assign P35[5] = IN1[8]&IN2[27];
  assign P36[4] = IN1[8]&IN2[28];
  assign P37[3] = IN1[8]&IN2[29];
  assign P38[2] = IN1[8]&IN2[30];
  assign P39[1] = IN1[8]&IN2[31];
  assign P40[0] = IN1[8]&IN2[32];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[8] = IN1[9]&IN2[24];
  assign P34[7] = IN1[9]&IN2[25];
  assign P35[6] = IN1[9]&IN2[26];
  assign P36[5] = IN1[9]&IN2[27];
  assign P37[4] = IN1[9]&IN2[28];
  assign P38[3] = IN1[9]&IN2[29];
  assign P39[2] = IN1[9]&IN2[30];
  assign P40[1] = IN1[9]&IN2[31];
  assign P41[0] = IN1[9]&IN2[32];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[9] = IN1[10]&IN2[23];
  assign P34[8] = IN1[10]&IN2[24];
  assign P35[7] = IN1[10]&IN2[25];
  assign P36[6] = IN1[10]&IN2[26];
  assign P37[5] = IN1[10]&IN2[27];
  assign P38[4] = IN1[10]&IN2[28];
  assign P39[3] = IN1[10]&IN2[29];
  assign P40[2] = IN1[10]&IN2[30];
  assign P41[1] = IN1[10]&IN2[31];
  assign P42[0] = IN1[10]&IN2[32];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [10:0] IN11;
  input [10:0] IN12;
  input [10:0] IN13;
  input [10:0] IN14;
  input [10:0] IN15;
  input [10:0] IN16;
  input [10:0] IN17;
  input [10:0] IN18;
  input [10:0] IN19;
  input [10:0] IN20;
  input [10:0] IN21;
  input [10:0] IN22;
  input [10:0] IN23;
  input [10:0] IN24;
  input [10:0] IN25;
  input [10:0] IN26;
  input [10:0] IN27;
  input [10:0] IN28;
  input [10:0] IN29;
  input [10:0] IN30;
  input [10:0] IN31;
  input [10:0] IN32;
  input [9:0] IN33;
  input [8:0] IN34;
  input [7:0] IN35;
  input [6:0] IN36;
  input [5:0] IN37;
  input [4:0] IN38;
  input [3:0] IN39;
  input [2:0] IN40;
  input [1:0] IN41;
  input [0:0] IN42;
  output [42:0] Out1;
  output [31:0] Out2;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w621;
  wire w622;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w669;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w717;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w764;
  wire w765;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w813;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w861;
  wire w862;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w909;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w933;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w957;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w981;
  wire w982;
  wire w984;
  wire w986;
  wire w988;
  wire w990;
  wire w992;
  wire w994;
  wire w996;
  wire w998;
  wire w1000;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w364);
  FullAdder U1 (w364, IN2[0], IN2[1], w365, w366);
  FullAdder U2 (w366, IN3[0], IN3[1], w367, w368);
  FullAdder U3 (w368, IN4[0], IN4[1], w369, w370);
  FullAdder U4 (w370, IN5[0], IN5[1], w371, w372);
  FullAdder U5 (w372, IN6[0], IN6[1], w373, w374);
  FullAdder U6 (w374, IN7[0], IN7[1], w375, w376);
  FullAdder U7 (w376, IN8[0], IN8[1], w377, w378);
  FullAdder U8 (w378, IN9[0], IN9[1], w379, w380);
  FullAdder U9 (w380, IN10[0], IN10[1], w381, w382);
  HalfAdder U10 (w365, IN2[2], Out1[2], w384);
  FullAdder U11 (w384, w367, IN3[2], w385, w386);
  FullAdder U12 (w386, w369, IN4[2], w387, w388);
  FullAdder U13 (w388, w371, IN5[2], w389, w390);
  FullAdder U14 (w390, w373, IN6[2], w391, w392);
  FullAdder U15 (w392, w375, IN7[2], w393, w394);
  FullAdder U16 (w394, w377, IN8[2], w395, w396);
  FullAdder U17 (w396, w379, IN9[2], w397, w398);
  FullAdder U18 (w398, w381, IN10[2], w399, w400);
  FullAdder U19 (w400, w382, IN11[0], w401, w402);
  HalfAdder U20 (w385, IN3[3], Out1[3], w404);
  FullAdder U21 (w404, w387, IN4[3], w405, w406);
  FullAdder U22 (w406, w389, IN5[3], w407, w408);
  FullAdder U23 (w408, w391, IN6[3], w409, w410);
  FullAdder U24 (w410, w393, IN7[3], w411, w412);
  FullAdder U25 (w412, w395, IN8[3], w413, w414);
  FullAdder U26 (w414, w397, IN9[3], w415, w416);
  FullAdder U27 (w416, w399, IN10[3], w417, w418);
  FullAdder U28 (w418, w401, IN11[1], w419, w420);
  FullAdder U29 (w420, w402, IN12[0], w421, w422);
  HalfAdder U30 (w405, IN4[4], Out1[4], w424);
  FullAdder U31 (w424, w407, IN5[4], w425, w426);
  FullAdder U32 (w426, w409, IN6[4], w427, w428);
  FullAdder U33 (w428, w411, IN7[4], w429, w430);
  FullAdder U34 (w430, w413, IN8[4], w431, w432);
  FullAdder U35 (w432, w415, IN9[4], w433, w434);
  FullAdder U36 (w434, w417, IN10[4], w435, w436);
  FullAdder U37 (w436, w419, IN11[2], w437, w438);
  FullAdder U38 (w438, w421, IN12[1], w439, w440);
  FullAdder U39 (w440, w422, IN13[0], w441, w442);
  HalfAdder U40 (w425, IN5[5], Out1[5], w444);
  FullAdder U41 (w444, w427, IN6[5], w445, w446);
  FullAdder U42 (w446, w429, IN7[5], w447, w448);
  FullAdder U43 (w448, w431, IN8[5], w449, w450);
  FullAdder U44 (w450, w433, IN9[5], w451, w452);
  FullAdder U45 (w452, w435, IN10[5], w453, w454);
  FullAdder U46 (w454, w437, IN11[3], w455, w456);
  FullAdder U47 (w456, w439, IN12[2], w457, w458);
  FullAdder U48 (w458, w441, IN13[1], w459, w460);
  FullAdder U49 (w460, w442, IN14[0], w461, w462);
  HalfAdder U50 (w445, IN6[6], Out1[6], w464);
  FullAdder U51 (w464, w447, IN7[6], w465, w466);
  FullAdder U52 (w466, w449, IN8[6], w467, w468);
  FullAdder U53 (w468, w451, IN9[6], w469, w470);
  FullAdder U54 (w470, w453, IN10[6], w471, w472);
  FullAdder U55 (w472, w455, IN11[4], w473, w474);
  FullAdder U56 (w474, w457, IN12[3], w475, w476);
  FullAdder U57 (w476, w459, IN13[2], w477, w478);
  FullAdder U58 (w478, w461, IN14[1], w479, w480);
  FullAdder U59 (w480, w462, IN15[0], w481, w482);
  HalfAdder U60 (w465, IN7[7], Out1[7], w484);
  FullAdder U61 (w484, w467, IN8[7], w485, w486);
  FullAdder U62 (w486, w469, IN9[7], w487, w488);
  FullAdder U63 (w488, w471, IN10[7], w489, w490);
  FullAdder U64 (w490, w473, IN11[5], w491, w492);
  FullAdder U65 (w492, w475, IN12[4], w493, w494);
  FullAdder U66 (w494, w477, IN13[3], w495, w496);
  FullAdder U67 (w496, w479, IN14[2], w497, w498);
  FullAdder U68 (w498, w481, IN15[1], w499, w500);
  FullAdder U69 (w500, w482, IN16[0], w501, w502);
  HalfAdder U70 (w485, IN8[8], Out1[8], w504);
  FullAdder U71 (w504, w487, IN9[8], w505, w506);
  FullAdder U72 (w506, w489, IN10[8], w507, w508);
  FullAdder U73 (w508, w491, IN11[6], w509, w510);
  FullAdder U74 (w510, w493, IN12[5], w511, w512);
  FullAdder U75 (w512, w495, IN13[4], w513, w514);
  FullAdder U76 (w514, w497, IN14[3], w515, w516);
  FullAdder U77 (w516, w499, IN15[2], w517, w518);
  FullAdder U78 (w518, w501, IN16[1], w519, w520);
  FullAdder U79 (w520, w502, IN17[0], w521, w522);
  HalfAdder U80 (w505, IN9[9], Out1[9], w524);
  FullAdder U81 (w524, w507, IN10[9], w525, w526);
  FullAdder U82 (w526, w509, IN11[7], w527, w528);
  FullAdder U83 (w528, w511, IN12[6], w529, w530);
  FullAdder U84 (w530, w513, IN13[5], w531, w532);
  FullAdder U85 (w532, w515, IN14[4], w533, w534);
  FullAdder U86 (w534, w517, IN15[3], w535, w536);
  FullAdder U87 (w536, w519, IN16[2], w537, w538);
  FullAdder U88 (w538, w521, IN17[1], w539, w540);
  FullAdder U89 (w540, w522, IN18[0], w541, w542);
  HalfAdder U90 (w525, IN10[10], Out1[10], w544);
  FullAdder U91 (w544, w527, IN11[8], w545, w546);
  FullAdder U92 (w546, w529, IN12[7], w547, w548);
  FullAdder U93 (w548, w531, IN13[6], w549, w550);
  FullAdder U94 (w550, w533, IN14[5], w551, w552);
  FullAdder U95 (w552, w535, IN15[4], w553, w554);
  FullAdder U96 (w554, w537, IN16[3], w555, w556);
  FullAdder U97 (w556, w539, IN17[2], w557, w558);
  FullAdder U98 (w558, w541, IN18[1], w559, w560);
  FullAdder U99 (w560, w542, IN19[0], w561, w562);
  HalfAdder U100 (w545, IN11[9], Out1[11], w564);
  FullAdder U101 (w564, w547, IN12[8], w565, w566);
  FullAdder U102 (w566, w549, IN13[7], w567, w568);
  FullAdder U103 (w568, w551, IN14[6], w569, w570);
  FullAdder U104 (w570, w553, IN15[5], w571, w572);
  FullAdder U105 (w572, w555, IN16[4], w573, w574);
  FullAdder U106 (w574, w557, IN17[3], w575, w576);
  FullAdder U107 (w576, w559, IN18[2], w577, w578);
  FullAdder U108 (w578, w561, IN19[1], w579, w580);
  FullAdder U109 (w580, w562, IN20[0], w581, w582);
  HalfAdder U110 (w565, IN12[9], Out1[12], w584);
  FullAdder U111 (w584, w567, IN13[8], w585, w586);
  FullAdder U112 (w586, w569, IN14[7], w587, w588);
  FullAdder U113 (w588, w571, IN15[6], w589, w590);
  FullAdder U114 (w590, w573, IN16[5], w591, w592);
  FullAdder U115 (w592, w575, IN17[4], w593, w594);
  FullAdder U116 (w594, w577, IN18[3], w595, w596);
  FullAdder U117 (w596, w579, IN19[2], w597, w598);
  FullAdder U118 (w598, w581, IN20[1], w599, w600);
  FullAdder U119 (w600, w582, IN21[0], w601, w602);
  HalfAdder U120 (w585, IN13[9], Out1[13], w604);
  FullAdder U121 (w604, w587, IN14[8], w605, w606);
  FullAdder U122 (w606, w589, IN15[7], w607, w608);
  FullAdder U123 (w608, w591, IN16[6], w609, w610);
  FullAdder U124 (w610, w593, IN17[5], w611, w612);
  FullAdder U125 (w612, w595, IN18[4], w613, w614);
  FullAdder U126 (w614, w597, IN19[3], w615, w616);
  FullAdder U127 (w616, w599, IN20[2], w617, w618);
  FullAdder U128 (w618, w601, IN21[1], w619, w620);
  FullAdder U129 (w620, w602, IN22[0], w621, w622);
  HalfAdder U130 (w605, IN14[9], Out1[14], w624);
  FullAdder U131 (w624, w607, IN15[8], w625, w626);
  FullAdder U132 (w626, w609, IN16[7], w627, w628);
  FullAdder U133 (w628, w611, IN17[6], w629, w630);
  FullAdder U134 (w630, w613, IN18[5], w631, w632);
  FullAdder U135 (w632, w615, IN19[4], w633, w634);
  FullAdder U136 (w634, w617, IN20[3], w635, w636);
  FullAdder U137 (w636, w619, IN21[2], w637, w638);
  FullAdder U138 (w638, w621, IN22[1], w639, w640);
  FullAdder U139 (w640, w622, IN23[0], w641, w642);
  HalfAdder U140 (w625, IN15[9], Out1[15], w644);
  FullAdder U141 (w644, w627, IN16[8], w645, w646);
  FullAdder U142 (w646, w629, IN17[7], w647, w648);
  FullAdder U143 (w648, w631, IN18[6], w649, w650);
  FullAdder U144 (w650, w633, IN19[5], w651, w652);
  FullAdder U145 (w652, w635, IN20[4], w653, w654);
  FullAdder U146 (w654, w637, IN21[3], w655, w656);
  FullAdder U147 (w656, w639, IN22[2], w657, w658);
  FullAdder U148 (w658, w641, IN23[1], w659, w660);
  FullAdder U149 (w660, w642, IN24[0], w661, w662);
  HalfAdder U150 (w645, IN16[9], Out1[16], w664);
  FullAdder U151 (w664, w647, IN17[8], w665, w666);
  FullAdder U152 (w666, w649, IN18[7], w667, w668);
  FullAdder U153 (w668, w651, IN19[6], w669, w670);
  FullAdder U154 (w670, w653, IN20[5], w671, w672);
  FullAdder U155 (w672, w655, IN21[4], w673, w674);
  FullAdder U156 (w674, w657, IN22[3], w675, w676);
  FullAdder U157 (w676, w659, IN23[2], w677, w678);
  FullAdder U158 (w678, w661, IN24[1], w679, w680);
  FullAdder U159 (w680, w662, IN25[0], w681, w682);
  HalfAdder U160 (w665, IN17[9], Out1[17], w684);
  FullAdder U161 (w684, w667, IN18[8], w685, w686);
  FullAdder U162 (w686, w669, IN19[7], w687, w688);
  FullAdder U163 (w688, w671, IN20[6], w689, w690);
  FullAdder U164 (w690, w673, IN21[5], w691, w692);
  FullAdder U165 (w692, w675, IN22[4], w693, w694);
  FullAdder U166 (w694, w677, IN23[3], w695, w696);
  FullAdder U167 (w696, w679, IN24[2], w697, w698);
  FullAdder U168 (w698, w681, IN25[1], w699, w700);
  FullAdder U169 (w700, w682, IN26[0], w701, w702);
  HalfAdder U170 (w685, IN18[9], Out1[18], w704);
  FullAdder U171 (w704, w687, IN19[8], w705, w706);
  FullAdder U172 (w706, w689, IN20[7], w707, w708);
  FullAdder U173 (w708, w691, IN21[6], w709, w710);
  FullAdder U174 (w710, w693, IN22[5], w711, w712);
  FullAdder U175 (w712, w695, IN23[4], w713, w714);
  FullAdder U176 (w714, w697, IN24[3], w715, w716);
  FullAdder U177 (w716, w699, IN25[2], w717, w718);
  FullAdder U178 (w718, w701, IN26[1], w719, w720);
  FullAdder U179 (w720, w702, IN27[0], w721, w722);
  HalfAdder U180 (w705, IN19[9], Out1[19], w724);
  FullAdder U181 (w724, w707, IN20[8], w725, w726);
  FullAdder U182 (w726, w709, IN21[7], w727, w728);
  FullAdder U183 (w728, w711, IN22[6], w729, w730);
  FullAdder U184 (w730, w713, IN23[5], w731, w732);
  FullAdder U185 (w732, w715, IN24[4], w733, w734);
  FullAdder U186 (w734, w717, IN25[3], w735, w736);
  FullAdder U187 (w736, w719, IN26[2], w737, w738);
  FullAdder U188 (w738, w721, IN27[1], w739, w740);
  FullAdder U189 (w740, w722, IN28[0], w741, w742);
  HalfAdder U190 (w725, IN20[9], Out1[20], w744);
  FullAdder U191 (w744, w727, IN21[8], w745, w746);
  FullAdder U192 (w746, w729, IN22[7], w747, w748);
  FullAdder U193 (w748, w731, IN23[6], w749, w750);
  FullAdder U194 (w750, w733, IN24[5], w751, w752);
  FullAdder U195 (w752, w735, IN25[4], w753, w754);
  FullAdder U196 (w754, w737, IN26[3], w755, w756);
  FullAdder U197 (w756, w739, IN27[2], w757, w758);
  FullAdder U198 (w758, w741, IN28[1], w759, w760);
  FullAdder U199 (w760, w742, IN29[0], w761, w762);
  HalfAdder U200 (w745, IN21[9], Out1[21], w764);
  FullAdder U201 (w764, w747, IN22[8], w765, w766);
  FullAdder U202 (w766, w749, IN23[7], w767, w768);
  FullAdder U203 (w768, w751, IN24[6], w769, w770);
  FullAdder U204 (w770, w753, IN25[5], w771, w772);
  FullAdder U205 (w772, w755, IN26[4], w773, w774);
  FullAdder U206 (w774, w757, IN27[3], w775, w776);
  FullAdder U207 (w776, w759, IN28[2], w777, w778);
  FullAdder U208 (w778, w761, IN29[1], w779, w780);
  FullAdder U209 (w780, w762, IN30[0], w781, w782);
  HalfAdder U210 (w765, IN22[9], Out1[22], w784);
  FullAdder U211 (w784, w767, IN23[8], w785, w786);
  FullAdder U212 (w786, w769, IN24[7], w787, w788);
  FullAdder U213 (w788, w771, IN25[6], w789, w790);
  FullAdder U214 (w790, w773, IN26[5], w791, w792);
  FullAdder U215 (w792, w775, IN27[4], w793, w794);
  FullAdder U216 (w794, w777, IN28[3], w795, w796);
  FullAdder U217 (w796, w779, IN29[2], w797, w798);
  FullAdder U218 (w798, w781, IN30[1], w799, w800);
  FullAdder U219 (w800, w782, IN31[0], w801, w802);
  HalfAdder U220 (w785, IN23[9], Out1[23], w804);
  FullAdder U221 (w804, w787, IN24[8], w805, w806);
  FullAdder U222 (w806, w789, IN25[7], w807, w808);
  FullAdder U223 (w808, w791, IN26[6], w809, w810);
  FullAdder U224 (w810, w793, IN27[5], w811, w812);
  FullAdder U225 (w812, w795, IN28[4], w813, w814);
  FullAdder U226 (w814, w797, IN29[3], w815, w816);
  FullAdder U227 (w816, w799, IN30[2], w817, w818);
  FullAdder U228 (w818, w801, IN31[1], w819, w820);
  FullAdder U229 (w820, w802, IN32[0], w821, w822);
  HalfAdder U230 (w805, IN24[9], Out1[24], w824);
  FullAdder U231 (w824, w807, IN25[8], w825, w826);
  FullAdder U232 (w826, w809, IN26[7], w827, w828);
  FullAdder U233 (w828, w811, IN27[6], w829, w830);
  FullAdder U234 (w830, w813, IN28[5], w831, w832);
  FullAdder U235 (w832, w815, IN29[4], w833, w834);
  FullAdder U236 (w834, w817, IN30[3], w835, w836);
  FullAdder U237 (w836, w819, IN31[2], w837, w838);
  FullAdder U238 (w838, w821, IN32[1], w839, w840);
  FullAdder U239 (w840, w822, IN33[0], w841, w842);
  HalfAdder U240 (w825, IN25[9], Out1[25], w844);
  FullAdder U241 (w844, w827, IN26[8], w845, w846);
  FullAdder U242 (w846, w829, IN27[7], w847, w848);
  FullAdder U243 (w848, w831, IN28[6], w849, w850);
  FullAdder U244 (w850, w833, IN29[5], w851, w852);
  FullAdder U245 (w852, w835, IN30[4], w853, w854);
  FullAdder U246 (w854, w837, IN31[3], w855, w856);
  FullAdder U247 (w856, w839, IN32[2], w857, w858);
  FullAdder U248 (w858, w841, IN33[1], w859, w860);
  FullAdder U249 (w860, w842, IN34[0], w861, w862);
  HalfAdder U250 (w845, IN26[9], Out1[26], w864);
  FullAdder U251 (w864, w847, IN27[8], w865, w866);
  FullAdder U252 (w866, w849, IN28[7], w867, w868);
  FullAdder U253 (w868, w851, IN29[6], w869, w870);
  FullAdder U254 (w870, w853, IN30[5], w871, w872);
  FullAdder U255 (w872, w855, IN31[4], w873, w874);
  FullAdder U256 (w874, w857, IN32[3], w875, w876);
  FullAdder U257 (w876, w859, IN33[2], w877, w878);
  FullAdder U258 (w878, w861, IN34[1], w879, w880);
  FullAdder U259 (w880, w862, IN35[0], w881, w882);
  HalfAdder U260 (w865, IN27[9], Out1[27], w884);
  FullAdder U261 (w884, w867, IN28[8], w885, w886);
  FullAdder U262 (w886, w869, IN29[7], w887, w888);
  FullAdder U263 (w888, w871, IN30[6], w889, w890);
  FullAdder U264 (w890, w873, IN31[5], w891, w892);
  FullAdder U265 (w892, w875, IN32[4], w893, w894);
  FullAdder U266 (w894, w877, IN33[3], w895, w896);
  FullAdder U267 (w896, w879, IN34[2], w897, w898);
  FullAdder U268 (w898, w881, IN35[1], w899, w900);
  FullAdder U269 (w900, w882, IN36[0], w901, w902);
  HalfAdder U270 (w885, IN28[9], Out1[28], w904);
  FullAdder U271 (w904, w887, IN29[8], w905, w906);
  FullAdder U272 (w906, w889, IN30[7], w907, w908);
  FullAdder U273 (w908, w891, IN31[6], w909, w910);
  FullAdder U274 (w910, w893, IN32[5], w911, w912);
  FullAdder U275 (w912, w895, IN33[4], w913, w914);
  FullAdder U276 (w914, w897, IN34[3], w915, w916);
  FullAdder U277 (w916, w899, IN35[2], w917, w918);
  FullAdder U278 (w918, w901, IN36[1], w919, w920);
  FullAdder U279 (w920, w902, IN37[0], w921, w922);
  HalfAdder U280 (w905, IN29[9], Out1[29], w924);
  FullAdder U281 (w924, w907, IN30[8], w925, w926);
  FullAdder U282 (w926, w909, IN31[7], w927, w928);
  FullAdder U283 (w928, w911, IN32[6], w929, w930);
  FullAdder U284 (w930, w913, IN33[5], w931, w932);
  FullAdder U285 (w932, w915, IN34[4], w933, w934);
  FullAdder U286 (w934, w917, IN35[3], w935, w936);
  FullAdder U287 (w936, w919, IN36[2], w937, w938);
  FullAdder U288 (w938, w921, IN37[1], w939, w940);
  FullAdder U289 (w940, w922, IN38[0], w941, w942);
  HalfAdder U290 (w925, IN30[9], Out1[30], w944);
  FullAdder U291 (w944, w927, IN31[8], w945, w946);
  FullAdder U292 (w946, w929, IN32[7], w947, w948);
  FullAdder U293 (w948, w931, IN33[6], w949, w950);
  FullAdder U294 (w950, w933, IN34[5], w951, w952);
  FullAdder U295 (w952, w935, IN35[4], w953, w954);
  FullAdder U296 (w954, w937, IN36[3], w955, w956);
  FullAdder U297 (w956, w939, IN37[2], w957, w958);
  FullAdder U298 (w958, w941, IN38[1], w959, w960);
  FullAdder U299 (w960, w942, IN39[0], w961, w962);
  HalfAdder U300 (w945, IN31[9], Out1[31], w964);
  FullAdder U301 (w964, w947, IN32[8], w965, w966);
  FullAdder U302 (w966, w949, IN33[7], w967, w968);
  FullAdder U303 (w968, w951, IN34[6], w969, w970);
  FullAdder U304 (w970, w953, IN35[5], w971, w972);
  FullAdder U305 (w972, w955, IN36[4], w973, w974);
  FullAdder U306 (w974, w957, IN37[3], w975, w976);
  FullAdder U307 (w976, w959, IN38[2], w977, w978);
  FullAdder U308 (w978, w961, IN39[1], w979, w980);
  FullAdder U309 (w980, w962, IN40[0], w981, w982);
  HalfAdder U310 (w965, IN32[9], Out1[32], w984);
  FullAdder U311 (w984, w967, IN33[8], Out1[33], w986);
  FullAdder U312 (w986, w969, IN34[7], Out1[34], w988);
  FullAdder U313 (w988, w971, IN35[6], Out1[35], w990);
  FullAdder U314 (w990, w973, IN36[5], Out1[36], w992);
  FullAdder U315 (w992, w975, IN37[4], Out1[37], w994);
  FullAdder U316 (w994, w977, IN38[3], Out1[38], w996);
  FullAdder U317 (w996, w979, IN39[2], Out1[39], w998);
  FullAdder U318 (w998, w981, IN40[1], Out1[40], w1000);
  FullAdder U319 (w1000, w982, IN41[0], Out1[41], Out1[42]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN11[10];
  assign Out2[1] = IN12[10];
  assign Out2[2] = IN13[10];
  assign Out2[3] = IN14[10];
  assign Out2[4] = IN15[10];
  assign Out2[5] = IN16[10];
  assign Out2[6] = IN17[10];
  assign Out2[7] = IN18[10];
  assign Out2[8] = IN19[10];
  assign Out2[9] = IN20[10];
  assign Out2[10] = IN21[10];
  assign Out2[11] = IN22[10];
  assign Out2[12] = IN23[10];
  assign Out2[13] = IN24[10];
  assign Out2[14] = IN25[10];
  assign Out2[15] = IN26[10];
  assign Out2[16] = IN27[10];
  assign Out2[17] = IN28[10];
  assign Out2[18] = IN29[10];
  assign Out2[19] = IN30[10];
  assign Out2[20] = IN31[10];
  assign Out2[21] = IN32[10];
  assign Out2[22] = IN33[9];
  assign Out2[23] = IN34[8];
  assign Out2[24] = IN35[7];
  assign Out2[25] = IN36[6];
  assign Out2[26] = IN37[5];
  assign Out2[27] = IN38[4];
  assign Out2[28] = IN39[3];
  assign Out2[29] = IN40[2];
  assign Out2[30] = IN41[1];
  assign Out2[31] = IN42[0];

endmodule
module RC_32_32(IN1, IN2, Out);
  input [31:0] IN1;
  input [31:0] IN2;
  output [32:0] Out;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w65);
  FullAdder U1 (IN1[1], IN2[1], w65, Out[1], w67);
  FullAdder U2 (IN1[2], IN2[2], w67, Out[2], w69);
  FullAdder U3 (IN1[3], IN2[3], w69, Out[3], w71);
  FullAdder U4 (IN1[4], IN2[4], w71, Out[4], w73);
  FullAdder U5 (IN1[5], IN2[5], w73, Out[5], w75);
  FullAdder U6 (IN1[6], IN2[6], w75, Out[6], w77);
  FullAdder U7 (IN1[7], IN2[7], w77, Out[7], w79);
  FullAdder U8 (IN1[8], IN2[8], w79, Out[8], w81);
  FullAdder U9 (IN1[9], IN2[9], w81, Out[9], w83);
  FullAdder U10 (IN1[10], IN2[10], w83, Out[10], w85);
  FullAdder U11 (IN1[11], IN2[11], w85, Out[11], w87);
  FullAdder U12 (IN1[12], IN2[12], w87, Out[12], w89);
  FullAdder U13 (IN1[13], IN2[13], w89, Out[13], w91);
  FullAdder U14 (IN1[14], IN2[14], w91, Out[14], w93);
  FullAdder U15 (IN1[15], IN2[15], w93, Out[15], w95);
  FullAdder U16 (IN1[16], IN2[16], w95, Out[16], w97);
  FullAdder U17 (IN1[17], IN2[17], w97, Out[17], w99);
  FullAdder U18 (IN1[18], IN2[18], w99, Out[18], w101);
  FullAdder U19 (IN1[19], IN2[19], w101, Out[19], w103);
  FullAdder U20 (IN1[20], IN2[20], w103, Out[20], w105);
  FullAdder U21 (IN1[21], IN2[21], w105, Out[21], w107);
  FullAdder U22 (IN1[22], IN2[22], w107, Out[22], w109);
  FullAdder U23 (IN1[23], IN2[23], w109, Out[23], w111);
  FullAdder U24 (IN1[24], IN2[24], w111, Out[24], w113);
  FullAdder U25 (IN1[25], IN2[25], w113, Out[25], w115);
  FullAdder U26 (IN1[26], IN2[26], w115, Out[26], w117);
  FullAdder U27 (IN1[27], IN2[27], w117, Out[27], w119);
  FullAdder U28 (IN1[28], IN2[28], w119, Out[28], w121);
  FullAdder U29 (IN1[29], IN2[29], w121, Out[29], w123);
  FullAdder U30 (IN1[30], IN2[30], w123, Out[30], w125);
  FullAdder U31 (IN1[31], IN2[31], w125, Out[31], Out[32]);

endmodule
module NR_11_33(IN1, IN2, Out);
  input [10:0] IN1;
  input [32:0] IN2;
  output [43:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [10:0] P11;
  wire [10:0] P12;
  wire [10:0] P13;
  wire [10:0] P14;
  wire [10:0] P15;
  wire [10:0] P16;
  wire [10:0] P17;
  wire [10:0] P18;
  wire [10:0] P19;
  wire [10:0] P20;
  wire [10:0] P21;
  wire [10:0] P22;
  wire [10:0] P23;
  wire [10:0] P24;
  wire [10:0] P25;
  wire [10:0] P26;
  wire [10:0] P27;
  wire [10:0] P28;
  wire [10:0] P29;
  wire [10:0] P30;
  wire [10:0] P31;
  wire [10:0] P32;
  wire [9:0] P33;
  wire [8:0] P34;
  wire [7:0] P35;
  wire [6:0] P36;
  wire [5:0] P37;
  wire [4:0] P38;
  wire [3:0] P39;
  wire [2:0] P40;
  wire [1:0] P41;
  wire [0:0] P42;
  wire [42:0] R1;
  wire [31:0] R2;
  wire [43:0] aOut;
  U_SP_11_33 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, R1, R2);
  RC_32_32 S2 (R1[42:11], R2, aOut[43:11]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign Out = aOut[43:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
