
module NR_1_50(
    input [0:0]IN1,
    input [49:0]IN2,
    output [49:0]Out
);
    assign Out = IN2;
endmodule
