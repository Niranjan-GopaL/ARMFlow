
module customAdder52_0(
    input [51 : 0] A,
    input [51 : 0] B,
    output [52 : 0] Sum
);

    assign Sum = A+B;

endmodule
