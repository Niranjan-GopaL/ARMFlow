//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 9
  second input length: 37
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_9_37(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  input [8:0] IN1;
  input [36:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [8:0] P9;
  output [8:0] P10;
  output [8:0] P11;
  output [8:0] P12;
  output [8:0] P13;
  output [8:0] P14;
  output [8:0] P15;
  output [8:0] P16;
  output [8:0] P17;
  output [8:0] P18;
  output [8:0] P19;
  output [8:0] P20;
  output [8:0] P21;
  output [8:0] P22;
  output [8:0] P23;
  output [8:0] P24;
  output [8:0] P25;
  output [8:0] P26;
  output [8:0] P27;
  output [8:0] P28;
  output [8:0] P29;
  output [8:0] P30;
  output [8:0] P31;
  output [8:0] P32;
  output [8:0] P33;
  output [8:0] P34;
  output [8:0] P35;
  output [8:0] P36;
  output [7:0] P37;
  output [6:0] P38;
  output [5:0] P39;
  output [4:0] P40;
  output [3:0] P41;
  output [2:0] P42;
  output [1:0] P43;
  output [0:0] P44;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[0] = IN1[1]&IN2[36];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[1] = IN1[2]&IN2[35];
  assign P38[0] = IN1[2]&IN2[36];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[2] = IN1[3]&IN2[34];
  assign P38[1] = IN1[3]&IN2[35];
  assign P39[0] = IN1[3]&IN2[36];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[3] = IN1[4]&IN2[33];
  assign P38[2] = IN1[4]&IN2[34];
  assign P39[1] = IN1[4]&IN2[35];
  assign P40[0] = IN1[4]&IN2[36];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[4] = IN1[5]&IN2[32];
  assign P38[3] = IN1[5]&IN2[33];
  assign P39[2] = IN1[5]&IN2[34];
  assign P40[1] = IN1[5]&IN2[35];
  assign P41[0] = IN1[5]&IN2[36];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[5] = IN1[6]&IN2[31];
  assign P38[4] = IN1[6]&IN2[32];
  assign P39[3] = IN1[6]&IN2[33];
  assign P40[2] = IN1[6]&IN2[34];
  assign P41[1] = IN1[6]&IN2[35];
  assign P42[0] = IN1[6]&IN2[36];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[6] = IN1[7]&IN2[30];
  assign P38[5] = IN1[7]&IN2[31];
  assign P39[4] = IN1[7]&IN2[32];
  assign P40[3] = IN1[7]&IN2[33];
  assign P41[2] = IN1[7]&IN2[34];
  assign P42[1] = IN1[7]&IN2[35];
  assign P43[0] = IN1[7]&IN2[36];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[7] = IN1[8]&IN2[29];
  assign P38[6] = IN1[8]&IN2[30];
  assign P39[5] = IN1[8]&IN2[31];
  assign P40[4] = IN1[8]&IN2[32];
  assign P41[3] = IN1[8]&IN2[33];
  assign P42[2] = IN1[8]&IN2[34];
  assign P43[1] = IN1[8]&IN2[35];
  assign P44[0] = IN1[8]&IN2[36];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [8:0] IN9;
  input [8:0] IN10;
  input [8:0] IN11;
  input [8:0] IN12;
  input [8:0] IN13;
  input [8:0] IN14;
  input [8:0] IN15;
  input [8:0] IN16;
  input [8:0] IN17;
  input [8:0] IN18;
  input [8:0] IN19;
  input [8:0] IN20;
  input [8:0] IN21;
  input [8:0] IN22;
  input [8:0] IN23;
  input [8:0] IN24;
  input [8:0] IN25;
  input [8:0] IN26;
  input [8:0] IN27;
  input [8:0] IN28;
  input [8:0] IN29;
  input [8:0] IN30;
  input [8:0] IN31;
  input [8:0] IN32;
  input [8:0] IN33;
  input [8:0] IN34;
  input [8:0] IN35;
  input [8:0] IN36;
  input [7:0] IN37;
  input [6:0] IN38;
  input [5:0] IN39;
  input [4:0] IN40;
  input [3:0] IN41;
  input [2:0] IN42;
  input [1:0] IN43;
  input [0:0] IN44;
  output [44:0] Out1;
  output [35:0] Out2;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w645;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w693;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w741;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w789;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w837;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w885;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w894;
  wire w896;
  wire w898;
  wire w900;
  wire w902;
  wire w904;
  wire w906;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w334);
  FullAdder U1 (w334, IN2[0], IN2[1], w335, w336);
  FullAdder U2 (w336, IN3[0], IN3[1], w337, w338);
  FullAdder U3 (w338, IN4[0], IN4[1], w339, w340);
  FullAdder U4 (w340, IN5[0], IN5[1], w341, w342);
  FullAdder U5 (w342, IN6[0], IN6[1], w343, w344);
  FullAdder U6 (w344, IN7[0], IN7[1], w345, w346);
  FullAdder U7 (w346, IN8[0], IN8[1], w347, w348);
  HalfAdder U8 (w335, IN2[2], Out1[2], w350);
  FullAdder U9 (w350, w337, IN3[2], w351, w352);
  FullAdder U10 (w352, w339, IN4[2], w353, w354);
  FullAdder U11 (w354, w341, IN5[2], w355, w356);
  FullAdder U12 (w356, w343, IN6[2], w357, w358);
  FullAdder U13 (w358, w345, IN7[2], w359, w360);
  FullAdder U14 (w360, w347, IN8[2], w361, w362);
  FullAdder U15 (w362, w348, IN9[0], w363, w364);
  HalfAdder U16 (w351, IN3[3], Out1[3], w366);
  FullAdder U17 (w366, w353, IN4[3], w367, w368);
  FullAdder U18 (w368, w355, IN5[3], w369, w370);
  FullAdder U19 (w370, w357, IN6[3], w371, w372);
  FullAdder U20 (w372, w359, IN7[3], w373, w374);
  FullAdder U21 (w374, w361, IN8[3], w375, w376);
  FullAdder U22 (w376, w363, IN9[1], w377, w378);
  FullAdder U23 (w378, w364, IN10[0], w379, w380);
  HalfAdder U24 (w367, IN4[4], Out1[4], w382);
  FullAdder U25 (w382, w369, IN5[4], w383, w384);
  FullAdder U26 (w384, w371, IN6[4], w385, w386);
  FullAdder U27 (w386, w373, IN7[4], w387, w388);
  FullAdder U28 (w388, w375, IN8[4], w389, w390);
  FullAdder U29 (w390, w377, IN9[2], w391, w392);
  FullAdder U30 (w392, w379, IN10[1], w393, w394);
  FullAdder U31 (w394, w380, IN11[0], w395, w396);
  HalfAdder U32 (w383, IN5[5], Out1[5], w398);
  FullAdder U33 (w398, w385, IN6[5], w399, w400);
  FullAdder U34 (w400, w387, IN7[5], w401, w402);
  FullAdder U35 (w402, w389, IN8[5], w403, w404);
  FullAdder U36 (w404, w391, IN9[3], w405, w406);
  FullAdder U37 (w406, w393, IN10[2], w407, w408);
  FullAdder U38 (w408, w395, IN11[1], w409, w410);
  FullAdder U39 (w410, w396, IN12[0], w411, w412);
  HalfAdder U40 (w399, IN6[6], Out1[6], w414);
  FullAdder U41 (w414, w401, IN7[6], w415, w416);
  FullAdder U42 (w416, w403, IN8[6], w417, w418);
  FullAdder U43 (w418, w405, IN9[4], w419, w420);
  FullAdder U44 (w420, w407, IN10[3], w421, w422);
  FullAdder U45 (w422, w409, IN11[2], w423, w424);
  FullAdder U46 (w424, w411, IN12[1], w425, w426);
  FullAdder U47 (w426, w412, IN13[0], w427, w428);
  HalfAdder U48 (w415, IN7[7], Out1[7], w430);
  FullAdder U49 (w430, w417, IN8[7], w431, w432);
  FullAdder U50 (w432, w419, IN9[5], w433, w434);
  FullAdder U51 (w434, w421, IN10[4], w435, w436);
  FullAdder U52 (w436, w423, IN11[3], w437, w438);
  FullAdder U53 (w438, w425, IN12[2], w439, w440);
  FullAdder U54 (w440, w427, IN13[1], w441, w442);
  FullAdder U55 (w442, w428, IN14[0], w443, w444);
  HalfAdder U56 (w431, IN8[8], Out1[8], w446);
  FullAdder U57 (w446, w433, IN9[6], w447, w448);
  FullAdder U58 (w448, w435, IN10[5], w449, w450);
  FullAdder U59 (w450, w437, IN11[4], w451, w452);
  FullAdder U60 (w452, w439, IN12[3], w453, w454);
  FullAdder U61 (w454, w441, IN13[2], w455, w456);
  FullAdder U62 (w456, w443, IN14[1], w457, w458);
  FullAdder U63 (w458, w444, IN15[0], w459, w460);
  HalfAdder U64 (w447, IN9[7], Out1[9], w462);
  FullAdder U65 (w462, w449, IN10[6], w463, w464);
  FullAdder U66 (w464, w451, IN11[5], w465, w466);
  FullAdder U67 (w466, w453, IN12[4], w467, w468);
  FullAdder U68 (w468, w455, IN13[3], w469, w470);
  FullAdder U69 (w470, w457, IN14[2], w471, w472);
  FullAdder U70 (w472, w459, IN15[1], w473, w474);
  FullAdder U71 (w474, w460, IN16[0], w475, w476);
  HalfAdder U72 (w463, IN10[7], Out1[10], w478);
  FullAdder U73 (w478, w465, IN11[6], w479, w480);
  FullAdder U74 (w480, w467, IN12[5], w481, w482);
  FullAdder U75 (w482, w469, IN13[4], w483, w484);
  FullAdder U76 (w484, w471, IN14[3], w485, w486);
  FullAdder U77 (w486, w473, IN15[2], w487, w488);
  FullAdder U78 (w488, w475, IN16[1], w489, w490);
  FullAdder U79 (w490, w476, IN17[0], w491, w492);
  HalfAdder U80 (w479, IN11[7], Out1[11], w494);
  FullAdder U81 (w494, w481, IN12[6], w495, w496);
  FullAdder U82 (w496, w483, IN13[5], w497, w498);
  FullAdder U83 (w498, w485, IN14[4], w499, w500);
  FullAdder U84 (w500, w487, IN15[3], w501, w502);
  FullAdder U85 (w502, w489, IN16[2], w503, w504);
  FullAdder U86 (w504, w491, IN17[1], w505, w506);
  FullAdder U87 (w506, w492, IN18[0], w507, w508);
  HalfAdder U88 (w495, IN12[7], Out1[12], w510);
  FullAdder U89 (w510, w497, IN13[6], w511, w512);
  FullAdder U90 (w512, w499, IN14[5], w513, w514);
  FullAdder U91 (w514, w501, IN15[4], w515, w516);
  FullAdder U92 (w516, w503, IN16[3], w517, w518);
  FullAdder U93 (w518, w505, IN17[2], w519, w520);
  FullAdder U94 (w520, w507, IN18[1], w521, w522);
  FullAdder U95 (w522, w508, IN19[0], w523, w524);
  HalfAdder U96 (w511, IN13[7], Out1[13], w526);
  FullAdder U97 (w526, w513, IN14[6], w527, w528);
  FullAdder U98 (w528, w515, IN15[5], w529, w530);
  FullAdder U99 (w530, w517, IN16[4], w531, w532);
  FullAdder U100 (w532, w519, IN17[3], w533, w534);
  FullAdder U101 (w534, w521, IN18[2], w535, w536);
  FullAdder U102 (w536, w523, IN19[1], w537, w538);
  FullAdder U103 (w538, w524, IN20[0], w539, w540);
  HalfAdder U104 (w527, IN14[7], Out1[14], w542);
  FullAdder U105 (w542, w529, IN15[6], w543, w544);
  FullAdder U106 (w544, w531, IN16[5], w545, w546);
  FullAdder U107 (w546, w533, IN17[4], w547, w548);
  FullAdder U108 (w548, w535, IN18[3], w549, w550);
  FullAdder U109 (w550, w537, IN19[2], w551, w552);
  FullAdder U110 (w552, w539, IN20[1], w553, w554);
  FullAdder U111 (w554, w540, IN21[0], w555, w556);
  HalfAdder U112 (w543, IN15[7], Out1[15], w558);
  FullAdder U113 (w558, w545, IN16[6], w559, w560);
  FullAdder U114 (w560, w547, IN17[5], w561, w562);
  FullAdder U115 (w562, w549, IN18[4], w563, w564);
  FullAdder U116 (w564, w551, IN19[3], w565, w566);
  FullAdder U117 (w566, w553, IN20[2], w567, w568);
  FullAdder U118 (w568, w555, IN21[1], w569, w570);
  FullAdder U119 (w570, w556, IN22[0], w571, w572);
  HalfAdder U120 (w559, IN16[7], Out1[16], w574);
  FullAdder U121 (w574, w561, IN17[6], w575, w576);
  FullAdder U122 (w576, w563, IN18[5], w577, w578);
  FullAdder U123 (w578, w565, IN19[4], w579, w580);
  FullAdder U124 (w580, w567, IN20[3], w581, w582);
  FullAdder U125 (w582, w569, IN21[2], w583, w584);
  FullAdder U126 (w584, w571, IN22[1], w585, w586);
  FullAdder U127 (w586, w572, IN23[0], w587, w588);
  HalfAdder U128 (w575, IN17[7], Out1[17], w590);
  FullAdder U129 (w590, w577, IN18[6], w591, w592);
  FullAdder U130 (w592, w579, IN19[5], w593, w594);
  FullAdder U131 (w594, w581, IN20[4], w595, w596);
  FullAdder U132 (w596, w583, IN21[3], w597, w598);
  FullAdder U133 (w598, w585, IN22[2], w599, w600);
  FullAdder U134 (w600, w587, IN23[1], w601, w602);
  FullAdder U135 (w602, w588, IN24[0], w603, w604);
  HalfAdder U136 (w591, IN18[7], Out1[18], w606);
  FullAdder U137 (w606, w593, IN19[6], w607, w608);
  FullAdder U138 (w608, w595, IN20[5], w609, w610);
  FullAdder U139 (w610, w597, IN21[4], w611, w612);
  FullAdder U140 (w612, w599, IN22[3], w613, w614);
  FullAdder U141 (w614, w601, IN23[2], w615, w616);
  FullAdder U142 (w616, w603, IN24[1], w617, w618);
  FullAdder U143 (w618, w604, IN25[0], w619, w620);
  HalfAdder U144 (w607, IN19[7], Out1[19], w622);
  FullAdder U145 (w622, w609, IN20[6], w623, w624);
  FullAdder U146 (w624, w611, IN21[5], w625, w626);
  FullAdder U147 (w626, w613, IN22[4], w627, w628);
  FullAdder U148 (w628, w615, IN23[3], w629, w630);
  FullAdder U149 (w630, w617, IN24[2], w631, w632);
  FullAdder U150 (w632, w619, IN25[1], w633, w634);
  FullAdder U151 (w634, w620, IN26[0], w635, w636);
  HalfAdder U152 (w623, IN20[7], Out1[20], w638);
  FullAdder U153 (w638, w625, IN21[6], w639, w640);
  FullAdder U154 (w640, w627, IN22[5], w641, w642);
  FullAdder U155 (w642, w629, IN23[4], w643, w644);
  FullAdder U156 (w644, w631, IN24[3], w645, w646);
  FullAdder U157 (w646, w633, IN25[2], w647, w648);
  FullAdder U158 (w648, w635, IN26[1], w649, w650);
  FullAdder U159 (w650, w636, IN27[0], w651, w652);
  HalfAdder U160 (w639, IN21[7], Out1[21], w654);
  FullAdder U161 (w654, w641, IN22[6], w655, w656);
  FullAdder U162 (w656, w643, IN23[5], w657, w658);
  FullAdder U163 (w658, w645, IN24[4], w659, w660);
  FullAdder U164 (w660, w647, IN25[3], w661, w662);
  FullAdder U165 (w662, w649, IN26[2], w663, w664);
  FullAdder U166 (w664, w651, IN27[1], w665, w666);
  FullAdder U167 (w666, w652, IN28[0], w667, w668);
  HalfAdder U168 (w655, IN22[7], Out1[22], w670);
  FullAdder U169 (w670, w657, IN23[6], w671, w672);
  FullAdder U170 (w672, w659, IN24[5], w673, w674);
  FullAdder U171 (w674, w661, IN25[4], w675, w676);
  FullAdder U172 (w676, w663, IN26[3], w677, w678);
  FullAdder U173 (w678, w665, IN27[2], w679, w680);
  FullAdder U174 (w680, w667, IN28[1], w681, w682);
  FullAdder U175 (w682, w668, IN29[0], w683, w684);
  HalfAdder U176 (w671, IN23[7], Out1[23], w686);
  FullAdder U177 (w686, w673, IN24[6], w687, w688);
  FullAdder U178 (w688, w675, IN25[5], w689, w690);
  FullAdder U179 (w690, w677, IN26[4], w691, w692);
  FullAdder U180 (w692, w679, IN27[3], w693, w694);
  FullAdder U181 (w694, w681, IN28[2], w695, w696);
  FullAdder U182 (w696, w683, IN29[1], w697, w698);
  FullAdder U183 (w698, w684, IN30[0], w699, w700);
  HalfAdder U184 (w687, IN24[7], Out1[24], w702);
  FullAdder U185 (w702, w689, IN25[6], w703, w704);
  FullAdder U186 (w704, w691, IN26[5], w705, w706);
  FullAdder U187 (w706, w693, IN27[4], w707, w708);
  FullAdder U188 (w708, w695, IN28[3], w709, w710);
  FullAdder U189 (w710, w697, IN29[2], w711, w712);
  FullAdder U190 (w712, w699, IN30[1], w713, w714);
  FullAdder U191 (w714, w700, IN31[0], w715, w716);
  HalfAdder U192 (w703, IN25[7], Out1[25], w718);
  FullAdder U193 (w718, w705, IN26[6], w719, w720);
  FullAdder U194 (w720, w707, IN27[5], w721, w722);
  FullAdder U195 (w722, w709, IN28[4], w723, w724);
  FullAdder U196 (w724, w711, IN29[3], w725, w726);
  FullAdder U197 (w726, w713, IN30[2], w727, w728);
  FullAdder U198 (w728, w715, IN31[1], w729, w730);
  FullAdder U199 (w730, w716, IN32[0], w731, w732);
  HalfAdder U200 (w719, IN26[7], Out1[26], w734);
  FullAdder U201 (w734, w721, IN27[6], w735, w736);
  FullAdder U202 (w736, w723, IN28[5], w737, w738);
  FullAdder U203 (w738, w725, IN29[4], w739, w740);
  FullAdder U204 (w740, w727, IN30[3], w741, w742);
  FullAdder U205 (w742, w729, IN31[2], w743, w744);
  FullAdder U206 (w744, w731, IN32[1], w745, w746);
  FullAdder U207 (w746, w732, IN33[0], w747, w748);
  HalfAdder U208 (w735, IN27[7], Out1[27], w750);
  FullAdder U209 (w750, w737, IN28[6], w751, w752);
  FullAdder U210 (w752, w739, IN29[5], w753, w754);
  FullAdder U211 (w754, w741, IN30[4], w755, w756);
  FullAdder U212 (w756, w743, IN31[3], w757, w758);
  FullAdder U213 (w758, w745, IN32[2], w759, w760);
  FullAdder U214 (w760, w747, IN33[1], w761, w762);
  FullAdder U215 (w762, w748, IN34[0], w763, w764);
  HalfAdder U216 (w751, IN28[7], Out1[28], w766);
  FullAdder U217 (w766, w753, IN29[6], w767, w768);
  FullAdder U218 (w768, w755, IN30[5], w769, w770);
  FullAdder U219 (w770, w757, IN31[4], w771, w772);
  FullAdder U220 (w772, w759, IN32[3], w773, w774);
  FullAdder U221 (w774, w761, IN33[2], w775, w776);
  FullAdder U222 (w776, w763, IN34[1], w777, w778);
  FullAdder U223 (w778, w764, IN35[0], w779, w780);
  HalfAdder U224 (w767, IN29[7], Out1[29], w782);
  FullAdder U225 (w782, w769, IN30[6], w783, w784);
  FullAdder U226 (w784, w771, IN31[5], w785, w786);
  FullAdder U227 (w786, w773, IN32[4], w787, w788);
  FullAdder U228 (w788, w775, IN33[3], w789, w790);
  FullAdder U229 (w790, w777, IN34[2], w791, w792);
  FullAdder U230 (w792, w779, IN35[1], w793, w794);
  FullAdder U231 (w794, w780, IN36[0], w795, w796);
  HalfAdder U232 (w783, IN30[7], Out1[30], w798);
  FullAdder U233 (w798, w785, IN31[6], w799, w800);
  FullAdder U234 (w800, w787, IN32[5], w801, w802);
  FullAdder U235 (w802, w789, IN33[4], w803, w804);
  FullAdder U236 (w804, w791, IN34[3], w805, w806);
  FullAdder U237 (w806, w793, IN35[2], w807, w808);
  FullAdder U238 (w808, w795, IN36[1], w809, w810);
  FullAdder U239 (w810, w796, IN37[0], w811, w812);
  HalfAdder U240 (w799, IN31[7], Out1[31], w814);
  FullAdder U241 (w814, w801, IN32[6], w815, w816);
  FullAdder U242 (w816, w803, IN33[5], w817, w818);
  FullAdder U243 (w818, w805, IN34[4], w819, w820);
  FullAdder U244 (w820, w807, IN35[3], w821, w822);
  FullAdder U245 (w822, w809, IN36[2], w823, w824);
  FullAdder U246 (w824, w811, IN37[1], w825, w826);
  FullAdder U247 (w826, w812, IN38[0], w827, w828);
  HalfAdder U248 (w815, IN32[7], Out1[32], w830);
  FullAdder U249 (w830, w817, IN33[6], w831, w832);
  FullAdder U250 (w832, w819, IN34[5], w833, w834);
  FullAdder U251 (w834, w821, IN35[4], w835, w836);
  FullAdder U252 (w836, w823, IN36[3], w837, w838);
  FullAdder U253 (w838, w825, IN37[2], w839, w840);
  FullAdder U254 (w840, w827, IN38[1], w841, w842);
  FullAdder U255 (w842, w828, IN39[0], w843, w844);
  HalfAdder U256 (w831, IN33[7], Out1[33], w846);
  FullAdder U257 (w846, w833, IN34[6], w847, w848);
  FullAdder U258 (w848, w835, IN35[5], w849, w850);
  FullAdder U259 (w850, w837, IN36[4], w851, w852);
  FullAdder U260 (w852, w839, IN37[3], w853, w854);
  FullAdder U261 (w854, w841, IN38[2], w855, w856);
  FullAdder U262 (w856, w843, IN39[1], w857, w858);
  FullAdder U263 (w858, w844, IN40[0], w859, w860);
  HalfAdder U264 (w847, IN34[7], Out1[34], w862);
  FullAdder U265 (w862, w849, IN35[6], w863, w864);
  FullAdder U266 (w864, w851, IN36[5], w865, w866);
  FullAdder U267 (w866, w853, IN37[4], w867, w868);
  FullAdder U268 (w868, w855, IN38[3], w869, w870);
  FullAdder U269 (w870, w857, IN39[2], w871, w872);
  FullAdder U270 (w872, w859, IN40[1], w873, w874);
  FullAdder U271 (w874, w860, IN41[0], w875, w876);
  HalfAdder U272 (w863, IN35[7], Out1[35], w878);
  FullAdder U273 (w878, w865, IN36[6], w879, w880);
  FullAdder U274 (w880, w867, IN37[5], w881, w882);
  FullAdder U275 (w882, w869, IN38[4], w883, w884);
  FullAdder U276 (w884, w871, IN39[3], w885, w886);
  FullAdder U277 (w886, w873, IN40[2], w887, w888);
  FullAdder U278 (w888, w875, IN41[1], w889, w890);
  FullAdder U279 (w890, w876, IN42[0], w891, w892);
  HalfAdder U280 (w879, IN36[7], Out1[36], w894);
  FullAdder U281 (w894, w881, IN37[6], Out1[37], w896);
  FullAdder U282 (w896, w883, IN38[5], Out1[38], w898);
  FullAdder U283 (w898, w885, IN39[4], Out1[39], w900);
  FullAdder U284 (w900, w887, IN40[3], Out1[40], w902);
  FullAdder U285 (w902, w889, IN41[2], Out1[41], w904);
  FullAdder U286 (w904, w891, IN42[1], Out1[42], w906);
  FullAdder U287 (w906, w892, IN43[0], Out1[43], Out1[44]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN9[8];
  assign Out2[1] = IN10[8];
  assign Out2[2] = IN11[8];
  assign Out2[3] = IN12[8];
  assign Out2[4] = IN13[8];
  assign Out2[5] = IN14[8];
  assign Out2[6] = IN15[8];
  assign Out2[7] = IN16[8];
  assign Out2[8] = IN17[8];
  assign Out2[9] = IN18[8];
  assign Out2[10] = IN19[8];
  assign Out2[11] = IN20[8];
  assign Out2[12] = IN21[8];
  assign Out2[13] = IN22[8];
  assign Out2[14] = IN23[8];
  assign Out2[15] = IN24[8];
  assign Out2[16] = IN25[8];
  assign Out2[17] = IN26[8];
  assign Out2[18] = IN27[8];
  assign Out2[19] = IN28[8];
  assign Out2[20] = IN29[8];
  assign Out2[21] = IN30[8];
  assign Out2[22] = IN31[8];
  assign Out2[23] = IN32[8];
  assign Out2[24] = IN33[8];
  assign Out2[25] = IN34[8];
  assign Out2[26] = IN35[8];
  assign Out2[27] = IN36[8];
  assign Out2[28] = IN37[7];
  assign Out2[29] = IN38[6];
  assign Out2[30] = IN39[5];
  assign Out2[31] = IN40[4];
  assign Out2[32] = IN41[3];
  assign Out2[33] = IN42[2];
  assign Out2[34] = IN43[1];
  assign Out2[35] = IN44[0];

endmodule
module RC_36_36(IN1, IN2, Out);
  input [35:0] IN1;
  input [35:0] IN2;
  output [36:0] Out;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w73);
  FullAdder U1 (IN1[1], IN2[1], w73, Out[1], w75);
  FullAdder U2 (IN1[2], IN2[2], w75, Out[2], w77);
  FullAdder U3 (IN1[3], IN2[3], w77, Out[3], w79);
  FullAdder U4 (IN1[4], IN2[4], w79, Out[4], w81);
  FullAdder U5 (IN1[5], IN2[5], w81, Out[5], w83);
  FullAdder U6 (IN1[6], IN2[6], w83, Out[6], w85);
  FullAdder U7 (IN1[7], IN2[7], w85, Out[7], w87);
  FullAdder U8 (IN1[8], IN2[8], w87, Out[8], w89);
  FullAdder U9 (IN1[9], IN2[9], w89, Out[9], w91);
  FullAdder U10 (IN1[10], IN2[10], w91, Out[10], w93);
  FullAdder U11 (IN1[11], IN2[11], w93, Out[11], w95);
  FullAdder U12 (IN1[12], IN2[12], w95, Out[12], w97);
  FullAdder U13 (IN1[13], IN2[13], w97, Out[13], w99);
  FullAdder U14 (IN1[14], IN2[14], w99, Out[14], w101);
  FullAdder U15 (IN1[15], IN2[15], w101, Out[15], w103);
  FullAdder U16 (IN1[16], IN2[16], w103, Out[16], w105);
  FullAdder U17 (IN1[17], IN2[17], w105, Out[17], w107);
  FullAdder U18 (IN1[18], IN2[18], w107, Out[18], w109);
  FullAdder U19 (IN1[19], IN2[19], w109, Out[19], w111);
  FullAdder U20 (IN1[20], IN2[20], w111, Out[20], w113);
  FullAdder U21 (IN1[21], IN2[21], w113, Out[21], w115);
  FullAdder U22 (IN1[22], IN2[22], w115, Out[22], w117);
  FullAdder U23 (IN1[23], IN2[23], w117, Out[23], w119);
  FullAdder U24 (IN1[24], IN2[24], w119, Out[24], w121);
  FullAdder U25 (IN1[25], IN2[25], w121, Out[25], w123);
  FullAdder U26 (IN1[26], IN2[26], w123, Out[26], w125);
  FullAdder U27 (IN1[27], IN2[27], w125, Out[27], w127);
  FullAdder U28 (IN1[28], IN2[28], w127, Out[28], w129);
  FullAdder U29 (IN1[29], IN2[29], w129, Out[29], w131);
  FullAdder U30 (IN1[30], IN2[30], w131, Out[30], w133);
  FullAdder U31 (IN1[31], IN2[31], w133, Out[31], w135);
  FullAdder U32 (IN1[32], IN2[32], w135, Out[32], w137);
  FullAdder U33 (IN1[33], IN2[33], w137, Out[33], w139);
  FullAdder U34 (IN1[34], IN2[34], w139, Out[34], w141);
  FullAdder U35 (IN1[35], IN2[35], w141, Out[35], Out[36]);

endmodule
module NR_9_37(IN1, IN2, Out);
  input [8:0] IN1;
  input [36:0] IN2;
  output [45:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [8:0] P9;
  wire [8:0] P10;
  wire [8:0] P11;
  wire [8:0] P12;
  wire [8:0] P13;
  wire [8:0] P14;
  wire [8:0] P15;
  wire [8:0] P16;
  wire [8:0] P17;
  wire [8:0] P18;
  wire [8:0] P19;
  wire [8:0] P20;
  wire [8:0] P21;
  wire [8:0] P22;
  wire [8:0] P23;
  wire [8:0] P24;
  wire [8:0] P25;
  wire [8:0] P26;
  wire [8:0] P27;
  wire [8:0] P28;
  wire [8:0] P29;
  wire [8:0] P30;
  wire [8:0] P31;
  wire [8:0] P32;
  wire [8:0] P33;
  wire [8:0] P34;
  wire [8:0] P35;
  wire [8:0] P36;
  wire [7:0] P37;
  wire [6:0] P38;
  wire [5:0] P39;
  wire [4:0] P40;
  wire [3:0] P41;
  wire [2:0] P42;
  wire [1:0] P43;
  wire [0:0] P44;
  wire [44:0] R1;
  wire [35:0] R2;
  wire [45:0] aOut;
  U_SP_9_37 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, R1, R2);
  RC_36_36 S2 (R1[44:9], R2, aOut[45:9]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign Out = aOut[45:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
