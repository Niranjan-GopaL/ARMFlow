//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 13
  second input length: 33
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_13_33(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  input [12:0] IN1;
  input [32:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  output [12:0] P17;
  output [12:0] P18;
  output [12:0] P19;
  output [12:0] P20;
  output [12:0] P21;
  output [12:0] P22;
  output [12:0] P23;
  output [12:0] P24;
  output [12:0] P25;
  output [12:0] P26;
  output [12:0] P27;
  output [12:0] P28;
  output [12:0] P29;
  output [12:0] P30;
  output [12:0] P31;
  output [12:0] P32;
  output [11:0] P33;
  output [10:0] P34;
  output [9:0] P35;
  output [8:0] P36;
  output [7:0] P37;
  output [6:0] P38;
  output [5:0] P39;
  output [4:0] P40;
  output [3:0] P41;
  output [2:0] P42;
  output [1:0] P43;
  output [0:0] P44;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[0] = IN1[1]&IN2[32];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[1] = IN1[2]&IN2[31];
  assign P34[0] = IN1[2]&IN2[32];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[2] = IN1[3]&IN2[30];
  assign P34[1] = IN1[3]&IN2[31];
  assign P35[0] = IN1[3]&IN2[32];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[3] = IN1[4]&IN2[29];
  assign P34[2] = IN1[4]&IN2[30];
  assign P35[1] = IN1[4]&IN2[31];
  assign P36[0] = IN1[4]&IN2[32];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[4] = IN1[5]&IN2[28];
  assign P34[3] = IN1[5]&IN2[29];
  assign P35[2] = IN1[5]&IN2[30];
  assign P36[1] = IN1[5]&IN2[31];
  assign P37[0] = IN1[5]&IN2[32];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[5] = IN1[6]&IN2[27];
  assign P34[4] = IN1[6]&IN2[28];
  assign P35[3] = IN1[6]&IN2[29];
  assign P36[2] = IN1[6]&IN2[30];
  assign P37[1] = IN1[6]&IN2[31];
  assign P38[0] = IN1[6]&IN2[32];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[6] = IN1[7]&IN2[26];
  assign P34[5] = IN1[7]&IN2[27];
  assign P35[4] = IN1[7]&IN2[28];
  assign P36[3] = IN1[7]&IN2[29];
  assign P37[2] = IN1[7]&IN2[30];
  assign P38[1] = IN1[7]&IN2[31];
  assign P39[0] = IN1[7]&IN2[32];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[7] = IN1[8]&IN2[25];
  assign P34[6] = IN1[8]&IN2[26];
  assign P35[5] = IN1[8]&IN2[27];
  assign P36[4] = IN1[8]&IN2[28];
  assign P37[3] = IN1[8]&IN2[29];
  assign P38[2] = IN1[8]&IN2[30];
  assign P39[1] = IN1[8]&IN2[31];
  assign P40[0] = IN1[8]&IN2[32];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[8] = IN1[9]&IN2[24];
  assign P34[7] = IN1[9]&IN2[25];
  assign P35[6] = IN1[9]&IN2[26];
  assign P36[5] = IN1[9]&IN2[27];
  assign P37[4] = IN1[9]&IN2[28];
  assign P38[3] = IN1[9]&IN2[29];
  assign P39[2] = IN1[9]&IN2[30];
  assign P40[1] = IN1[9]&IN2[31];
  assign P41[0] = IN1[9]&IN2[32];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[9] = IN1[10]&IN2[23];
  assign P34[8] = IN1[10]&IN2[24];
  assign P35[7] = IN1[10]&IN2[25];
  assign P36[6] = IN1[10]&IN2[26];
  assign P37[5] = IN1[10]&IN2[27];
  assign P38[4] = IN1[10]&IN2[28];
  assign P39[3] = IN1[10]&IN2[29];
  assign P40[2] = IN1[10]&IN2[30];
  assign P41[1] = IN1[10]&IN2[31];
  assign P42[0] = IN1[10]&IN2[32];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[10] = IN1[11]&IN2[22];
  assign P34[9] = IN1[11]&IN2[23];
  assign P35[8] = IN1[11]&IN2[24];
  assign P36[7] = IN1[11]&IN2[25];
  assign P37[6] = IN1[11]&IN2[26];
  assign P38[5] = IN1[11]&IN2[27];
  assign P39[4] = IN1[11]&IN2[28];
  assign P40[3] = IN1[11]&IN2[29];
  assign P41[2] = IN1[11]&IN2[30];
  assign P42[1] = IN1[11]&IN2[31];
  assign P43[0] = IN1[11]&IN2[32];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[11] = IN1[12]&IN2[21];
  assign P34[10] = IN1[12]&IN2[22];
  assign P35[9] = IN1[12]&IN2[23];
  assign P36[8] = IN1[12]&IN2[24];
  assign P37[7] = IN1[12]&IN2[25];
  assign P38[6] = IN1[12]&IN2[26];
  assign P39[5] = IN1[12]&IN2[27];
  assign P40[4] = IN1[12]&IN2[28];
  assign P41[3] = IN1[12]&IN2[29];
  assign P42[2] = IN1[12]&IN2[30];
  assign P43[1] = IN1[12]&IN2[31];
  assign P44[0] = IN1[12]&IN2[32];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [12:0] IN13;
  input [12:0] IN14;
  input [12:0] IN15;
  input [12:0] IN16;
  input [12:0] IN17;
  input [12:0] IN18;
  input [12:0] IN19;
  input [12:0] IN20;
  input [12:0] IN21;
  input [12:0] IN22;
  input [12:0] IN23;
  input [12:0] IN24;
  input [12:0] IN25;
  input [12:0] IN26;
  input [12:0] IN27;
  input [12:0] IN28;
  input [12:0] IN29;
  input [12:0] IN30;
  input [12:0] IN31;
  input [12:0] IN32;
  input [11:0] IN33;
  input [10:0] IN34;
  input [9:0] IN35;
  input [8:0] IN36;
  input [7:0] IN37;
  input [6:0] IN38;
  input [5:0] IN39;
  input [4:0] IN40;
  input [3:0] IN41;
  input [2:0] IN42;
  input [1:0] IN43;
  input [0:0] IN44;
  output [44:0] Out1;
  output [31:0] Out2;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;
  wire w620;
  wire w622;
  wire w623;
  wire w624;
  wire w625;
  wire w626;
  wire w627;
  wire w628;
  wire w629;
  wire w630;
  wire w631;
  wire w632;
  wire w633;
  wire w634;
  wire w635;
  wire w636;
  wire w637;
  wire w638;
  wire w639;
  wire w640;
  wire w641;
  wire w642;
  wire w643;
  wire w644;
  wire w646;
  wire w647;
  wire w648;
  wire w649;
  wire w650;
  wire w651;
  wire w652;
  wire w653;
  wire w654;
  wire w655;
  wire w656;
  wire w657;
  wire w658;
  wire w659;
  wire w660;
  wire w661;
  wire w662;
  wire w663;
  wire w664;
  wire w665;
  wire w666;
  wire w667;
  wire w668;
  wire w670;
  wire w671;
  wire w672;
  wire w673;
  wire w674;
  wire w675;
  wire w676;
  wire w677;
  wire w678;
  wire w679;
  wire w680;
  wire w681;
  wire w682;
  wire w683;
  wire w684;
  wire w685;
  wire w686;
  wire w687;
  wire w688;
  wire w689;
  wire w690;
  wire w691;
  wire w692;
  wire w694;
  wire w695;
  wire w696;
  wire w697;
  wire w698;
  wire w699;
  wire w700;
  wire w701;
  wire w702;
  wire w703;
  wire w704;
  wire w705;
  wire w706;
  wire w707;
  wire w708;
  wire w709;
  wire w710;
  wire w711;
  wire w712;
  wire w713;
  wire w714;
  wire w715;
  wire w716;
  wire w718;
  wire w719;
  wire w720;
  wire w721;
  wire w722;
  wire w723;
  wire w724;
  wire w725;
  wire w726;
  wire w727;
  wire w728;
  wire w729;
  wire w730;
  wire w731;
  wire w732;
  wire w733;
  wire w734;
  wire w735;
  wire w736;
  wire w737;
  wire w738;
  wire w739;
  wire w740;
  wire w742;
  wire w743;
  wire w744;
  wire w745;
  wire w746;
  wire w747;
  wire w748;
  wire w749;
  wire w750;
  wire w751;
  wire w752;
  wire w753;
  wire w754;
  wire w755;
  wire w756;
  wire w757;
  wire w758;
  wire w759;
  wire w760;
  wire w761;
  wire w762;
  wire w763;
  wire w764;
  wire w766;
  wire w767;
  wire w768;
  wire w769;
  wire w770;
  wire w771;
  wire w772;
  wire w773;
  wire w774;
  wire w775;
  wire w776;
  wire w777;
  wire w778;
  wire w779;
  wire w780;
  wire w781;
  wire w782;
  wire w783;
  wire w784;
  wire w785;
  wire w786;
  wire w787;
  wire w788;
  wire w790;
  wire w791;
  wire w792;
  wire w793;
  wire w794;
  wire w795;
  wire w796;
  wire w797;
  wire w798;
  wire w799;
  wire w800;
  wire w801;
  wire w802;
  wire w803;
  wire w804;
  wire w805;
  wire w806;
  wire w807;
  wire w808;
  wire w809;
  wire w810;
  wire w811;
  wire w812;
  wire w814;
  wire w815;
  wire w816;
  wire w817;
  wire w818;
  wire w819;
  wire w820;
  wire w821;
  wire w822;
  wire w823;
  wire w824;
  wire w825;
  wire w826;
  wire w827;
  wire w828;
  wire w829;
  wire w830;
  wire w831;
  wire w832;
  wire w833;
  wire w834;
  wire w835;
  wire w836;
  wire w838;
  wire w839;
  wire w840;
  wire w841;
  wire w842;
  wire w843;
  wire w844;
  wire w845;
  wire w846;
  wire w847;
  wire w848;
  wire w849;
  wire w850;
  wire w851;
  wire w852;
  wire w853;
  wire w854;
  wire w855;
  wire w856;
  wire w857;
  wire w858;
  wire w859;
  wire w860;
  wire w862;
  wire w863;
  wire w864;
  wire w865;
  wire w866;
  wire w867;
  wire w868;
  wire w869;
  wire w870;
  wire w871;
  wire w872;
  wire w873;
  wire w874;
  wire w875;
  wire w876;
  wire w877;
  wire w878;
  wire w879;
  wire w880;
  wire w881;
  wire w882;
  wire w883;
  wire w884;
  wire w886;
  wire w887;
  wire w888;
  wire w889;
  wire w890;
  wire w891;
  wire w892;
  wire w893;
  wire w894;
  wire w895;
  wire w896;
  wire w897;
  wire w898;
  wire w899;
  wire w900;
  wire w901;
  wire w902;
  wire w903;
  wire w904;
  wire w905;
  wire w906;
  wire w907;
  wire w908;
  wire w910;
  wire w911;
  wire w912;
  wire w913;
  wire w914;
  wire w915;
  wire w916;
  wire w917;
  wire w918;
  wire w919;
  wire w920;
  wire w921;
  wire w922;
  wire w923;
  wire w924;
  wire w925;
  wire w926;
  wire w927;
  wire w928;
  wire w929;
  wire w930;
  wire w931;
  wire w932;
  wire w934;
  wire w935;
  wire w936;
  wire w937;
  wire w938;
  wire w939;
  wire w940;
  wire w941;
  wire w942;
  wire w943;
  wire w944;
  wire w945;
  wire w946;
  wire w947;
  wire w948;
  wire w949;
  wire w950;
  wire w951;
  wire w952;
  wire w953;
  wire w954;
  wire w955;
  wire w956;
  wire w958;
  wire w959;
  wire w960;
  wire w961;
  wire w962;
  wire w963;
  wire w964;
  wire w965;
  wire w966;
  wire w967;
  wire w968;
  wire w969;
  wire w970;
  wire w971;
  wire w972;
  wire w973;
  wire w974;
  wire w975;
  wire w976;
  wire w977;
  wire w978;
  wire w979;
  wire w980;
  wire w982;
  wire w983;
  wire w984;
  wire w985;
  wire w986;
  wire w987;
  wire w988;
  wire w989;
  wire w990;
  wire w991;
  wire w992;
  wire w993;
  wire w994;
  wire w995;
  wire w996;
  wire w997;
  wire w998;
  wire w999;
  wire w1000;
  wire w1001;
  wire w1002;
  wire w1003;
  wire w1004;
  wire w1006;
  wire w1007;
  wire w1008;
  wire w1009;
  wire w1010;
  wire w1011;
  wire w1012;
  wire w1013;
  wire w1014;
  wire w1015;
  wire w1016;
  wire w1017;
  wire w1018;
  wire w1019;
  wire w1020;
  wire w1021;
  wire w1022;
  wire w1023;
  wire w1024;
  wire w1025;
  wire w1026;
  wire w1027;
  wire w1028;
  wire w1030;
  wire w1031;
  wire w1032;
  wire w1033;
  wire w1034;
  wire w1035;
  wire w1036;
  wire w1037;
  wire w1038;
  wire w1039;
  wire w1040;
  wire w1041;
  wire w1042;
  wire w1043;
  wire w1044;
  wire w1045;
  wire w1046;
  wire w1047;
  wire w1048;
  wire w1049;
  wire w1050;
  wire w1051;
  wire w1052;
  wire w1054;
  wire w1055;
  wire w1056;
  wire w1057;
  wire w1058;
  wire w1059;
  wire w1060;
  wire w1061;
  wire w1062;
  wire w1063;
  wire w1064;
  wire w1065;
  wire w1066;
  wire w1067;
  wire w1068;
  wire w1069;
  wire w1070;
  wire w1071;
  wire w1072;
  wire w1073;
  wire w1074;
  wire w1075;
  wire w1076;
  wire w1078;
  wire w1079;
  wire w1080;
  wire w1081;
  wire w1082;
  wire w1083;
  wire w1084;
  wire w1085;
  wire w1086;
  wire w1087;
  wire w1088;
  wire w1089;
  wire w1090;
  wire w1091;
  wire w1092;
  wire w1093;
  wire w1094;
  wire w1095;
  wire w1096;
  wire w1097;
  wire w1098;
  wire w1099;
  wire w1100;
  wire w1102;
  wire w1103;
  wire w1104;
  wire w1105;
  wire w1106;
  wire w1107;
  wire w1108;
  wire w1109;
  wire w1110;
  wire w1111;
  wire w1112;
  wire w1113;
  wire w1114;
  wire w1115;
  wire w1116;
  wire w1117;
  wire w1118;
  wire w1119;
  wire w1120;
  wire w1121;
  wire w1122;
  wire w1123;
  wire w1124;
  wire w1126;
  wire w1127;
  wire w1128;
  wire w1129;
  wire w1130;
  wire w1131;
  wire w1132;
  wire w1133;
  wire w1134;
  wire w1135;
  wire w1136;
  wire w1137;
  wire w1138;
  wire w1139;
  wire w1140;
  wire w1141;
  wire w1142;
  wire w1143;
  wire w1144;
  wire w1145;
  wire w1146;
  wire w1147;
  wire w1148;
  wire w1150;
  wire w1151;
  wire w1152;
  wire w1153;
  wire w1154;
  wire w1155;
  wire w1156;
  wire w1157;
  wire w1158;
  wire w1159;
  wire w1160;
  wire w1161;
  wire w1162;
  wire w1163;
  wire w1164;
  wire w1165;
  wire w1166;
  wire w1167;
  wire w1168;
  wire w1169;
  wire w1170;
  wire w1171;
  wire w1172;
  wire w1174;
  wire w1176;
  wire w1178;
  wire w1180;
  wire w1182;
  wire w1184;
  wire w1186;
  wire w1188;
  wire w1190;
  wire w1192;
  wire w1194;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w430);
  FullAdder U1 (w430, IN2[0], IN2[1], w431, w432);
  FullAdder U2 (w432, IN3[0], IN3[1], w433, w434);
  FullAdder U3 (w434, IN4[0], IN4[1], w435, w436);
  FullAdder U4 (w436, IN5[0], IN5[1], w437, w438);
  FullAdder U5 (w438, IN6[0], IN6[1], w439, w440);
  FullAdder U6 (w440, IN7[0], IN7[1], w441, w442);
  FullAdder U7 (w442, IN8[0], IN8[1], w443, w444);
  FullAdder U8 (w444, IN9[0], IN9[1], w445, w446);
  FullAdder U9 (w446, IN10[0], IN10[1], w447, w448);
  FullAdder U10 (w448, IN11[0], IN11[1], w449, w450);
  FullAdder U11 (w450, IN12[0], IN12[1], w451, w452);
  HalfAdder U12 (w431, IN2[2], Out1[2], w454);
  FullAdder U13 (w454, w433, IN3[2], w455, w456);
  FullAdder U14 (w456, w435, IN4[2], w457, w458);
  FullAdder U15 (w458, w437, IN5[2], w459, w460);
  FullAdder U16 (w460, w439, IN6[2], w461, w462);
  FullAdder U17 (w462, w441, IN7[2], w463, w464);
  FullAdder U18 (w464, w443, IN8[2], w465, w466);
  FullAdder U19 (w466, w445, IN9[2], w467, w468);
  FullAdder U20 (w468, w447, IN10[2], w469, w470);
  FullAdder U21 (w470, w449, IN11[2], w471, w472);
  FullAdder U22 (w472, w451, IN12[2], w473, w474);
  FullAdder U23 (w474, w452, IN13[0], w475, w476);
  HalfAdder U24 (w455, IN3[3], Out1[3], w478);
  FullAdder U25 (w478, w457, IN4[3], w479, w480);
  FullAdder U26 (w480, w459, IN5[3], w481, w482);
  FullAdder U27 (w482, w461, IN6[3], w483, w484);
  FullAdder U28 (w484, w463, IN7[3], w485, w486);
  FullAdder U29 (w486, w465, IN8[3], w487, w488);
  FullAdder U30 (w488, w467, IN9[3], w489, w490);
  FullAdder U31 (w490, w469, IN10[3], w491, w492);
  FullAdder U32 (w492, w471, IN11[3], w493, w494);
  FullAdder U33 (w494, w473, IN12[3], w495, w496);
  FullAdder U34 (w496, w475, IN13[1], w497, w498);
  FullAdder U35 (w498, w476, IN14[0], w499, w500);
  HalfAdder U36 (w479, IN4[4], Out1[4], w502);
  FullAdder U37 (w502, w481, IN5[4], w503, w504);
  FullAdder U38 (w504, w483, IN6[4], w505, w506);
  FullAdder U39 (w506, w485, IN7[4], w507, w508);
  FullAdder U40 (w508, w487, IN8[4], w509, w510);
  FullAdder U41 (w510, w489, IN9[4], w511, w512);
  FullAdder U42 (w512, w491, IN10[4], w513, w514);
  FullAdder U43 (w514, w493, IN11[4], w515, w516);
  FullAdder U44 (w516, w495, IN12[4], w517, w518);
  FullAdder U45 (w518, w497, IN13[2], w519, w520);
  FullAdder U46 (w520, w499, IN14[1], w521, w522);
  FullAdder U47 (w522, w500, IN15[0], w523, w524);
  HalfAdder U48 (w503, IN5[5], Out1[5], w526);
  FullAdder U49 (w526, w505, IN6[5], w527, w528);
  FullAdder U50 (w528, w507, IN7[5], w529, w530);
  FullAdder U51 (w530, w509, IN8[5], w531, w532);
  FullAdder U52 (w532, w511, IN9[5], w533, w534);
  FullAdder U53 (w534, w513, IN10[5], w535, w536);
  FullAdder U54 (w536, w515, IN11[5], w537, w538);
  FullAdder U55 (w538, w517, IN12[5], w539, w540);
  FullAdder U56 (w540, w519, IN13[3], w541, w542);
  FullAdder U57 (w542, w521, IN14[2], w543, w544);
  FullAdder U58 (w544, w523, IN15[1], w545, w546);
  FullAdder U59 (w546, w524, IN16[0], w547, w548);
  HalfAdder U60 (w527, IN6[6], Out1[6], w550);
  FullAdder U61 (w550, w529, IN7[6], w551, w552);
  FullAdder U62 (w552, w531, IN8[6], w553, w554);
  FullAdder U63 (w554, w533, IN9[6], w555, w556);
  FullAdder U64 (w556, w535, IN10[6], w557, w558);
  FullAdder U65 (w558, w537, IN11[6], w559, w560);
  FullAdder U66 (w560, w539, IN12[6], w561, w562);
  FullAdder U67 (w562, w541, IN13[4], w563, w564);
  FullAdder U68 (w564, w543, IN14[3], w565, w566);
  FullAdder U69 (w566, w545, IN15[2], w567, w568);
  FullAdder U70 (w568, w547, IN16[1], w569, w570);
  FullAdder U71 (w570, w548, IN17[0], w571, w572);
  HalfAdder U72 (w551, IN7[7], Out1[7], w574);
  FullAdder U73 (w574, w553, IN8[7], w575, w576);
  FullAdder U74 (w576, w555, IN9[7], w577, w578);
  FullAdder U75 (w578, w557, IN10[7], w579, w580);
  FullAdder U76 (w580, w559, IN11[7], w581, w582);
  FullAdder U77 (w582, w561, IN12[7], w583, w584);
  FullAdder U78 (w584, w563, IN13[5], w585, w586);
  FullAdder U79 (w586, w565, IN14[4], w587, w588);
  FullAdder U80 (w588, w567, IN15[3], w589, w590);
  FullAdder U81 (w590, w569, IN16[2], w591, w592);
  FullAdder U82 (w592, w571, IN17[1], w593, w594);
  FullAdder U83 (w594, w572, IN18[0], w595, w596);
  HalfAdder U84 (w575, IN8[8], Out1[8], w598);
  FullAdder U85 (w598, w577, IN9[8], w599, w600);
  FullAdder U86 (w600, w579, IN10[8], w601, w602);
  FullAdder U87 (w602, w581, IN11[8], w603, w604);
  FullAdder U88 (w604, w583, IN12[8], w605, w606);
  FullAdder U89 (w606, w585, IN13[6], w607, w608);
  FullAdder U90 (w608, w587, IN14[5], w609, w610);
  FullAdder U91 (w610, w589, IN15[4], w611, w612);
  FullAdder U92 (w612, w591, IN16[3], w613, w614);
  FullAdder U93 (w614, w593, IN17[2], w615, w616);
  FullAdder U94 (w616, w595, IN18[1], w617, w618);
  FullAdder U95 (w618, w596, IN19[0], w619, w620);
  HalfAdder U96 (w599, IN9[9], Out1[9], w622);
  FullAdder U97 (w622, w601, IN10[9], w623, w624);
  FullAdder U98 (w624, w603, IN11[9], w625, w626);
  FullAdder U99 (w626, w605, IN12[9], w627, w628);
  FullAdder U100 (w628, w607, IN13[7], w629, w630);
  FullAdder U101 (w630, w609, IN14[6], w631, w632);
  FullAdder U102 (w632, w611, IN15[5], w633, w634);
  FullAdder U103 (w634, w613, IN16[4], w635, w636);
  FullAdder U104 (w636, w615, IN17[3], w637, w638);
  FullAdder U105 (w638, w617, IN18[2], w639, w640);
  FullAdder U106 (w640, w619, IN19[1], w641, w642);
  FullAdder U107 (w642, w620, IN20[0], w643, w644);
  HalfAdder U108 (w623, IN10[10], Out1[10], w646);
  FullAdder U109 (w646, w625, IN11[10], w647, w648);
  FullAdder U110 (w648, w627, IN12[10], w649, w650);
  FullAdder U111 (w650, w629, IN13[8], w651, w652);
  FullAdder U112 (w652, w631, IN14[7], w653, w654);
  FullAdder U113 (w654, w633, IN15[6], w655, w656);
  FullAdder U114 (w656, w635, IN16[5], w657, w658);
  FullAdder U115 (w658, w637, IN17[4], w659, w660);
  FullAdder U116 (w660, w639, IN18[3], w661, w662);
  FullAdder U117 (w662, w641, IN19[2], w663, w664);
  FullAdder U118 (w664, w643, IN20[1], w665, w666);
  FullAdder U119 (w666, w644, IN21[0], w667, w668);
  HalfAdder U120 (w647, IN11[11], Out1[11], w670);
  FullAdder U121 (w670, w649, IN12[11], w671, w672);
  FullAdder U122 (w672, w651, IN13[9], w673, w674);
  FullAdder U123 (w674, w653, IN14[8], w675, w676);
  FullAdder U124 (w676, w655, IN15[7], w677, w678);
  FullAdder U125 (w678, w657, IN16[6], w679, w680);
  FullAdder U126 (w680, w659, IN17[5], w681, w682);
  FullAdder U127 (w682, w661, IN18[4], w683, w684);
  FullAdder U128 (w684, w663, IN19[3], w685, w686);
  FullAdder U129 (w686, w665, IN20[2], w687, w688);
  FullAdder U130 (w688, w667, IN21[1], w689, w690);
  FullAdder U131 (w690, w668, IN22[0], w691, w692);
  HalfAdder U132 (w671, IN12[12], Out1[12], w694);
  FullAdder U133 (w694, w673, IN13[10], w695, w696);
  FullAdder U134 (w696, w675, IN14[9], w697, w698);
  FullAdder U135 (w698, w677, IN15[8], w699, w700);
  FullAdder U136 (w700, w679, IN16[7], w701, w702);
  FullAdder U137 (w702, w681, IN17[6], w703, w704);
  FullAdder U138 (w704, w683, IN18[5], w705, w706);
  FullAdder U139 (w706, w685, IN19[4], w707, w708);
  FullAdder U140 (w708, w687, IN20[3], w709, w710);
  FullAdder U141 (w710, w689, IN21[2], w711, w712);
  FullAdder U142 (w712, w691, IN22[1], w713, w714);
  FullAdder U143 (w714, w692, IN23[0], w715, w716);
  HalfAdder U144 (w695, IN13[11], Out1[13], w718);
  FullAdder U145 (w718, w697, IN14[10], w719, w720);
  FullAdder U146 (w720, w699, IN15[9], w721, w722);
  FullAdder U147 (w722, w701, IN16[8], w723, w724);
  FullAdder U148 (w724, w703, IN17[7], w725, w726);
  FullAdder U149 (w726, w705, IN18[6], w727, w728);
  FullAdder U150 (w728, w707, IN19[5], w729, w730);
  FullAdder U151 (w730, w709, IN20[4], w731, w732);
  FullAdder U152 (w732, w711, IN21[3], w733, w734);
  FullAdder U153 (w734, w713, IN22[2], w735, w736);
  FullAdder U154 (w736, w715, IN23[1], w737, w738);
  FullAdder U155 (w738, w716, IN24[0], w739, w740);
  HalfAdder U156 (w719, IN14[11], Out1[14], w742);
  FullAdder U157 (w742, w721, IN15[10], w743, w744);
  FullAdder U158 (w744, w723, IN16[9], w745, w746);
  FullAdder U159 (w746, w725, IN17[8], w747, w748);
  FullAdder U160 (w748, w727, IN18[7], w749, w750);
  FullAdder U161 (w750, w729, IN19[6], w751, w752);
  FullAdder U162 (w752, w731, IN20[5], w753, w754);
  FullAdder U163 (w754, w733, IN21[4], w755, w756);
  FullAdder U164 (w756, w735, IN22[3], w757, w758);
  FullAdder U165 (w758, w737, IN23[2], w759, w760);
  FullAdder U166 (w760, w739, IN24[1], w761, w762);
  FullAdder U167 (w762, w740, IN25[0], w763, w764);
  HalfAdder U168 (w743, IN15[11], Out1[15], w766);
  FullAdder U169 (w766, w745, IN16[10], w767, w768);
  FullAdder U170 (w768, w747, IN17[9], w769, w770);
  FullAdder U171 (w770, w749, IN18[8], w771, w772);
  FullAdder U172 (w772, w751, IN19[7], w773, w774);
  FullAdder U173 (w774, w753, IN20[6], w775, w776);
  FullAdder U174 (w776, w755, IN21[5], w777, w778);
  FullAdder U175 (w778, w757, IN22[4], w779, w780);
  FullAdder U176 (w780, w759, IN23[3], w781, w782);
  FullAdder U177 (w782, w761, IN24[2], w783, w784);
  FullAdder U178 (w784, w763, IN25[1], w785, w786);
  FullAdder U179 (w786, w764, IN26[0], w787, w788);
  HalfAdder U180 (w767, IN16[11], Out1[16], w790);
  FullAdder U181 (w790, w769, IN17[10], w791, w792);
  FullAdder U182 (w792, w771, IN18[9], w793, w794);
  FullAdder U183 (w794, w773, IN19[8], w795, w796);
  FullAdder U184 (w796, w775, IN20[7], w797, w798);
  FullAdder U185 (w798, w777, IN21[6], w799, w800);
  FullAdder U186 (w800, w779, IN22[5], w801, w802);
  FullAdder U187 (w802, w781, IN23[4], w803, w804);
  FullAdder U188 (w804, w783, IN24[3], w805, w806);
  FullAdder U189 (w806, w785, IN25[2], w807, w808);
  FullAdder U190 (w808, w787, IN26[1], w809, w810);
  FullAdder U191 (w810, w788, IN27[0], w811, w812);
  HalfAdder U192 (w791, IN17[11], Out1[17], w814);
  FullAdder U193 (w814, w793, IN18[10], w815, w816);
  FullAdder U194 (w816, w795, IN19[9], w817, w818);
  FullAdder U195 (w818, w797, IN20[8], w819, w820);
  FullAdder U196 (w820, w799, IN21[7], w821, w822);
  FullAdder U197 (w822, w801, IN22[6], w823, w824);
  FullAdder U198 (w824, w803, IN23[5], w825, w826);
  FullAdder U199 (w826, w805, IN24[4], w827, w828);
  FullAdder U200 (w828, w807, IN25[3], w829, w830);
  FullAdder U201 (w830, w809, IN26[2], w831, w832);
  FullAdder U202 (w832, w811, IN27[1], w833, w834);
  FullAdder U203 (w834, w812, IN28[0], w835, w836);
  HalfAdder U204 (w815, IN18[11], Out1[18], w838);
  FullAdder U205 (w838, w817, IN19[10], w839, w840);
  FullAdder U206 (w840, w819, IN20[9], w841, w842);
  FullAdder U207 (w842, w821, IN21[8], w843, w844);
  FullAdder U208 (w844, w823, IN22[7], w845, w846);
  FullAdder U209 (w846, w825, IN23[6], w847, w848);
  FullAdder U210 (w848, w827, IN24[5], w849, w850);
  FullAdder U211 (w850, w829, IN25[4], w851, w852);
  FullAdder U212 (w852, w831, IN26[3], w853, w854);
  FullAdder U213 (w854, w833, IN27[2], w855, w856);
  FullAdder U214 (w856, w835, IN28[1], w857, w858);
  FullAdder U215 (w858, w836, IN29[0], w859, w860);
  HalfAdder U216 (w839, IN19[11], Out1[19], w862);
  FullAdder U217 (w862, w841, IN20[10], w863, w864);
  FullAdder U218 (w864, w843, IN21[9], w865, w866);
  FullAdder U219 (w866, w845, IN22[8], w867, w868);
  FullAdder U220 (w868, w847, IN23[7], w869, w870);
  FullAdder U221 (w870, w849, IN24[6], w871, w872);
  FullAdder U222 (w872, w851, IN25[5], w873, w874);
  FullAdder U223 (w874, w853, IN26[4], w875, w876);
  FullAdder U224 (w876, w855, IN27[3], w877, w878);
  FullAdder U225 (w878, w857, IN28[2], w879, w880);
  FullAdder U226 (w880, w859, IN29[1], w881, w882);
  FullAdder U227 (w882, w860, IN30[0], w883, w884);
  HalfAdder U228 (w863, IN20[11], Out1[20], w886);
  FullAdder U229 (w886, w865, IN21[10], w887, w888);
  FullAdder U230 (w888, w867, IN22[9], w889, w890);
  FullAdder U231 (w890, w869, IN23[8], w891, w892);
  FullAdder U232 (w892, w871, IN24[7], w893, w894);
  FullAdder U233 (w894, w873, IN25[6], w895, w896);
  FullAdder U234 (w896, w875, IN26[5], w897, w898);
  FullAdder U235 (w898, w877, IN27[4], w899, w900);
  FullAdder U236 (w900, w879, IN28[3], w901, w902);
  FullAdder U237 (w902, w881, IN29[2], w903, w904);
  FullAdder U238 (w904, w883, IN30[1], w905, w906);
  FullAdder U239 (w906, w884, IN31[0], w907, w908);
  HalfAdder U240 (w887, IN21[11], Out1[21], w910);
  FullAdder U241 (w910, w889, IN22[10], w911, w912);
  FullAdder U242 (w912, w891, IN23[9], w913, w914);
  FullAdder U243 (w914, w893, IN24[8], w915, w916);
  FullAdder U244 (w916, w895, IN25[7], w917, w918);
  FullAdder U245 (w918, w897, IN26[6], w919, w920);
  FullAdder U246 (w920, w899, IN27[5], w921, w922);
  FullAdder U247 (w922, w901, IN28[4], w923, w924);
  FullAdder U248 (w924, w903, IN29[3], w925, w926);
  FullAdder U249 (w926, w905, IN30[2], w927, w928);
  FullAdder U250 (w928, w907, IN31[1], w929, w930);
  FullAdder U251 (w930, w908, IN32[0], w931, w932);
  HalfAdder U252 (w911, IN22[11], Out1[22], w934);
  FullAdder U253 (w934, w913, IN23[10], w935, w936);
  FullAdder U254 (w936, w915, IN24[9], w937, w938);
  FullAdder U255 (w938, w917, IN25[8], w939, w940);
  FullAdder U256 (w940, w919, IN26[7], w941, w942);
  FullAdder U257 (w942, w921, IN27[6], w943, w944);
  FullAdder U258 (w944, w923, IN28[5], w945, w946);
  FullAdder U259 (w946, w925, IN29[4], w947, w948);
  FullAdder U260 (w948, w927, IN30[3], w949, w950);
  FullAdder U261 (w950, w929, IN31[2], w951, w952);
  FullAdder U262 (w952, w931, IN32[1], w953, w954);
  FullAdder U263 (w954, w932, IN33[0], w955, w956);
  HalfAdder U264 (w935, IN23[11], Out1[23], w958);
  FullAdder U265 (w958, w937, IN24[10], w959, w960);
  FullAdder U266 (w960, w939, IN25[9], w961, w962);
  FullAdder U267 (w962, w941, IN26[8], w963, w964);
  FullAdder U268 (w964, w943, IN27[7], w965, w966);
  FullAdder U269 (w966, w945, IN28[6], w967, w968);
  FullAdder U270 (w968, w947, IN29[5], w969, w970);
  FullAdder U271 (w970, w949, IN30[4], w971, w972);
  FullAdder U272 (w972, w951, IN31[3], w973, w974);
  FullAdder U273 (w974, w953, IN32[2], w975, w976);
  FullAdder U274 (w976, w955, IN33[1], w977, w978);
  FullAdder U275 (w978, w956, IN34[0], w979, w980);
  HalfAdder U276 (w959, IN24[11], Out1[24], w982);
  FullAdder U277 (w982, w961, IN25[10], w983, w984);
  FullAdder U278 (w984, w963, IN26[9], w985, w986);
  FullAdder U279 (w986, w965, IN27[8], w987, w988);
  FullAdder U280 (w988, w967, IN28[7], w989, w990);
  FullAdder U281 (w990, w969, IN29[6], w991, w992);
  FullAdder U282 (w992, w971, IN30[5], w993, w994);
  FullAdder U283 (w994, w973, IN31[4], w995, w996);
  FullAdder U284 (w996, w975, IN32[3], w997, w998);
  FullAdder U285 (w998, w977, IN33[2], w999, w1000);
  FullAdder U286 (w1000, w979, IN34[1], w1001, w1002);
  FullAdder U287 (w1002, w980, IN35[0], w1003, w1004);
  HalfAdder U288 (w983, IN25[11], Out1[25], w1006);
  FullAdder U289 (w1006, w985, IN26[10], w1007, w1008);
  FullAdder U290 (w1008, w987, IN27[9], w1009, w1010);
  FullAdder U291 (w1010, w989, IN28[8], w1011, w1012);
  FullAdder U292 (w1012, w991, IN29[7], w1013, w1014);
  FullAdder U293 (w1014, w993, IN30[6], w1015, w1016);
  FullAdder U294 (w1016, w995, IN31[5], w1017, w1018);
  FullAdder U295 (w1018, w997, IN32[4], w1019, w1020);
  FullAdder U296 (w1020, w999, IN33[3], w1021, w1022);
  FullAdder U297 (w1022, w1001, IN34[2], w1023, w1024);
  FullAdder U298 (w1024, w1003, IN35[1], w1025, w1026);
  FullAdder U299 (w1026, w1004, IN36[0], w1027, w1028);
  HalfAdder U300 (w1007, IN26[11], Out1[26], w1030);
  FullAdder U301 (w1030, w1009, IN27[10], w1031, w1032);
  FullAdder U302 (w1032, w1011, IN28[9], w1033, w1034);
  FullAdder U303 (w1034, w1013, IN29[8], w1035, w1036);
  FullAdder U304 (w1036, w1015, IN30[7], w1037, w1038);
  FullAdder U305 (w1038, w1017, IN31[6], w1039, w1040);
  FullAdder U306 (w1040, w1019, IN32[5], w1041, w1042);
  FullAdder U307 (w1042, w1021, IN33[4], w1043, w1044);
  FullAdder U308 (w1044, w1023, IN34[3], w1045, w1046);
  FullAdder U309 (w1046, w1025, IN35[2], w1047, w1048);
  FullAdder U310 (w1048, w1027, IN36[1], w1049, w1050);
  FullAdder U311 (w1050, w1028, IN37[0], w1051, w1052);
  HalfAdder U312 (w1031, IN27[11], Out1[27], w1054);
  FullAdder U313 (w1054, w1033, IN28[10], w1055, w1056);
  FullAdder U314 (w1056, w1035, IN29[9], w1057, w1058);
  FullAdder U315 (w1058, w1037, IN30[8], w1059, w1060);
  FullAdder U316 (w1060, w1039, IN31[7], w1061, w1062);
  FullAdder U317 (w1062, w1041, IN32[6], w1063, w1064);
  FullAdder U318 (w1064, w1043, IN33[5], w1065, w1066);
  FullAdder U319 (w1066, w1045, IN34[4], w1067, w1068);
  FullAdder U320 (w1068, w1047, IN35[3], w1069, w1070);
  FullAdder U321 (w1070, w1049, IN36[2], w1071, w1072);
  FullAdder U322 (w1072, w1051, IN37[1], w1073, w1074);
  FullAdder U323 (w1074, w1052, IN38[0], w1075, w1076);
  HalfAdder U324 (w1055, IN28[11], Out1[28], w1078);
  FullAdder U325 (w1078, w1057, IN29[10], w1079, w1080);
  FullAdder U326 (w1080, w1059, IN30[9], w1081, w1082);
  FullAdder U327 (w1082, w1061, IN31[8], w1083, w1084);
  FullAdder U328 (w1084, w1063, IN32[7], w1085, w1086);
  FullAdder U329 (w1086, w1065, IN33[6], w1087, w1088);
  FullAdder U330 (w1088, w1067, IN34[5], w1089, w1090);
  FullAdder U331 (w1090, w1069, IN35[4], w1091, w1092);
  FullAdder U332 (w1092, w1071, IN36[3], w1093, w1094);
  FullAdder U333 (w1094, w1073, IN37[2], w1095, w1096);
  FullAdder U334 (w1096, w1075, IN38[1], w1097, w1098);
  FullAdder U335 (w1098, w1076, IN39[0], w1099, w1100);
  HalfAdder U336 (w1079, IN29[11], Out1[29], w1102);
  FullAdder U337 (w1102, w1081, IN30[10], w1103, w1104);
  FullAdder U338 (w1104, w1083, IN31[9], w1105, w1106);
  FullAdder U339 (w1106, w1085, IN32[8], w1107, w1108);
  FullAdder U340 (w1108, w1087, IN33[7], w1109, w1110);
  FullAdder U341 (w1110, w1089, IN34[6], w1111, w1112);
  FullAdder U342 (w1112, w1091, IN35[5], w1113, w1114);
  FullAdder U343 (w1114, w1093, IN36[4], w1115, w1116);
  FullAdder U344 (w1116, w1095, IN37[3], w1117, w1118);
  FullAdder U345 (w1118, w1097, IN38[2], w1119, w1120);
  FullAdder U346 (w1120, w1099, IN39[1], w1121, w1122);
  FullAdder U347 (w1122, w1100, IN40[0], w1123, w1124);
  HalfAdder U348 (w1103, IN30[11], Out1[30], w1126);
  FullAdder U349 (w1126, w1105, IN31[10], w1127, w1128);
  FullAdder U350 (w1128, w1107, IN32[9], w1129, w1130);
  FullAdder U351 (w1130, w1109, IN33[8], w1131, w1132);
  FullAdder U352 (w1132, w1111, IN34[7], w1133, w1134);
  FullAdder U353 (w1134, w1113, IN35[6], w1135, w1136);
  FullAdder U354 (w1136, w1115, IN36[5], w1137, w1138);
  FullAdder U355 (w1138, w1117, IN37[4], w1139, w1140);
  FullAdder U356 (w1140, w1119, IN38[3], w1141, w1142);
  FullAdder U357 (w1142, w1121, IN39[2], w1143, w1144);
  FullAdder U358 (w1144, w1123, IN40[1], w1145, w1146);
  FullAdder U359 (w1146, w1124, IN41[0], w1147, w1148);
  HalfAdder U360 (w1127, IN31[11], Out1[31], w1150);
  FullAdder U361 (w1150, w1129, IN32[10], w1151, w1152);
  FullAdder U362 (w1152, w1131, IN33[9], w1153, w1154);
  FullAdder U363 (w1154, w1133, IN34[8], w1155, w1156);
  FullAdder U364 (w1156, w1135, IN35[7], w1157, w1158);
  FullAdder U365 (w1158, w1137, IN36[6], w1159, w1160);
  FullAdder U366 (w1160, w1139, IN37[5], w1161, w1162);
  FullAdder U367 (w1162, w1141, IN38[4], w1163, w1164);
  FullAdder U368 (w1164, w1143, IN39[3], w1165, w1166);
  FullAdder U369 (w1166, w1145, IN40[2], w1167, w1168);
  FullAdder U370 (w1168, w1147, IN41[1], w1169, w1170);
  FullAdder U371 (w1170, w1148, IN42[0], w1171, w1172);
  HalfAdder U372 (w1151, IN32[11], Out1[32], w1174);
  FullAdder U373 (w1174, w1153, IN33[10], Out1[33], w1176);
  FullAdder U374 (w1176, w1155, IN34[9], Out1[34], w1178);
  FullAdder U375 (w1178, w1157, IN35[8], Out1[35], w1180);
  FullAdder U376 (w1180, w1159, IN36[7], Out1[36], w1182);
  FullAdder U377 (w1182, w1161, IN37[6], Out1[37], w1184);
  FullAdder U378 (w1184, w1163, IN38[5], Out1[38], w1186);
  FullAdder U379 (w1186, w1165, IN39[4], Out1[39], w1188);
  FullAdder U380 (w1188, w1167, IN40[3], Out1[40], w1190);
  FullAdder U381 (w1190, w1169, IN41[2], Out1[41], w1192);
  FullAdder U382 (w1192, w1171, IN42[1], Out1[42], w1194);
  FullAdder U383 (w1194, w1172, IN43[0], Out1[43], Out1[44]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN13[12];
  assign Out2[1] = IN14[12];
  assign Out2[2] = IN15[12];
  assign Out2[3] = IN16[12];
  assign Out2[4] = IN17[12];
  assign Out2[5] = IN18[12];
  assign Out2[6] = IN19[12];
  assign Out2[7] = IN20[12];
  assign Out2[8] = IN21[12];
  assign Out2[9] = IN22[12];
  assign Out2[10] = IN23[12];
  assign Out2[11] = IN24[12];
  assign Out2[12] = IN25[12];
  assign Out2[13] = IN26[12];
  assign Out2[14] = IN27[12];
  assign Out2[15] = IN28[12];
  assign Out2[16] = IN29[12];
  assign Out2[17] = IN30[12];
  assign Out2[18] = IN31[12];
  assign Out2[19] = IN32[12];
  assign Out2[20] = IN33[11];
  assign Out2[21] = IN34[10];
  assign Out2[22] = IN35[9];
  assign Out2[23] = IN36[8];
  assign Out2[24] = IN37[7];
  assign Out2[25] = IN38[6];
  assign Out2[26] = IN39[5];
  assign Out2[27] = IN40[4];
  assign Out2[28] = IN41[3];
  assign Out2[29] = IN42[2];
  assign Out2[30] = IN43[1];
  assign Out2[31] = IN44[0];

endmodule
module RC_32_32(IN1, IN2, Out);
  input [31:0] IN1;
  input [31:0] IN2;
  output [32:0] Out;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w65);
  FullAdder U1 (IN1[1], IN2[1], w65, Out[1], w67);
  FullAdder U2 (IN1[2], IN2[2], w67, Out[2], w69);
  FullAdder U3 (IN1[3], IN2[3], w69, Out[3], w71);
  FullAdder U4 (IN1[4], IN2[4], w71, Out[4], w73);
  FullAdder U5 (IN1[5], IN2[5], w73, Out[5], w75);
  FullAdder U6 (IN1[6], IN2[6], w75, Out[6], w77);
  FullAdder U7 (IN1[7], IN2[7], w77, Out[7], w79);
  FullAdder U8 (IN1[8], IN2[8], w79, Out[8], w81);
  FullAdder U9 (IN1[9], IN2[9], w81, Out[9], w83);
  FullAdder U10 (IN1[10], IN2[10], w83, Out[10], w85);
  FullAdder U11 (IN1[11], IN2[11], w85, Out[11], w87);
  FullAdder U12 (IN1[12], IN2[12], w87, Out[12], w89);
  FullAdder U13 (IN1[13], IN2[13], w89, Out[13], w91);
  FullAdder U14 (IN1[14], IN2[14], w91, Out[14], w93);
  FullAdder U15 (IN1[15], IN2[15], w93, Out[15], w95);
  FullAdder U16 (IN1[16], IN2[16], w95, Out[16], w97);
  FullAdder U17 (IN1[17], IN2[17], w97, Out[17], w99);
  FullAdder U18 (IN1[18], IN2[18], w99, Out[18], w101);
  FullAdder U19 (IN1[19], IN2[19], w101, Out[19], w103);
  FullAdder U20 (IN1[20], IN2[20], w103, Out[20], w105);
  FullAdder U21 (IN1[21], IN2[21], w105, Out[21], w107);
  FullAdder U22 (IN1[22], IN2[22], w107, Out[22], w109);
  FullAdder U23 (IN1[23], IN2[23], w109, Out[23], w111);
  FullAdder U24 (IN1[24], IN2[24], w111, Out[24], w113);
  FullAdder U25 (IN1[25], IN2[25], w113, Out[25], w115);
  FullAdder U26 (IN1[26], IN2[26], w115, Out[26], w117);
  FullAdder U27 (IN1[27], IN2[27], w117, Out[27], w119);
  FullAdder U28 (IN1[28], IN2[28], w119, Out[28], w121);
  FullAdder U29 (IN1[29], IN2[29], w121, Out[29], w123);
  FullAdder U30 (IN1[30], IN2[30], w123, Out[30], w125);
  FullAdder U31 (IN1[31], IN2[31], w125, Out[31], Out[32]);

endmodule
module NR_13_33(IN1, IN2, Out);
  input [12:0] IN1;
  input [32:0] IN2;
  output [45:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [12:0] P13;
  wire [12:0] P14;
  wire [12:0] P15;
  wire [12:0] P16;
  wire [12:0] P17;
  wire [12:0] P18;
  wire [12:0] P19;
  wire [12:0] P20;
  wire [12:0] P21;
  wire [12:0] P22;
  wire [12:0] P23;
  wire [12:0] P24;
  wire [12:0] P25;
  wire [12:0] P26;
  wire [12:0] P27;
  wire [12:0] P28;
  wire [12:0] P29;
  wire [12:0] P30;
  wire [12:0] P31;
  wire [12:0] P32;
  wire [11:0] P33;
  wire [10:0] P34;
  wire [9:0] P35;
  wire [8:0] P36;
  wire [7:0] P37;
  wire [6:0] P38;
  wire [5:0] P39;
  wire [4:0] P40;
  wire [3:0] P41;
  wire [2:0] P42;
  wire [1:0] P43;
  wire [0:0] P44;
  wire [44:0] R1;
  wire [31:0] R2;
  wire [45:0] aOut;
  U_SP_13_33 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, R1, R2);
  RC_32_32 S2 (R1[44:13], R2, aOut[45:13]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign Out = aOut[45:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
