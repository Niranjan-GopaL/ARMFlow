
module customAdder42_0(
    input [41 : 0] A,
    input [41 : 0] B,
    output [42 : 0] Sum
);

    assign Sum = A+B;

endmodule
