//Compilation time: 2025-03-17 16:17:21
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 41
  second input length: 54
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Array [AR]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule
module FullAdderProp(X, Y, Z, S, C, P);
  output C;
  output S;
  output P;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
  assign P = X ^ Y;
endmodule
module HalfAdder(X, Y, S, C);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule
module ConstatntOne(O);
  output O;
  assign O = 1;
endmodule
module Counter(X1, X2, X3, X4, X5, X6, X7, S3, S2, S1);
output S1;
output S2;
output S3;
input X1;
input X2;
input X3;
input X4;
input X5;
input X6;
input X7;
wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
assign W1 = X1 ^ X2 ^ X3;
assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
assign W5 = ~ ( X4 & X5 & X6 & X7 );
assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
assign S3 = W1 ^ W2;
assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule
module U_SP_41_54(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93);
  input [40:0] IN1;
  input [53:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [16:0] P16;
  output [17:0] P17;
  output [18:0] P18;
  output [19:0] P19;
  output [20:0] P20;
  output [21:0] P21;
  output [22:0] P22;
  output [23:0] P23;
  output [24:0] P24;
  output [25:0] P25;
  output [26:0] P26;
  output [27:0] P27;
  output [28:0] P28;
  output [29:0] P29;
  output [30:0] P30;
  output [31:0] P31;
  output [32:0] P32;
  output [33:0] P33;
  output [34:0] P34;
  output [35:0] P35;
  output [36:0] P36;
  output [37:0] P37;
  output [38:0] P38;
  output [39:0] P39;
  output [40:0] P40;
  output [40:0] P41;
  output [40:0] P42;
  output [40:0] P43;
  output [40:0] P44;
  output [40:0] P45;
  output [40:0] P46;
  output [40:0] P47;
  output [40:0] P48;
  output [40:0] P49;
  output [40:0] P50;
  output [40:0] P51;
  output [40:0] P52;
  output [40:0] P53;
  output [39:0] P54;
  output [38:0] P55;
  output [37:0] P56;
  output [36:0] P57;
  output [35:0] P58;
  output [34:0] P59;
  output [33:0] P60;
  output [32:0] P61;
  output [31:0] P62;
  output [30:0] P63;
  output [29:0] P64;
  output [28:0] P65;
  output [27:0] P66;
  output [26:0] P67;
  output [25:0] P68;
  output [24:0] P69;
  output [23:0] P70;
  output [22:0] P71;
  output [21:0] P72;
  output [20:0] P73;
  output [19:0] P74;
  output [18:0] P75;
  output [17:0] P76;
  output [16:0] P77;
  output [15:0] P78;
  output [14:0] P79;
  output [13:0] P80;
  output [12:0] P81;
  output [11:0] P82;
  output [10:0] P83;
  output [9:0] P84;
  output [8:0] P85;
  output [7:0] P86;
  output [6:0] P87;
  output [5:0] P88;
  output [4:0] P89;
  output [3:0] P90;
  output [2:0] P91;
  output [1:0] P92;
  output [0:0] P93;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P16[0] = IN1[0]&IN2[16];
  assign P17[0] = IN1[0]&IN2[17];
  assign P18[0] = IN1[0]&IN2[18];
  assign P19[0] = IN1[0]&IN2[19];
  assign P20[0] = IN1[0]&IN2[20];
  assign P21[0] = IN1[0]&IN2[21];
  assign P22[0] = IN1[0]&IN2[22];
  assign P23[0] = IN1[0]&IN2[23];
  assign P24[0] = IN1[0]&IN2[24];
  assign P25[0] = IN1[0]&IN2[25];
  assign P26[0] = IN1[0]&IN2[26];
  assign P27[0] = IN1[0]&IN2[27];
  assign P28[0] = IN1[0]&IN2[28];
  assign P29[0] = IN1[0]&IN2[29];
  assign P30[0] = IN1[0]&IN2[30];
  assign P31[0] = IN1[0]&IN2[31];
  assign P32[0] = IN1[0]&IN2[32];
  assign P33[0] = IN1[0]&IN2[33];
  assign P34[0] = IN1[0]&IN2[34];
  assign P35[0] = IN1[0]&IN2[35];
  assign P36[0] = IN1[0]&IN2[36];
  assign P37[0] = IN1[0]&IN2[37];
  assign P38[0] = IN1[0]&IN2[38];
  assign P39[0] = IN1[0]&IN2[39];
  assign P40[0] = IN1[0]&IN2[40];
  assign P41[0] = IN1[0]&IN2[41];
  assign P42[0] = IN1[0]&IN2[42];
  assign P43[0] = IN1[0]&IN2[43];
  assign P44[0] = IN1[0]&IN2[44];
  assign P45[0] = IN1[0]&IN2[45];
  assign P46[0] = IN1[0]&IN2[46];
  assign P47[0] = IN1[0]&IN2[47];
  assign P48[0] = IN1[0]&IN2[48];
  assign P49[0] = IN1[0]&IN2[49];
  assign P50[0] = IN1[0]&IN2[50];
  assign P51[0] = IN1[0]&IN2[51];
  assign P52[0] = IN1[0]&IN2[52];
  assign P53[0] = IN1[0]&IN2[53];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[1] = IN1[1]&IN2[15];
  assign P17[1] = IN1[1]&IN2[16];
  assign P18[1] = IN1[1]&IN2[17];
  assign P19[1] = IN1[1]&IN2[18];
  assign P20[1] = IN1[1]&IN2[19];
  assign P21[1] = IN1[1]&IN2[20];
  assign P22[1] = IN1[1]&IN2[21];
  assign P23[1] = IN1[1]&IN2[22];
  assign P24[1] = IN1[1]&IN2[23];
  assign P25[1] = IN1[1]&IN2[24];
  assign P26[1] = IN1[1]&IN2[25];
  assign P27[1] = IN1[1]&IN2[26];
  assign P28[1] = IN1[1]&IN2[27];
  assign P29[1] = IN1[1]&IN2[28];
  assign P30[1] = IN1[1]&IN2[29];
  assign P31[1] = IN1[1]&IN2[30];
  assign P32[1] = IN1[1]&IN2[31];
  assign P33[1] = IN1[1]&IN2[32];
  assign P34[1] = IN1[1]&IN2[33];
  assign P35[1] = IN1[1]&IN2[34];
  assign P36[1] = IN1[1]&IN2[35];
  assign P37[1] = IN1[1]&IN2[36];
  assign P38[1] = IN1[1]&IN2[37];
  assign P39[1] = IN1[1]&IN2[38];
  assign P40[1] = IN1[1]&IN2[39];
  assign P41[1] = IN1[1]&IN2[40];
  assign P42[1] = IN1[1]&IN2[41];
  assign P43[1] = IN1[1]&IN2[42];
  assign P44[1] = IN1[1]&IN2[43];
  assign P45[1] = IN1[1]&IN2[44];
  assign P46[1] = IN1[1]&IN2[45];
  assign P47[1] = IN1[1]&IN2[46];
  assign P48[1] = IN1[1]&IN2[47];
  assign P49[1] = IN1[1]&IN2[48];
  assign P50[1] = IN1[1]&IN2[49];
  assign P51[1] = IN1[1]&IN2[50];
  assign P52[1] = IN1[1]&IN2[51];
  assign P53[1] = IN1[1]&IN2[52];
  assign P54[0] = IN1[1]&IN2[53];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[2] = IN1[2]&IN2[14];
  assign P17[2] = IN1[2]&IN2[15];
  assign P18[2] = IN1[2]&IN2[16];
  assign P19[2] = IN1[2]&IN2[17];
  assign P20[2] = IN1[2]&IN2[18];
  assign P21[2] = IN1[2]&IN2[19];
  assign P22[2] = IN1[2]&IN2[20];
  assign P23[2] = IN1[2]&IN2[21];
  assign P24[2] = IN1[2]&IN2[22];
  assign P25[2] = IN1[2]&IN2[23];
  assign P26[2] = IN1[2]&IN2[24];
  assign P27[2] = IN1[2]&IN2[25];
  assign P28[2] = IN1[2]&IN2[26];
  assign P29[2] = IN1[2]&IN2[27];
  assign P30[2] = IN1[2]&IN2[28];
  assign P31[2] = IN1[2]&IN2[29];
  assign P32[2] = IN1[2]&IN2[30];
  assign P33[2] = IN1[2]&IN2[31];
  assign P34[2] = IN1[2]&IN2[32];
  assign P35[2] = IN1[2]&IN2[33];
  assign P36[2] = IN1[2]&IN2[34];
  assign P37[2] = IN1[2]&IN2[35];
  assign P38[2] = IN1[2]&IN2[36];
  assign P39[2] = IN1[2]&IN2[37];
  assign P40[2] = IN1[2]&IN2[38];
  assign P41[2] = IN1[2]&IN2[39];
  assign P42[2] = IN1[2]&IN2[40];
  assign P43[2] = IN1[2]&IN2[41];
  assign P44[2] = IN1[2]&IN2[42];
  assign P45[2] = IN1[2]&IN2[43];
  assign P46[2] = IN1[2]&IN2[44];
  assign P47[2] = IN1[2]&IN2[45];
  assign P48[2] = IN1[2]&IN2[46];
  assign P49[2] = IN1[2]&IN2[47];
  assign P50[2] = IN1[2]&IN2[48];
  assign P51[2] = IN1[2]&IN2[49];
  assign P52[2] = IN1[2]&IN2[50];
  assign P53[2] = IN1[2]&IN2[51];
  assign P54[1] = IN1[2]&IN2[52];
  assign P55[0] = IN1[2]&IN2[53];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[3] = IN1[3]&IN2[13];
  assign P17[3] = IN1[3]&IN2[14];
  assign P18[3] = IN1[3]&IN2[15];
  assign P19[3] = IN1[3]&IN2[16];
  assign P20[3] = IN1[3]&IN2[17];
  assign P21[3] = IN1[3]&IN2[18];
  assign P22[3] = IN1[3]&IN2[19];
  assign P23[3] = IN1[3]&IN2[20];
  assign P24[3] = IN1[3]&IN2[21];
  assign P25[3] = IN1[3]&IN2[22];
  assign P26[3] = IN1[3]&IN2[23];
  assign P27[3] = IN1[3]&IN2[24];
  assign P28[3] = IN1[3]&IN2[25];
  assign P29[3] = IN1[3]&IN2[26];
  assign P30[3] = IN1[3]&IN2[27];
  assign P31[3] = IN1[3]&IN2[28];
  assign P32[3] = IN1[3]&IN2[29];
  assign P33[3] = IN1[3]&IN2[30];
  assign P34[3] = IN1[3]&IN2[31];
  assign P35[3] = IN1[3]&IN2[32];
  assign P36[3] = IN1[3]&IN2[33];
  assign P37[3] = IN1[3]&IN2[34];
  assign P38[3] = IN1[3]&IN2[35];
  assign P39[3] = IN1[3]&IN2[36];
  assign P40[3] = IN1[3]&IN2[37];
  assign P41[3] = IN1[3]&IN2[38];
  assign P42[3] = IN1[3]&IN2[39];
  assign P43[3] = IN1[3]&IN2[40];
  assign P44[3] = IN1[3]&IN2[41];
  assign P45[3] = IN1[3]&IN2[42];
  assign P46[3] = IN1[3]&IN2[43];
  assign P47[3] = IN1[3]&IN2[44];
  assign P48[3] = IN1[3]&IN2[45];
  assign P49[3] = IN1[3]&IN2[46];
  assign P50[3] = IN1[3]&IN2[47];
  assign P51[3] = IN1[3]&IN2[48];
  assign P52[3] = IN1[3]&IN2[49];
  assign P53[3] = IN1[3]&IN2[50];
  assign P54[2] = IN1[3]&IN2[51];
  assign P55[1] = IN1[3]&IN2[52];
  assign P56[0] = IN1[3]&IN2[53];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[4] = IN1[4]&IN2[12];
  assign P17[4] = IN1[4]&IN2[13];
  assign P18[4] = IN1[4]&IN2[14];
  assign P19[4] = IN1[4]&IN2[15];
  assign P20[4] = IN1[4]&IN2[16];
  assign P21[4] = IN1[4]&IN2[17];
  assign P22[4] = IN1[4]&IN2[18];
  assign P23[4] = IN1[4]&IN2[19];
  assign P24[4] = IN1[4]&IN2[20];
  assign P25[4] = IN1[4]&IN2[21];
  assign P26[4] = IN1[4]&IN2[22];
  assign P27[4] = IN1[4]&IN2[23];
  assign P28[4] = IN1[4]&IN2[24];
  assign P29[4] = IN1[4]&IN2[25];
  assign P30[4] = IN1[4]&IN2[26];
  assign P31[4] = IN1[4]&IN2[27];
  assign P32[4] = IN1[4]&IN2[28];
  assign P33[4] = IN1[4]&IN2[29];
  assign P34[4] = IN1[4]&IN2[30];
  assign P35[4] = IN1[4]&IN2[31];
  assign P36[4] = IN1[4]&IN2[32];
  assign P37[4] = IN1[4]&IN2[33];
  assign P38[4] = IN1[4]&IN2[34];
  assign P39[4] = IN1[4]&IN2[35];
  assign P40[4] = IN1[4]&IN2[36];
  assign P41[4] = IN1[4]&IN2[37];
  assign P42[4] = IN1[4]&IN2[38];
  assign P43[4] = IN1[4]&IN2[39];
  assign P44[4] = IN1[4]&IN2[40];
  assign P45[4] = IN1[4]&IN2[41];
  assign P46[4] = IN1[4]&IN2[42];
  assign P47[4] = IN1[4]&IN2[43];
  assign P48[4] = IN1[4]&IN2[44];
  assign P49[4] = IN1[4]&IN2[45];
  assign P50[4] = IN1[4]&IN2[46];
  assign P51[4] = IN1[4]&IN2[47];
  assign P52[4] = IN1[4]&IN2[48];
  assign P53[4] = IN1[4]&IN2[49];
  assign P54[3] = IN1[4]&IN2[50];
  assign P55[2] = IN1[4]&IN2[51];
  assign P56[1] = IN1[4]&IN2[52];
  assign P57[0] = IN1[4]&IN2[53];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[5] = IN1[5]&IN2[11];
  assign P17[5] = IN1[5]&IN2[12];
  assign P18[5] = IN1[5]&IN2[13];
  assign P19[5] = IN1[5]&IN2[14];
  assign P20[5] = IN1[5]&IN2[15];
  assign P21[5] = IN1[5]&IN2[16];
  assign P22[5] = IN1[5]&IN2[17];
  assign P23[5] = IN1[5]&IN2[18];
  assign P24[5] = IN1[5]&IN2[19];
  assign P25[5] = IN1[5]&IN2[20];
  assign P26[5] = IN1[5]&IN2[21];
  assign P27[5] = IN1[5]&IN2[22];
  assign P28[5] = IN1[5]&IN2[23];
  assign P29[5] = IN1[5]&IN2[24];
  assign P30[5] = IN1[5]&IN2[25];
  assign P31[5] = IN1[5]&IN2[26];
  assign P32[5] = IN1[5]&IN2[27];
  assign P33[5] = IN1[5]&IN2[28];
  assign P34[5] = IN1[5]&IN2[29];
  assign P35[5] = IN1[5]&IN2[30];
  assign P36[5] = IN1[5]&IN2[31];
  assign P37[5] = IN1[5]&IN2[32];
  assign P38[5] = IN1[5]&IN2[33];
  assign P39[5] = IN1[5]&IN2[34];
  assign P40[5] = IN1[5]&IN2[35];
  assign P41[5] = IN1[5]&IN2[36];
  assign P42[5] = IN1[5]&IN2[37];
  assign P43[5] = IN1[5]&IN2[38];
  assign P44[5] = IN1[5]&IN2[39];
  assign P45[5] = IN1[5]&IN2[40];
  assign P46[5] = IN1[5]&IN2[41];
  assign P47[5] = IN1[5]&IN2[42];
  assign P48[5] = IN1[5]&IN2[43];
  assign P49[5] = IN1[5]&IN2[44];
  assign P50[5] = IN1[5]&IN2[45];
  assign P51[5] = IN1[5]&IN2[46];
  assign P52[5] = IN1[5]&IN2[47];
  assign P53[5] = IN1[5]&IN2[48];
  assign P54[4] = IN1[5]&IN2[49];
  assign P55[3] = IN1[5]&IN2[50];
  assign P56[2] = IN1[5]&IN2[51];
  assign P57[1] = IN1[5]&IN2[52];
  assign P58[0] = IN1[5]&IN2[53];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[6] = IN1[6]&IN2[10];
  assign P17[6] = IN1[6]&IN2[11];
  assign P18[6] = IN1[6]&IN2[12];
  assign P19[6] = IN1[6]&IN2[13];
  assign P20[6] = IN1[6]&IN2[14];
  assign P21[6] = IN1[6]&IN2[15];
  assign P22[6] = IN1[6]&IN2[16];
  assign P23[6] = IN1[6]&IN2[17];
  assign P24[6] = IN1[6]&IN2[18];
  assign P25[6] = IN1[6]&IN2[19];
  assign P26[6] = IN1[6]&IN2[20];
  assign P27[6] = IN1[6]&IN2[21];
  assign P28[6] = IN1[6]&IN2[22];
  assign P29[6] = IN1[6]&IN2[23];
  assign P30[6] = IN1[6]&IN2[24];
  assign P31[6] = IN1[6]&IN2[25];
  assign P32[6] = IN1[6]&IN2[26];
  assign P33[6] = IN1[6]&IN2[27];
  assign P34[6] = IN1[6]&IN2[28];
  assign P35[6] = IN1[6]&IN2[29];
  assign P36[6] = IN1[6]&IN2[30];
  assign P37[6] = IN1[6]&IN2[31];
  assign P38[6] = IN1[6]&IN2[32];
  assign P39[6] = IN1[6]&IN2[33];
  assign P40[6] = IN1[6]&IN2[34];
  assign P41[6] = IN1[6]&IN2[35];
  assign P42[6] = IN1[6]&IN2[36];
  assign P43[6] = IN1[6]&IN2[37];
  assign P44[6] = IN1[6]&IN2[38];
  assign P45[6] = IN1[6]&IN2[39];
  assign P46[6] = IN1[6]&IN2[40];
  assign P47[6] = IN1[6]&IN2[41];
  assign P48[6] = IN1[6]&IN2[42];
  assign P49[6] = IN1[6]&IN2[43];
  assign P50[6] = IN1[6]&IN2[44];
  assign P51[6] = IN1[6]&IN2[45];
  assign P52[6] = IN1[6]&IN2[46];
  assign P53[6] = IN1[6]&IN2[47];
  assign P54[5] = IN1[6]&IN2[48];
  assign P55[4] = IN1[6]&IN2[49];
  assign P56[3] = IN1[6]&IN2[50];
  assign P57[2] = IN1[6]&IN2[51];
  assign P58[1] = IN1[6]&IN2[52];
  assign P59[0] = IN1[6]&IN2[53];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[7] = IN1[7]&IN2[9];
  assign P17[7] = IN1[7]&IN2[10];
  assign P18[7] = IN1[7]&IN2[11];
  assign P19[7] = IN1[7]&IN2[12];
  assign P20[7] = IN1[7]&IN2[13];
  assign P21[7] = IN1[7]&IN2[14];
  assign P22[7] = IN1[7]&IN2[15];
  assign P23[7] = IN1[7]&IN2[16];
  assign P24[7] = IN1[7]&IN2[17];
  assign P25[7] = IN1[7]&IN2[18];
  assign P26[7] = IN1[7]&IN2[19];
  assign P27[7] = IN1[7]&IN2[20];
  assign P28[7] = IN1[7]&IN2[21];
  assign P29[7] = IN1[7]&IN2[22];
  assign P30[7] = IN1[7]&IN2[23];
  assign P31[7] = IN1[7]&IN2[24];
  assign P32[7] = IN1[7]&IN2[25];
  assign P33[7] = IN1[7]&IN2[26];
  assign P34[7] = IN1[7]&IN2[27];
  assign P35[7] = IN1[7]&IN2[28];
  assign P36[7] = IN1[7]&IN2[29];
  assign P37[7] = IN1[7]&IN2[30];
  assign P38[7] = IN1[7]&IN2[31];
  assign P39[7] = IN1[7]&IN2[32];
  assign P40[7] = IN1[7]&IN2[33];
  assign P41[7] = IN1[7]&IN2[34];
  assign P42[7] = IN1[7]&IN2[35];
  assign P43[7] = IN1[7]&IN2[36];
  assign P44[7] = IN1[7]&IN2[37];
  assign P45[7] = IN1[7]&IN2[38];
  assign P46[7] = IN1[7]&IN2[39];
  assign P47[7] = IN1[7]&IN2[40];
  assign P48[7] = IN1[7]&IN2[41];
  assign P49[7] = IN1[7]&IN2[42];
  assign P50[7] = IN1[7]&IN2[43];
  assign P51[7] = IN1[7]&IN2[44];
  assign P52[7] = IN1[7]&IN2[45];
  assign P53[7] = IN1[7]&IN2[46];
  assign P54[6] = IN1[7]&IN2[47];
  assign P55[5] = IN1[7]&IN2[48];
  assign P56[4] = IN1[7]&IN2[49];
  assign P57[3] = IN1[7]&IN2[50];
  assign P58[2] = IN1[7]&IN2[51];
  assign P59[1] = IN1[7]&IN2[52];
  assign P60[0] = IN1[7]&IN2[53];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[8] = IN1[8]&IN2[8];
  assign P17[8] = IN1[8]&IN2[9];
  assign P18[8] = IN1[8]&IN2[10];
  assign P19[8] = IN1[8]&IN2[11];
  assign P20[8] = IN1[8]&IN2[12];
  assign P21[8] = IN1[8]&IN2[13];
  assign P22[8] = IN1[8]&IN2[14];
  assign P23[8] = IN1[8]&IN2[15];
  assign P24[8] = IN1[8]&IN2[16];
  assign P25[8] = IN1[8]&IN2[17];
  assign P26[8] = IN1[8]&IN2[18];
  assign P27[8] = IN1[8]&IN2[19];
  assign P28[8] = IN1[8]&IN2[20];
  assign P29[8] = IN1[8]&IN2[21];
  assign P30[8] = IN1[8]&IN2[22];
  assign P31[8] = IN1[8]&IN2[23];
  assign P32[8] = IN1[8]&IN2[24];
  assign P33[8] = IN1[8]&IN2[25];
  assign P34[8] = IN1[8]&IN2[26];
  assign P35[8] = IN1[8]&IN2[27];
  assign P36[8] = IN1[8]&IN2[28];
  assign P37[8] = IN1[8]&IN2[29];
  assign P38[8] = IN1[8]&IN2[30];
  assign P39[8] = IN1[8]&IN2[31];
  assign P40[8] = IN1[8]&IN2[32];
  assign P41[8] = IN1[8]&IN2[33];
  assign P42[8] = IN1[8]&IN2[34];
  assign P43[8] = IN1[8]&IN2[35];
  assign P44[8] = IN1[8]&IN2[36];
  assign P45[8] = IN1[8]&IN2[37];
  assign P46[8] = IN1[8]&IN2[38];
  assign P47[8] = IN1[8]&IN2[39];
  assign P48[8] = IN1[8]&IN2[40];
  assign P49[8] = IN1[8]&IN2[41];
  assign P50[8] = IN1[8]&IN2[42];
  assign P51[8] = IN1[8]&IN2[43];
  assign P52[8] = IN1[8]&IN2[44];
  assign P53[8] = IN1[8]&IN2[45];
  assign P54[7] = IN1[8]&IN2[46];
  assign P55[6] = IN1[8]&IN2[47];
  assign P56[5] = IN1[8]&IN2[48];
  assign P57[4] = IN1[8]&IN2[49];
  assign P58[3] = IN1[8]&IN2[50];
  assign P59[2] = IN1[8]&IN2[51];
  assign P60[1] = IN1[8]&IN2[52];
  assign P61[0] = IN1[8]&IN2[53];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[9] = IN1[9]&IN2[7];
  assign P17[9] = IN1[9]&IN2[8];
  assign P18[9] = IN1[9]&IN2[9];
  assign P19[9] = IN1[9]&IN2[10];
  assign P20[9] = IN1[9]&IN2[11];
  assign P21[9] = IN1[9]&IN2[12];
  assign P22[9] = IN1[9]&IN2[13];
  assign P23[9] = IN1[9]&IN2[14];
  assign P24[9] = IN1[9]&IN2[15];
  assign P25[9] = IN1[9]&IN2[16];
  assign P26[9] = IN1[9]&IN2[17];
  assign P27[9] = IN1[9]&IN2[18];
  assign P28[9] = IN1[9]&IN2[19];
  assign P29[9] = IN1[9]&IN2[20];
  assign P30[9] = IN1[9]&IN2[21];
  assign P31[9] = IN1[9]&IN2[22];
  assign P32[9] = IN1[9]&IN2[23];
  assign P33[9] = IN1[9]&IN2[24];
  assign P34[9] = IN1[9]&IN2[25];
  assign P35[9] = IN1[9]&IN2[26];
  assign P36[9] = IN1[9]&IN2[27];
  assign P37[9] = IN1[9]&IN2[28];
  assign P38[9] = IN1[9]&IN2[29];
  assign P39[9] = IN1[9]&IN2[30];
  assign P40[9] = IN1[9]&IN2[31];
  assign P41[9] = IN1[9]&IN2[32];
  assign P42[9] = IN1[9]&IN2[33];
  assign P43[9] = IN1[9]&IN2[34];
  assign P44[9] = IN1[9]&IN2[35];
  assign P45[9] = IN1[9]&IN2[36];
  assign P46[9] = IN1[9]&IN2[37];
  assign P47[9] = IN1[9]&IN2[38];
  assign P48[9] = IN1[9]&IN2[39];
  assign P49[9] = IN1[9]&IN2[40];
  assign P50[9] = IN1[9]&IN2[41];
  assign P51[9] = IN1[9]&IN2[42];
  assign P52[9] = IN1[9]&IN2[43];
  assign P53[9] = IN1[9]&IN2[44];
  assign P54[8] = IN1[9]&IN2[45];
  assign P55[7] = IN1[9]&IN2[46];
  assign P56[6] = IN1[9]&IN2[47];
  assign P57[5] = IN1[9]&IN2[48];
  assign P58[4] = IN1[9]&IN2[49];
  assign P59[3] = IN1[9]&IN2[50];
  assign P60[2] = IN1[9]&IN2[51];
  assign P61[1] = IN1[9]&IN2[52];
  assign P62[0] = IN1[9]&IN2[53];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[10] = IN1[10]&IN2[6];
  assign P17[10] = IN1[10]&IN2[7];
  assign P18[10] = IN1[10]&IN2[8];
  assign P19[10] = IN1[10]&IN2[9];
  assign P20[10] = IN1[10]&IN2[10];
  assign P21[10] = IN1[10]&IN2[11];
  assign P22[10] = IN1[10]&IN2[12];
  assign P23[10] = IN1[10]&IN2[13];
  assign P24[10] = IN1[10]&IN2[14];
  assign P25[10] = IN1[10]&IN2[15];
  assign P26[10] = IN1[10]&IN2[16];
  assign P27[10] = IN1[10]&IN2[17];
  assign P28[10] = IN1[10]&IN2[18];
  assign P29[10] = IN1[10]&IN2[19];
  assign P30[10] = IN1[10]&IN2[20];
  assign P31[10] = IN1[10]&IN2[21];
  assign P32[10] = IN1[10]&IN2[22];
  assign P33[10] = IN1[10]&IN2[23];
  assign P34[10] = IN1[10]&IN2[24];
  assign P35[10] = IN1[10]&IN2[25];
  assign P36[10] = IN1[10]&IN2[26];
  assign P37[10] = IN1[10]&IN2[27];
  assign P38[10] = IN1[10]&IN2[28];
  assign P39[10] = IN1[10]&IN2[29];
  assign P40[10] = IN1[10]&IN2[30];
  assign P41[10] = IN1[10]&IN2[31];
  assign P42[10] = IN1[10]&IN2[32];
  assign P43[10] = IN1[10]&IN2[33];
  assign P44[10] = IN1[10]&IN2[34];
  assign P45[10] = IN1[10]&IN2[35];
  assign P46[10] = IN1[10]&IN2[36];
  assign P47[10] = IN1[10]&IN2[37];
  assign P48[10] = IN1[10]&IN2[38];
  assign P49[10] = IN1[10]&IN2[39];
  assign P50[10] = IN1[10]&IN2[40];
  assign P51[10] = IN1[10]&IN2[41];
  assign P52[10] = IN1[10]&IN2[42];
  assign P53[10] = IN1[10]&IN2[43];
  assign P54[9] = IN1[10]&IN2[44];
  assign P55[8] = IN1[10]&IN2[45];
  assign P56[7] = IN1[10]&IN2[46];
  assign P57[6] = IN1[10]&IN2[47];
  assign P58[5] = IN1[10]&IN2[48];
  assign P59[4] = IN1[10]&IN2[49];
  assign P60[3] = IN1[10]&IN2[50];
  assign P61[2] = IN1[10]&IN2[51];
  assign P62[1] = IN1[10]&IN2[52];
  assign P63[0] = IN1[10]&IN2[53];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[11] = IN1[11]&IN2[5];
  assign P17[11] = IN1[11]&IN2[6];
  assign P18[11] = IN1[11]&IN2[7];
  assign P19[11] = IN1[11]&IN2[8];
  assign P20[11] = IN1[11]&IN2[9];
  assign P21[11] = IN1[11]&IN2[10];
  assign P22[11] = IN1[11]&IN2[11];
  assign P23[11] = IN1[11]&IN2[12];
  assign P24[11] = IN1[11]&IN2[13];
  assign P25[11] = IN1[11]&IN2[14];
  assign P26[11] = IN1[11]&IN2[15];
  assign P27[11] = IN1[11]&IN2[16];
  assign P28[11] = IN1[11]&IN2[17];
  assign P29[11] = IN1[11]&IN2[18];
  assign P30[11] = IN1[11]&IN2[19];
  assign P31[11] = IN1[11]&IN2[20];
  assign P32[11] = IN1[11]&IN2[21];
  assign P33[11] = IN1[11]&IN2[22];
  assign P34[11] = IN1[11]&IN2[23];
  assign P35[11] = IN1[11]&IN2[24];
  assign P36[11] = IN1[11]&IN2[25];
  assign P37[11] = IN1[11]&IN2[26];
  assign P38[11] = IN1[11]&IN2[27];
  assign P39[11] = IN1[11]&IN2[28];
  assign P40[11] = IN1[11]&IN2[29];
  assign P41[11] = IN1[11]&IN2[30];
  assign P42[11] = IN1[11]&IN2[31];
  assign P43[11] = IN1[11]&IN2[32];
  assign P44[11] = IN1[11]&IN2[33];
  assign P45[11] = IN1[11]&IN2[34];
  assign P46[11] = IN1[11]&IN2[35];
  assign P47[11] = IN1[11]&IN2[36];
  assign P48[11] = IN1[11]&IN2[37];
  assign P49[11] = IN1[11]&IN2[38];
  assign P50[11] = IN1[11]&IN2[39];
  assign P51[11] = IN1[11]&IN2[40];
  assign P52[11] = IN1[11]&IN2[41];
  assign P53[11] = IN1[11]&IN2[42];
  assign P54[10] = IN1[11]&IN2[43];
  assign P55[9] = IN1[11]&IN2[44];
  assign P56[8] = IN1[11]&IN2[45];
  assign P57[7] = IN1[11]&IN2[46];
  assign P58[6] = IN1[11]&IN2[47];
  assign P59[5] = IN1[11]&IN2[48];
  assign P60[4] = IN1[11]&IN2[49];
  assign P61[3] = IN1[11]&IN2[50];
  assign P62[2] = IN1[11]&IN2[51];
  assign P63[1] = IN1[11]&IN2[52];
  assign P64[0] = IN1[11]&IN2[53];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[12] = IN1[12]&IN2[4];
  assign P17[12] = IN1[12]&IN2[5];
  assign P18[12] = IN1[12]&IN2[6];
  assign P19[12] = IN1[12]&IN2[7];
  assign P20[12] = IN1[12]&IN2[8];
  assign P21[12] = IN1[12]&IN2[9];
  assign P22[12] = IN1[12]&IN2[10];
  assign P23[12] = IN1[12]&IN2[11];
  assign P24[12] = IN1[12]&IN2[12];
  assign P25[12] = IN1[12]&IN2[13];
  assign P26[12] = IN1[12]&IN2[14];
  assign P27[12] = IN1[12]&IN2[15];
  assign P28[12] = IN1[12]&IN2[16];
  assign P29[12] = IN1[12]&IN2[17];
  assign P30[12] = IN1[12]&IN2[18];
  assign P31[12] = IN1[12]&IN2[19];
  assign P32[12] = IN1[12]&IN2[20];
  assign P33[12] = IN1[12]&IN2[21];
  assign P34[12] = IN1[12]&IN2[22];
  assign P35[12] = IN1[12]&IN2[23];
  assign P36[12] = IN1[12]&IN2[24];
  assign P37[12] = IN1[12]&IN2[25];
  assign P38[12] = IN1[12]&IN2[26];
  assign P39[12] = IN1[12]&IN2[27];
  assign P40[12] = IN1[12]&IN2[28];
  assign P41[12] = IN1[12]&IN2[29];
  assign P42[12] = IN1[12]&IN2[30];
  assign P43[12] = IN1[12]&IN2[31];
  assign P44[12] = IN1[12]&IN2[32];
  assign P45[12] = IN1[12]&IN2[33];
  assign P46[12] = IN1[12]&IN2[34];
  assign P47[12] = IN1[12]&IN2[35];
  assign P48[12] = IN1[12]&IN2[36];
  assign P49[12] = IN1[12]&IN2[37];
  assign P50[12] = IN1[12]&IN2[38];
  assign P51[12] = IN1[12]&IN2[39];
  assign P52[12] = IN1[12]&IN2[40];
  assign P53[12] = IN1[12]&IN2[41];
  assign P54[11] = IN1[12]&IN2[42];
  assign P55[10] = IN1[12]&IN2[43];
  assign P56[9] = IN1[12]&IN2[44];
  assign P57[8] = IN1[12]&IN2[45];
  assign P58[7] = IN1[12]&IN2[46];
  assign P59[6] = IN1[12]&IN2[47];
  assign P60[5] = IN1[12]&IN2[48];
  assign P61[4] = IN1[12]&IN2[49];
  assign P62[3] = IN1[12]&IN2[50];
  assign P63[2] = IN1[12]&IN2[51];
  assign P64[1] = IN1[12]&IN2[52];
  assign P65[0] = IN1[12]&IN2[53];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[13] = IN1[13]&IN2[3];
  assign P17[13] = IN1[13]&IN2[4];
  assign P18[13] = IN1[13]&IN2[5];
  assign P19[13] = IN1[13]&IN2[6];
  assign P20[13] = IN1[13]&IN2[7];
  assign P21[13] = IN1[13]&IN2[8];
  assign P22[13] = IN1[13]&IN2[9];
  assign P23[13] = IN1[13]&IN2[10];
  assign P24[13] = IN1[13]&IN2[11];
  assign P25[13] = IN1[13]&IN2[12];
  assign P26[13] = IN1[13]&IN2[13];
  assign P27[13] = IN1[13]&IN2[14];
  assign P28[13] = IN1[13]&IN2[15];
  assign P29[13] = IN1[13]&IN2[16];
  assign P30[13] = IN1[13]&IN2[17];
  assign P31[13] = IN1[13]&IN2[18];
  assign P32[13] = IN1[13]&IN2[19];
  assign P33[13] = IN1[13]&IN2[20];
  assign P34[13] = IN1[13]&IN2[21];
  assign P35[13] = IN1[13]&IN2[22];
  assign P36[13] = IN1[13]&IN2[23];
  assign P37[13] = IN1[13]&IN2[24];
  assign P38[13] = IN1[13]&IN2[25];
  assign P39[13] = IN1[13]&IN2[26];
  assign P40[13] = IN1[13]&IN2[27];
  assign P41[13] = IN1[13]&IN2[28];
  assign P42[13] = IN1[13]&IN2[29];
  assign P43[13] = IN1[13]&IN2[30];
  assign P44[13] = IN1[13]&IN2[31];
  assign P45[13] = IN1[13]&IN2[32];
  assign P46[13] = IN1[13]&IN2[33];
  assign P47[13] = IN1[13]&IN2[34];
  assign P48[13] = IN1[13]&IN2[35];
  assign P49[13] = IN1[13]&IN2[36];
  assign P50[13] = IN1[13]&IN2[37];
  assign P51[13] = IN1[13]&IN2[38];
  assign P52[13] = IN1[13]&IN2[39];
  assign P53[13] = IN1[13]&IN2[40];
  assign P54[12] = IN1[13]&IN2[41];
  assign P55[11] = IN1[13]&IN2[42];
  assign P56[10] = IN1[13]&IN2[43];
  assign P57[9] = IN1[13]&IN2[44];
  assign P58[8] = IN1[13]&IN2[45];
  assign P59[7] = IN1[13]&IN2[46];
  assign P60[6] = IN1[13]&IN2[47];
  assign P61[5] = IN1[13]&IN2[48];
  assign P62[4] = IN1[13]&IN2[49];
  assign P63[3] = IN1[13]&IN2[50];
  assign P64[2] = IN1[13]&IN2[51];
  assign P65[1] = IN1[13]&IN2[52];
  assign P66[0] = IN1[13]&IN2[53];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[14] = IN1[14]&IN2[2];
  assign P17[14] = IN1[14]&IN2[3];
  assign P18[14] = IN1[14]&IN2[4];
  assign P19[14] = IN1[14]&IN2[5];
  assign P20[14] = IN1[14]&IN2[6];
  assign P21[14] = IN1[14]&IN2[7];
  assign P22[14] = IN1[14]&IN2[8];
  assign P23[14] = IN1[14]&IN2[9];
  assign P24[14] = IN1[14]&IN2[10];
  assign P25[14] = IN1[14]&IN2[11];
  assign P26[14] = IN1[14]&IN2[12];
  assign P27[14] = IN1[14]&IN2[13];
  assign P28[14] = IN1[14]&IN2[14];
  assign P29[14] = IN1[14]&IN2[15];
  assign P30[14] = IN1[14]&IN2[16];
  assign P31[14] = IN1[14]&IN2[17];
  assign P32[14] = IN1[14]&IN2[18];
  assign P33[14] = IN1[14]&IN2[19];
  assign P34[14] = IN1[14]&IN2[20];
  assign P35[14] = IN1[14]&IN2[21];
  assign P36[14] = IN1[14]&IN2[22];
  assign P37[14] = IN1[14]&IN2[23];
  assign P38[14] = IN1[14]&IN2[24];
  assign P39[14] = IN1[14]&IN2[25];
  assign P40[14] = IN1[14]&IN2[26];
  assign P41[14] = IN1[14]&IN2[27];
  assign P42[14] = IN1[14]&IN2[28];
  assign P43[14] = IN1[14]&IN2[29];
  assign P44[14] = IN1[14]&IN2[30];
  assign P45[14] = IN1[14]&IN2[31];
  assign P46[14] = IN1[14]&IN2[32];
  assign P47[14] = IN1[14]&IN2[33];
  assign P48[14] = IN1[14]&IN2[34];
  assign P49[14] = IN1[14]&IN2[35];
  assign P50[14] = IN1[14]&IN2[36];
  assign P51[14] = IN1[14]&IN2[37];
  assign P52[14] = IN1[14]&IN2[38];
  assign P53[14] = IN1[14]&IN2[39];
  assign P54[13] = IN1[14]&IN2[40];
  assign P55[12] = IN1[14]&IN2[41];
  assign P56[11] = IN1[14]&IN2[42];
  assign P57[10] = IN1[14]&IN2[43];
  assign P58[9] = IN1[14]&IN2[44];
  assign P59[8] = IN1[14]&IN2[45];
  assign P60[7] = IN1[14]&IN2[46];
  assign P61[6] = IN1[14]&IN2[47];
  assign P62[5] = IN1[14]&IN2[48];
  assign P63[4] = IN1[14]&IN2[49];
  assign P64[3] = IN1[14]&IN2[50];
  assign P65[2] = IN1[14]&IN2[51];
  assign P66[1] = IN1[14]&IN2[52];
  assign P67[0] = IN1[14]&IN2[53];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[15] = IN1[15]&IN2[1];
  assign P17[15] = IN1[15]&IN2[2];
  assign P18[15] = IN1[15]&IN2[3];
  assign P19[15] = IN1[15]&IN2[4];
  assign P20[15] = IN1[15]&IN2[5];
  assign P21[15] = IN1[15]&IN2[6];
  assign P22[15] = IN1[15]&IN2[7];
  assign P23[15] = IN1[15]&IN2[8];
  assign P24[15] = IN1[15]&IN2[9];
  assign P25[15] = IN1[15]&IN2[10];
  assign P26[15] = IN1[15]&IN2[11];
  assign P27[15] = IN1[15]&IN2[12];
  assign P28[15] = IN1[15]&IN2[13];
  assign P29[15] = IN1[15]&IN2[14];
  assign P30[15] = IN1[15]&IN2[15];
  assign P31[15] = IN1[15]&IN2[16];
  assign P32[15] = IN1[15]&IN2[17];
  assign P33[15] = IN1[15]&IN2[18];
  assign P34[15] = IN1[15]&IN2[19];
  assign P35[15] = IN1[15]&IN2[20];
  assign P36[15] = IN1[15]&IN2[21];
  assign P37[15] = IN1[15]&IN2[22];
  assign P38[15] = IN1[15]&IN2[23];
  assign P39[15] = IN1[15]&IN2[24];
  assign P40[15] = IN1[15]&IN2[25];
  assign P41[15] = IN1[15]&IN2[26];
  assign P42[15] = IN1[15]&IN2[27];
  assign P43[15] = IN1[15]&IN2[28];
  assign P44[15] = IN1[15]&IN2[29];
  assign P45[15] = IN1[15]&IN2[30];
  assign P46[15] = IN1[15]&IN2[31];
  assign P47[15] = IN1[15]&IN2[32];
  assign P48[15] = IN1[15]&IN2[33];
  assign P49[15] = IN1[15]&IN2[34];
  assign P50[15] = IN1[15]&IN2[35];
  assign P51[15] = IN1[15]&IN2[36];
  assign P52[15] = IN1[15]&IN2[37];
  assign P53[15] = IN1[15]&IN2[38];
  assign P54[14] = IN1[15]&IN2[39];
  assign P55[13] = IN1[15]&IN2[40];
  assign P56[12] = IN1[15]&IN2[41];
  assign P57[11] = IN1[15]&IN2[42];
  assign P58[10] = IN1[15]&IN2[43];
  assign P59[9] = IN1[15]&IN2[44];
  assign P60[8] = IN1[15]&IN2[45];
  assign P61[7] = IN1[15]&IN2[46];
  assign P62[6] = IN1[15]&IN2[47];
  assign P63[5] = IN1[15]&IN2[48];
  assign P64[4] = IN1[15]&IN2[49];
  assign P65[3] = IN1[15]&IN2[50];
  assign P66[2] = IN1[15]&IN2[51];
  assign P67[1] = IN1[15]&IN2[52];
  assign P68[0] = IN1[15]&IN2[53];
  assign P16[16] = IN1[16]&IN2[0];
  assign P17[16] = IN1[16]&IN2[1];
  assign P18[16] = IN1[16]&IN2[2];
  assign P19[16] = IN1[16]&IN2[3];
  assign P20[16] = IN1[16]&IN2[4];
  assign P21[16] = IN1[16]&IN2[5];
  assign P22[16] = IN1[16]&IN2[6];
  assign P23[16] = IN1[16]&IN2[7];
  assign P24[16] = IN1[16]&IN2[8];
  assign P25[16] = IN1[16]&IN2[9];
  assign P26[16] = IN1[16]&IN2[10];
  assign P27[16] = IN1[16]&IN2[11];
  assign P28[16] = IN1[16]&IN2[12];
  assign P29[16] = IN1[16]&IN2[13];
  assign P30[16] = IN1[16]&IN2[14];
  assign P31[16] = IN1[16]&IN2[15];
  assign P32[16] = IN1[16]&IN2[16];
  assign P33[16] = IN1[16]&IN2[17];
  assign P34[16] = IN1[16]&IN2[18];
  assign P35[16] = IN1[16]&IN2[19];
  assign P36[16] = IN1[16]&IN2[20];
  assign P37[16] = IN1[16]&IN2[21];
  assign P38[16] = IN1[16]&IN2[22];
  assign P39[16] = IN1[16]&IN2[23];
  assign P40[16] = IN1[16]&IN2[24];
  assign P41[16] = IN1[16]&IN2[25];
  assign P42[16] = IN1[16]&IN2[26];
  assign P43[16] = IN1[16]&IN2[27];
  assign P44[16] = IN1[16]&IN2[28];
  assign P45[16] = IN1[16]&IN2[29];
  assign P46[16] = IN1[16]&IN2[30];
  assign P47[16] = IN1[16]&IN2[31];
  assign P48[16] = IN1[16]&IN2[32];
  assign P49[16] = IN1[16]&IN2[33];
  assign P50[16] = IN1[16]&IN2[34];
  assign P51[16] = IN1[16]&IN2[35];
  assign P52[16] = IN1[16]&IN2[36];
  assign P53[16] = IN1[16]&IN2[37];
  assign P54[15] = IN1[16]&IN2[38];
  assign P55[14] = IN1[16]&IN2[39];
  assign P56[13] = IN1[16]&IN2[40];
  assign P57[12] = IN1[16]&IN2[41];
  assign P58[11] = IN1[16]&IN2[42];
  assign P59[10] = IN1[16]&IN2[43];
  assign P60[9] = IN1[16]&IN2[44];
  assign P61[8] = IN1[16]&IN2[45];
  assign P62[7] = IN1[16]&IN2[46];
  assign P63[6] = IN1[16]&IN2[47];
  assign P64[5] = IN1[16]&IN2[48];
  assign P65[4] = IN1[16]&IN2[49];
  assign P66[3] = IN1[16]&IN2[50];
  assign P67[2] = IN1[16]&IN2[51];
  assign P68[1] = IN1[16]&IN2[52];
  assign P69[0] = IN1[16]&IN2[53];
  assign P17[17] = IN1[17]&IN2[0];
  assign P18[17] = IN1[17]&IN2[1];
  assign P19[17] = IN1[17]&IN2[2];
  assign P20[17] = IN1[17]&IN2[3];
  assign P21[17] = IN1[17]&IN2[4];
  assign P22[17] = IN1[17]&IN2[5];
  assign P23[17] = IN1[17]&IN2[6];
  assign P24[17] = IN1[17]&IN2[7];
  assign P25[17] = IN1[17]&IN2[8];
  assign P26[17] = IN1[17]&IN2[9];
  assign P27[17] = IN1[17]&IN2[10];
  assign P28[17] = IN1[17]&IN2[11];
  assign P29[17] = IN1[17]&IN2[12];
  assign P30[17] = IN1[17]&IN2[13];
  assign P31[17] = IN1[17]&IN2[14];
  assign P32[17] = IN1[17]&IN2[15];
  assign P33[17] = IN1[17]&IN2[16];
  assign P34[17] = IN1[17]&IN2[17];
  assign P35[17] = IN1[17]&IN2[18];
  assign P36[17] = IN1[17]&IN2[19];
  assign P37[17] = IN1[17]&IN2[20];
  assign P38[17] = IN1[17]&IN2[21];
  assign P39[17] = IN1[17]&IN2[22];
  assign P40[17] = IN1[17]&IN2[23];
  assign P41[17] = IN1[17]&IN2[24];
  assign P42[17] = IN1[17]&IN2[25];
  assign P43[17] = IN1[17]&IN2[26];
  assign P44[17] = IN1[17]&IN2[27];
  assign P45[17] = IN1[17]&IN2[28];
  assign P46[17] = IN1[17]&IN2[29];
  assign P47[17] = IN1[17]&IN2[30];
  assign P48[17] = IN1[17]&IN2[31];
  assign P49[17] = IN1[17]&IN2[32];
  assign P50[17] = IN1[17]&IN2[33];
  assign P51[17] = IN1[17]&IN2[34];
  assign P52[17] = IN1[17]&IN2[35];
  assign P53[17] = IN1[17]&IN2[36];
  assign P54[16] = IN1[17]&IN2[37];
  assign P55[15] = IN1[17]&IN2[38];
  assign P56[14] = IN1[17]&IN2[39];
  assign P57[13] = IN1[17]&IN2[40];
  assign P58[12] = IN1[17]&IN2[41];
  assign P59[11] = IN1[17]&IN2[42];
  assign P60[10] = IN1[17]&IN2[43];
  assign P61[9] = IN1[17]&IN2[44];
  assign P62[8] = IN1[17]&IN2[45];
  assign P63[7] = IN1[17]&IN2[46];
  assign P64[6] = IN1[17]&IN2[47];
  assign P65[5] = IN1[17]&IN2[48];
  assign P66[4] = IN1[17]&IN2[49];
  assign P67[3] = IN1[17]&IN2[50];
  assign P68[2] = IN1[17]&IN2[51];
  assign P69[1] = IN1[17]&IN2[52];
  assign P70[0] = IN1[17]&IN2[53];
  assign P18[18] = IN1[18]&IN2[0];
  assign P19[18] = IN1[18]&IN2[1];
  assign P20[18] = IN1[18]&IN2[2];
  assign P21[18] = IN1[18]&IN2[3];
  assign P22[18] = IN1[18]&IN2[4];
  assign P23[18] = IN1[18]&IN2[5];
  assign P24[18] = IN1[18]&IN2[6];
  assign P25[18] = IN1[18]&IN2[7];
  assign P26[18] = IN1[18]&IN2[8];
  assign P27[18] = IN1[18]&IN2[9];
  assign P28[18] = IN1[18]&IN2[10];
  assign P29[18] = IN1[18]&IN2[11];
  assign P30[18] = IN1[18]&IN2[12];
  assign P31[18] = IN1[18]&IN2[13];
  assign P32[18] = IN1[18]&IN2[14];
  assign P33[18] = IN1[18]&IN2[15];
  assign P34[18] = IN1[18]&IN2[16];
  assign P35[18] = IN1[18]&IN2[17];
  assign P36[18] = IN1[18]&IN2[18];
  assign P37[18] = IN1[18]&IN2[19];
  assign P38[18] = IN1[18]&IN2[20];
  assign P39[18] = IN1[18]&IN2[21];
  assign P40[18] = IN1[18]&IN2[22];
  assign P41[18] = IN1[18]&IN2[23];
  assign P42[18] = IN1[18]&IN2[24];
  assign P43[18] = IN1[18]&IN2[25];
  assign P44[18] = IN1[18]&IN2[26];
  assign P45[18] = IN1[18]&IN2[27];
  assign P46[18] = IN1[18]&IN2[28];
  assign P47[18] = IN1[18]&IN2[29];
  assign P48[18] = IN1[18]&IN2[30];
  assign P49[18] = IN1[18]&IN2[31];
  assign P50[18] = IN1[18]&IN2[32];
  assign P51[18] = IN1[18]&IN2[33];
  assign P52[18] = IN1[18]&IN2[34];
  assign P53[18] = IN1[18]&IN2[35];
  assign P54[17] = IN1[18]&IN2[36];
  assign P55[16] = IN1[18]&IN2[37];
  assign P56[15] = IN1[18]&IN2[38];
  assign P57[14] = IN1[18]&IN2[39];
  assign P58[13] = IN1[18]&IN2[40];
  assign P59[12] = IN1[18]&IN2[41];
  assign P60[11] = IN1[18]&IN2[42];
  assign P61[10] = IN1[18]&IN2[43];
  assign P62[9] = IN1[18]&IN2[44];
  assign P63[8] = IN1[18]&IN2[45];
  assign P64[7] = IN1[18]&IN2[46];
  assign P65[6] = IN1[18]&IN2[47];
  assign P66[5] = IN1[18]&IN2[48];
  assign P67[4] = IN1[18]&IN2[49];
  assign P68[3] = IN1[18]&IN2[50];
  assign P69[2] = IN1[18]&IN2[51];
  assign P70[1] = IN1[18]&IN2[52];
  assign P71[0] = IN1[18]&IN2[53];
  assign P19[19] = IN1[19]&IN2[0];
  assign P20[19] = IN1[19]&IN2[1];
  assign P21[19] = IN1[19]&IN2[2];
  assign P22[19] = IN1[19]&IN2[3];
  assign P23[19] = IN1[19]&IN2[4];
  assign P24[19] = IN1[19]&IN2[5];
  assign P25[19] = IN1[19]&IN2[6];
  assign P26[19] = IN1[19]&IN2[7];
  assign P27[19] = IN1[19]&IN2[8];
  assign P28[19] = IN1[19]&IN2[9];
  assign P29[19] = IN1[19]&IN2[10];
  assign P30[19] = IN1[19]&IN2[11];
  assign P31[19] = IN1[19]&IN2[12];
  assign P32[19] = IN1[19]&IN2[13];
  assign P33[19] = IN1[19]&IN2[14];
  assign P34[19] = IN1[19]&IN2[15];
  assign P35[19] = IN1[19]&IN2[16];
  assign P36[19] = IN1[19]&IN2[17];
  assign P37[19] = IN1[19]&IN2[18];
  assign P38[19] = IN1[19]&IN2[19];
  assign P39[19] = IN1[19]&IN2[20];
  assign P40[19] = IN1[19]&IN2[21];
  assign P41[19] = IN1[19]&IN2[22];
  assign P42[19] = IN1[19]&IN2[23];
  assign P43[19] = IN1[19]&IN2[24];
  assign P44[19] = IN1[19]&IN2[25];
  assign P45[19] = IN1[19]&IN2[26];
  assign P46[19] = IN1[19]&IN2[27];
  assign P47[19] = IN1[19]&IN2[28];
  assign P48[19] = IN1[19]&IN2[29];
  assign P49[19] = IN1[19]&IN2[30];
  assign P50[19] = IN1[19]&IN2[31];
  assign P51[19] = IN1[19]&IN2[32];
  assign P52[19] = IN1[19]&IN2[33];
  assign P53[19] = IN1[19]&IN2[34];
  assign P54[18] = IN1[19]&IN2[35];
  assign P55[17] = IN1[19]&IN2[36];
  assign P56[16] = IN1[19]&IN2[37];
  assign P57[15] = IN1[19]&IN2[38];
  assign P58[14] = IN1[19]&IN2[39];
  assign P59[13] = IN1[19]&IN2[40];
  assign P60[12] = IN1[19]&IN2[41];
  assign P61[11] = IN1[19]&IN2[42];
  assign P62[10] = IN1[19]&IN2[43];
  assign P63[9] = IN1[19]&IN2[44];
  assign P64[8] = IN1[19]&IN2[45];
  assign P65[7] = IN1[19]&IN2[46];
  assign P66[6] = IN1[19]&IN2[47];
  assign P67[5] = IN1[19]&IN2[48];
  assign P68[4] = IN1[19]&IN2[49];
  assign P69[3] = IN1[19]&IN2[50];
  assign P70[2] = IN1[19]&IN2[51];
  assign P71[1] = IN1[19]&IN2[52];
  assign P72[0] = IN1[19]&IN2[53];
  assign P20[20] = IN1[20]&IN2[0];
  assign P21[20] = IN1[20]&IN2[1];
  assign P22[20] = IN1[20]&IN2[2];
  assign P23[20] = IN1[20]&IN2[3];
  assign P24[20] = IN1[20]&IN2[4];
  assign P25[20] = IN1[20]&IN2[5];
  assign P26[20] = IN1[20]&IN2[6];
  assign P27[20] = IN1[20]&IN2[7];
  assign P28[20] = IN1[20]&IN2[8];
  assign P29[20] = IN1[20]&IN2[9];
  assign P30[20] = IN1[20]&IN2[10];
  assign P31[20] = IN1[20]&IN2[11];
  assign P32[20] = IN1[20]&IN2[12];
  assign P33[20] = IN1[20]&IN2[13];
  assign P34[20] = IN1[20]&IN2[14];
  assign P35[20] = IN1[20]&IN2[15];
  assign P36[20] = IN1[20]&IN2[16];
  assign P37[20] = IN1[20]&IN2[17];
  assign P38[20] = IN1[20]&IN2[18];
  assign P39[20] = IN1[20]&IN2[19];
  assign P40[20] = IN1[20]&IN2[20];
  assign P41[20] = IN1[20]&IN2[21];
  assign P42[20] = IN1[20]&IN2[22];
  assign P43[20] = IN1[20]&IN2[23];
  assign P44[20] = IN1[20]&IN2[24];
  assign P45[20] = IN1[20]&IN2[25];
  assign P46[20] = IN1[20]&IN2[26];
  assign P47[20] = IN1[20]&IN2[27];
  assign P48[20] = IN1[20]&IN2[28];
  assign P49[20] = IN1[20]&IN2[29];
  assign P50[20] = IN1[20]&IN2[30];
  assign P51[20] = IN1[20]&IN2[31];
  assign P52[20] = IN1[20]&IN2[32];
  assign P53[20] = IN1[20]&IN2[33];
  assign P54[19] = IN1[20]&IN2[34];
  assign P55[18] = IN1[20]&IN2[35];
  assign P56[17] = IN1[20]&IN2[36];
  assign P57[16] = IN1[20]&IN2[37];
  assign P58[15] = IN1[20]&IN2[38];
  assign P59[14] = IN1[20]&IN2[39];
  assign P60[13] = IN1[20]&IN2[40];
  assign P61[12] = IN1[20]&IN2[41];
  assign P62[11] = IN1[20]&IN2[42];
  assign P63[10] = IN1[20]&IN2[43];
  assign P64[9] = IN1[20]&IN2[44];
  assign P65[8] = IN1[20]&IN2[45];
  assign P66[7] = IN1[20]&IN2[46];
  assign P67[6] = IN1[20]&IN2[47];
  assign P68[5] = IN1[20]&IN2[48];
  assign P69[4] = IN1[20]&IN2[49];
  assign P70[3] = IN1[20]&IN2[50];
  assign P71[2] = IN1[20]&IN2[51];
  assign P72[1] = IN1[20]&IN2[52];
  assign P73[0] = IN1[20]&IN2[53];
  assign P21[21] = IN1[21]&IN2[0];
  assign P22[21] = IN1[21]&IN2[1];
  assign P23[21] = IN1[21]&IN2[2];
  assign P24[21] = IN1[21]&IN2[3];
  assign P25[21] = IN1[21]&IN2[4];
  assign P26[21] = IN1[21]&IN2[5];
  assign P27[21] = IN1[21]&IN2[6];
  assign P28[21] = IN1[21]&IN2[7];
  assign P29[21] = IN1[21]&IN2[8];
  assign P30[21] = IN1[21]&IN2[9];
  assign P31[21] = IN1[21]&IN2[10];
  assign P32[21] = IN1[21]&IN2[11];
  assign P33[21] = IN1[21]&IN2[12];
  assign P34[21] = IN1[21]&IN2[13];
  assign P35[21] = IN1[21]&IN2[14];
  assign P36[21] = IN1[21]&IN2[15];
  assign P37[21] = IN1[21]&IN2[16];
  assign P38[21] = IN1[21]&IN2[17];
  assign P39[21] = IN1[21]&IN2[18];
  assign P40[21] = IN1[21]&IN2[19];
  assign P41[21] = IN1[21]&IN2[20];
  assign P42[21] = IN1[21]&IN2[21];
  assign P43[21] = IN1[21]&IN2[22];
  assign P44[21] = IN1[21]&IN2[23];
  assign P45[21] = IN1[21]&IN2[24];
  assign P46[21] = IN1[21]&IN2[25];
  assign P47[21] = IN1[21]&IN2[26];
  assign P48[21] = IN1[21]&IN2[27];
  assign P49[21] = IN1[21]&IN2[28];
  assign P50[21] = IN1[21]&IN2[29];
  assign P51[21] = IN1[21]&IN2[30];
  assign P52[21] = IN1[21]&IN2[31];
  assign P53[21] = IN1[21]&IN2[32];
  assign P54[20] = IN1[21]&IN2[33];
  assign P55[19] = IN1[21]&IN2[34];
  assign P56[18] = IN1[21]&IN2[35];
  assign P57[17] = IN1[21]&IN2[36];
  assign P58[16] = IN1[21]&IN2[37];
  assign P59[15] = IN1[21]&IN2[38];
  assign P60[14] = IN1[21]&IN2[39];
  assign P61[13] = IN1[21]&IN2[40];
  assign P62[12] = IN1[21]&IN2[41];
  assign P63[11] = IN1[21]&IN2[42];
  assign P64[10] = IN1[21]&IN2[43];
  assign P65[9] = IN1[21]&IN2[44];
  assign P66[8] = IN1[21]&IN2[45];
  assign P67[7] = IN1[21]&IN2[46];
  assign P68[6] = IN1[21]&IN2[47];
  assign P69[5] = IN1[21]&IN2[48];
  assign P70[4] = IN1[21]&IN2[49];
  assign P71[3] = IN1[21]&IN2[50];
  assign P72[2] = IN1[21]&IN2[51];
  assign P73[1] = IN1[21]&IN2[52];
  assign P74[0] = IN1[21]&IN2[53];
  assign P22[22] = IN1[22]&IN2[0];
  assign P23[22] = IN1[22]&IN2[1];
  assign P24[22] = IN1[22]&IN2[2];
  assign P25[22] = IN1[22]&IN2[3];
  assign P26[22] = IN1[22]&IN2[4];
  assign P27[22] = IN1[22]&IN2[5];
  assign P28[22] = IN1[22]&IN2[6];
  assign P29[22] = IN1[22]&IN2[7];
  assign P30[22] = IN1[22]&IN2[8];
  assign P31[22] = IN1[22]&IN2[9];
  assign P32[22] = IN1[22]&IN2[10];
  assign P33[22] = IN1[22]&IN2[11];
  assign P34[22] = IN1[22]&IN2[12];
  assign P35[22] = IN1[22]&IN2[13];
  assign P36[22] = IN1[22]&IN2[14];
  assign P37[22] = IN1[22]&IN2[15];
  assign P38[22] = IN1[22]&IN2[16];
  assign P39[22] = IN1[22]&IN2[17];
  assign P40[22] = IN1[22]&IN2[18];
  assign P41[22] = IN1[22]&IN2[19];
  assign P42[22] = IN1[22]&IN2[20];
  assign P43[22] = IN1[22]&IN2[21];
  assign P44[22] = IN1[22]&IN2[22];
  assign P45[22] = IN1[22]&IN2[23];
  assign P46[22] = IN1[22]&IN2[24];
  assign P47[22] = IN1[22]&IN2[25];
  assign P48[22] = IN1[22]&IN2[26];
  assign P49[22] = IN1[22]&IN2[27];
  assign P50[22] = IN1[22]&IN2[28];
  assign P51[22] = IN1[22]&IN2[29];
  assign P52[22] = IN1[22]&IN2[30];
  assign P53[22] = IN1[22]&IN2[31];
  assign P54[21] = IN1[22]&IN2[32];
  assign P55[20] = IN1[22]&IN2[33];
  assign P56[19] = IN1[22]&IN2[34];
  assign P57[18] = IN1[22]&IN2[35];
  assign P58[17] = IN1[22]&IN2[36];
  assign P59[16] = IN1[22]&IN2[37];
  assign P60[15] = IN1[22]&IN2[38];
  assign P61[14] = IN1[22]&IN2[39];
  assign P62[13] = IN1[22]&IN2[40];
  assign P63[12] = IN1[22]&IN2[41];
  assign P64[11] = IN1[22]&IN2[42];
  assign P65[10] = IN1[22]&IN2[43];
  assign P66[9] = IN1[22]&IN2[44];
  assign P67[8] = IN1[22]&IN2[45];
  assign P68[7] = IN1[22]&IN2[46];
  assign P69[6] = IN1[22]&IN2[47];
  assign P70[5] = IN1[22]&IN2[48];
  assign P71[4] = IN1[22]&IN2[49];
  assign P72[3] = IN1[22]&IN2[50];
  assign P73[2] = IN1[22]&IN2[51];
  assign P74[1] = IN1[22]&IN2[52];
  assign P75[0] = IN1[22]&IN2[53];
  assign P23[23] = IN1[23]&IN2[0];
  assign P24[23] = IN1[23]&IN2[1];
  assign P25[23] = IN1[23]&IN2[2];
  assign P26[23] = IN1[23]&IN2[3];
  assign P27[23] = IN1[23]&IN2[4];
  assign P28[23] = IN1[23]&IN2[5];
  assign P29[23] = IN1[23]&IN2[6];
  assign P30[23] = IN1[23]&IN2[7];
  assign P31[23] = IN1[23]&IN2[8];
  assign P32[23] = IN1[23]&IN2[9];
  assign P33[23] = IN1[23]&IN2[10];
  assign P34[23] = IN1[23]&IN2[11];
  assign P35[23] = IN1[23]&IN2[12];
  assign P36[23] = IN1[23]&IN2[13];
  assign P37[23] = IN1[23]&IN2[14];
  assign P38[23] = IN1[23]&IN2[15];
  assign P39[23] = IN1[23]&IN2[16];
  assign P40[23] = IN1[23]&IN2[17];
  assign P41[23] = IN1[23]&IN2[18];
  assign P42[23] = IN1[23]&IN2[19];
  assign P43[23] = IN1[23]&IN2[20];
  assign P44[23] = IN1[23]&IN2[21];
  assign P45[23] = IN1[23]&IN2[22];
  assign P46[23] = IN1[23]&IN2[23];
  assign P47[23] = IN1[23]&IN2[24];
  assign P48[23] = IN1[23]&IN2[25];
  assign P49[23] = IN1[23]&IN2[26];
  assign P50[23] = IN1[23]&IN2[27];
  assign P51[23] = IN1[23]&IN2[28];
  assign P52[23] = IN1[23]&IN2[29];
  assign P53[23] = IN1[23]&IN2[30];
  assign P54[22] = IN1[23]&IN2[31];
  assign P55[21] = IN1[23]&IN2[32];
  assign P56[20] = IN1[23]&IN2[33];
  assign P57[19] = IN1[23]&IN2[34];
  assign P58[18] = IN1[23]&IN2[35];
  assign P59[17] = IN1[23]&IN2[36];
  assign P60[16] = IN1[23]&IN2[37];
  assign P61[15] = IN1[23]&IN2[38];
  assign P62[14] = IN1[23]&IN2[39];
  assign P63[13] = IN1[23]&IN2[40];
  assign P64[12] = IN1[23]&IN2[41];
  assign P65[11] = IN1[23]&IN2[42];
  assign P66[10] = IN1[23]&IN2[43];
  assign P67[9] = IN1[23]&IN2[44];
  assign P68[8] = IN1[23]&IN2[45];
  assign P69[7] = IN1[23]&IN2[46];
  assign P70[6] = IN1[23]&IN2[47];
  assign P71[5] = IN1[23]&IN2[48];
  assign P72[4] = IN1[23]&IN2[49];
  assign P73[3] = IN1[23]&IN2[50];
  assign P74[2] = IN1[23]&IN2[51];
  assign P75[1] = IN1[23]&IN2[52];
  assign P76[0] = IN1[23]&IN2[53];
  assign P24[24] = IN1[24]&IN2[0];
  assign P25[24] = IN1[24]&IN2[1];
  assign P26[24] = IN1[24]&IN2[2];
  assign P27[24] = IN1[24]&IN2[3];
  assign P28[24] = IN1[24]&IN2[4];
  assign P29[24] = IN1[24]&IN2[5];
  assign P30[24] = IN1[24]&IN2[6];
  assign P31[24] = IN1[24]&IN2[7];
  assign P32[24] = IN1[24]&IN2[8];
  assign P33[24] = IN1[24]&IN2[9];
  assign P34[24] = IN1[24]&IN2[10];
  assign P35[24] = IN1[24]&IN2[11];
  assign P36[24] = IN1[24]&IN2[12];
  assign P37[24] = IN1[24]&IN2[13];
  assign P38[24] = IN1[24]&IN2[14];
  assign P39[24] = IN1[24]&IN2[15];
  assign P40[24] = IN1[24]&IN2[16];
  assign P41[24] = IN1[24]&IN2[17];
  assign P42[24] = IN1[24]&IN2[18];
  assign P43[24] = IN1[24]&IN2[19];
  assign P44[24] = IN1[24]&IN2[20];
  assign P45[24] = IN1[24]&IN2[21];
  assign P46[24] = IN1[24]&IN2[22];
  assign P47[24] = IN1[24]&IN2[23];
  assign P48[24] = IN1[24]&IN2[24];
  assign P49[24] = IN1[24]&IN2[25];
  assign P50[24] = IN1[24]&IN2[26];
  assign P51[24] = IN1[24]&IN2[27];
  assign P52[24] = IN1[24]&IN2[28];
  assign P53[24] = IN1[24]&IN2[29];
  assign P54[23] = IN1[24]&IN2[30];
  assign P55[22] = IN1[24]&IN2[31];
  assign P56[21] = IN1[24]&IN2[32];
  assign P57[20] = IN1[24]&IN2[33];
  assign P58[19] = IN1[24]&IN2[34];
  assign P59[18] = IN1[24]&IN2[35];
  assign P60[17] = IN1[24]&IN2[36];
  assign P61[16] = IN1[24]&IN2[37];
  assign P62[15] = IN1[24]&IN2[38];
  assign P63[14] = IN1[24]&IN2[39];
  assign P64[13] = IN1[24]&IN2[40];
  assign P65[12] = IN1[24]&IN2[41];
  assign P66[11] = IN1[24]&IN2[42];
  assign P67[10] = IN1[24]&IN2[43];
  assign P68[9] = IN1[24]&IN2[44];
  assign P69[8] = IN1[24]&IN2[45];
  assign P70[7] = IN1[24]&IN2[46];
  assign P71[6] = IN1[24]&IN2[47];
  assign P72[5] = IN1[24]&IN2[48];
  assign P73[4] = IN1[24]&IN2[49];
  assign P74[3] = IN1[24]&IN2[50];
  assign P75[2] = IN1[24]&IN2[51];
  assign P76[1] = IN1[24]&IN2[52];
  assign P77[0] = IN1[24]&IN2[53];
  assign P25[25] = IN1[25]&IN2[0];
  assign P26[25] = IN1[25]&IN2[1];
  assign P27[25] = IN1[25]&IN2[2];
  assign P28[25] = IN1[25]&IN2[3];
  assign P29[25] = IN1[25]&IN2[4];
  assign P30[25] = IN1[25]&IN2[5];
  assign P31[25] = IN1[25]&IN2[6];
  assign P32[25] = IN1[25]&IN2[7];
  assign P33[25] = IN1[25]&IN2[8];
  assign P34[25] = IN1[25]&IN2[9];
  assign P35[25] = IN1[25]&IN2[10];
  assign P36[25] = IN1[25]&IN2[11];
  assign P37[25] = IN1[25]&IN2[12];
  assign P38[25] = IN1[25]&IN2[13];
  assign P39[25] = IN1[25]&IN2[14];
  assign P40[25] = IN1[25]&IN2[15];
  assign P41[25] = IN1[25]&IN2[16];
  assign P42[25] = IN1[25]&IN2[17];
  assign P43[25] = IN1[25]&IN2[18];
  assign P44[25] = IN1[25]&IN2[19];
  assign P45[25] = IN1[25]&IN2[20];
  assign P46[25] = IN1[25]&IN2[21];
  assign P47[25] = IN1[25]&IN2[22];
  assign P48[25] = IN1[25]&IN2[23];
  assign P49[25] = IN1[25]&IN2[24];
  assign P50[25] = IN1[25]&IN2[25];
  assign P51[25] = IN1[25]&IN2[26];
  assign P52[25] = IN1[25]&IN2[27];
  assign P53[25] = IN1[25]&IN2[28];
  assign P54[24] = IN1[25]&IN2[29];
  assign P55[23] = IN1[25]&IN2[30];
  assign P56[22] = IN1[25]&IN2[31];
  assign P57[21] = IN1[25]&IN2[32];
  assign P58[20] = IN1[25]&IN2[33];
  assign P59[19] = IN1[25]&IN2[34];
  assign P60[18] = IN1[25]&IN2[35];
  assign P61[17] = IN1[25]&IN2[36];
  assign P62[16] = IN1[25]&IN2[37];
  assign P63[15] = IN1[25]&IN2[38];
  assign P64[14] = IN1[25]&IN2[39];
  assign P65[13] = IN1[25]&IN2[40];
  assign P66[12] = IN1[25]&IN2[41];
  assign P67[11] = IN1[25]&IN2[42];
  assign P68[10] = IN1[25]&IN2[43];
  assign P69[9] = IN1[25]&IN2[44];
  assign P70[8] = IN1[25]&IN2[45];
  assign P71[7] = IN1[25]&IN2[46];
  assign P72[6] = IN1[25]&IN2[47];
  assign P73[5] = IN1[25]&IN2[48];
  assign P74[4] = IN1[25]&IN2[49];
  assign P75[3] = IN1[25]&IN2[50];
  assign P76[2] = IN1[25]&IN2[51];
  assign P77[1] = IN1[25]&IN2[52];
  assign P78[0] = IN1[25]&IN2[53];
  assign P26[26] = IN1[26]&IN2[0];
  assign P27[26] = IN1[26]&IN2[1];
  assign P28[26] = IN1[26]&IN2[2];
  assign P29[26] = IN1[26]&IN2[3];
  assign P30[26] = IN1[26]&IN2[4];
  assign P31[26] = IN1[26]&IN2[5];
  assign P32[26] = IN1[26]&IN2[6];
  assign P33[26] = IN1[26]&IN2[7];
  assign P34[26] = IN1[26]&IN2[8];
  assign P35[26] = IN1[26]&IN2[9];
  assign P36[26] = IN1[26]&IN2[10];
  assign P37[26] = IN1[26]&IN2[11];
  assign P38[26] = IN1[26]&IN2[12];
  assign P39[26] = IN1[26]&IN2[13];
  assign P40[26] = IN1[26]&IN2[14];
  assign P41[26] = IN1[26]&IN2[15];
  assign P42[26] = IN1[26]&IN2[16];
  assign P43[26] = IN1[26]&IN2[17];
  assign P44[26] = IN1[26]&IN2[18];
  assign P45[26] = IN1[26]&IN2[19];
  assign P46[26] = IN1[26]&IN2[20];
  assign P47[26] = IN1[26]&IN2[21];
  assign P48[26] = IN1[26]&IN2[22];
  assign P49[26] = IN1[26]&IN2[23];
  assign P50[26] = IN1[26]&IN2[24];
  assign P51[26] = IN1[26]&IN2[25];
  assign P52[26] = IN1[26]&IN2[26];
  assign P53[26] = IN1[26]&IN2[27];
  assign P54[25] = IN1[26]&IN2[28];
  assign P55[24] = IN1[26]&IN2[29];
  assign P56[23] = IN1[26]&IN2[30];
  assign P57[22] = IN1[26]&IN2[31];
  assign P58[21] = IN1[26]&IN2[32];
  assign P59[20] = IN1[26]&IN2[33];
  assign P60[19] = IN1[26]&IN2[34];
  assign P61[18] = IN1[26]&IN2[35];
  assign P62[17] = IN1[26]&IN2[36];
  assign P63[16] = IN1[26]&IN2[37];
  assign P64[15] = IN1[26]&IN2[38];
  assign P65[14] = IN1[26]&IN2[39];
  assign P66[13] = IN1[26]&IN2[40];
  assign P67[12] = IN1[26]&IN2[41];
  assign P68[11] = IN1[26]&IN2[42];
  assign P69[10] = IN1[26]&IN2[43];
  assign P70[9] = IN1[26]&IN2[44];
  assign P71[8] = IN1[26]&IN2[45];
  assign P72[7] = IN1[26]&IN2[46];
  assign P73[6] = IN1[26]&IN2[47];
  assign P74[5] = IN1[26]&IN2[48];
  assign P75[4] = IN1[26]&IN2[49];
  assign P76[3] = IN1[26]&IN2[50];
  assign P77[2] = IN1[26]&IN2[51];
  assign P78[1] = IN1[26]&IN2[52];
  assign P79[0] = IN1[26]&IN2[53];
  assign P27[27] = IN1[27]&IN2[0];
  assign P28[27] = IN1[27]&IN2[1];
  assign P29[27] = IN1[27]&IN2[2];
  assign P30[27] = IN1[27]&IN2[3];
  assign P31[27] = IN1[27]&IN2[4];
  assign P32[27] = IN1[27]&IN2[5];
  assign P33[27] = IN1[27]&IN2[6];
  assign P34[27] = IN1[27]&IN2[7];
  assign P35[27] = IN1[27]&IN2[8];
  assign P36[27] = IN1[27]&IN2[9];
  assign P37[27] = IN1[27]&IN2[10];
  assign P38[27] = IN1[27]&IN2[11];
  assign P39[27] = IN1[27]&IN2[12];
  assign P40[27] = IN1[27]&IN2[13];
  assign P41[27] = IN1[27]&IN2[14];
  assign P42[27] = IN1[27]&IN2[15];
  assign P43[27] = IN1[27]&IN2[16];
  assign P44[27] = IN1[27]&IN2[17];
  assign P45[27] = IN1[27]&IN2[18];
  assign P46[27] = IN1[27]&IN2[19];
  assign P47[27] = IN1[27]&IN2[20];
  assign P48[27] = IN1[27]&IN2[21];
  assign P49[27] = IN1[27]&IN2[22];
  assign P50[27] = IN1[27]&IN2[23];
  assign P51[27] = IN1[27]&IN2[24];
  assign P52[27] = IN1[27]&IN2[25];
  assign P53[27] = IN1[27]&IN2[26];
  assign P54[26] = IN1[27]&IN2[27];
  assign P55[25] = IN1[27]&IN2[28];
  assign P56[24] = IN1[27]&IN2[29];
  assign P57[23] = IN1[27]&IN2[30];
  assign P58[22] = IN1[27]&IN2[31];
  assign P59[21] = IN1[27]&IN2[32];
  assign P60[20] = IN1[27]&IN2[33];
  assign P61[19] = IN1[27]&IN2[34];
  assign P62[18] = IN1[27]&IN2[35];
  assign P63[17] = IN1[27]&IN2[36];
  assign P64[16] = IN1[27]&IN2[37];
  assign P65[15] = IN1[27]&IN2[38];
  assign P66[14] = IN1[27]&IN2[39];
  assign P67[13] = IN1[27]&IN2[40];
  assign P68[12] = IN1[27]&IN2[41];
  assign P69[11] = IN1[27]&IN2[42];
  assign P70[10] = IN1[27]&IN2[43];
  assign P71[9] = IN1[27]&IN2[44];
  assign P72[8] = IN1[27]&IN2[45];
  assign P73[7] = IN1[27]&IN2[46];
  assign P74[6] = IN1[27]&IN2[47];
  assign P75[5] = IN1[27]&IN2[48];
  assign P76[4] = IN1[27]&IN2[49];
  assign P77[3] = IN1[27]&IN2[50];
  assign P78[2] = IN1[27]&IN2[51];
  assign P79[1] = IN1[27]&IN2[52];
  assign P80[0] = IN1[27]&IN2[53];
  assign P28[28] = IN1[28]&IN2[0];
  assign P29[28] = IN1[28]&IN2[1];
  assign P30[28] = IN1[28]&IN2[2];
  assign P31[28] = IN1[28]&IN2[3];
  assign P32[28] = IN1[28]&IN2[4];
  assign P33[28] = IN1[28]&IN2[5];
  assign P34[28] = IN1[28]&IN2[6];
  assign P35[28] = IN1[28]&IN2[7];
  assign P36[28] = IN1[28]&IN2[8];
  assign P37[28] = IN1[28]&IN2[9];
  assign P38[28] = IN1[28]&IN2[10];
  assign P39[28] = IN1[28]&IN2[11];
  assign P40[28] = IN1[28]&IN2[12];
  assign P41[28] = IN1[28]&IN2[13];
  assign P42[28] = IN1[28]&IN2[14];
  assign P43[28] = IN1[28]&IN2[15];
  assign P44[28] = IN1[28]&IN2[16];
  assign P45[28] = IN1[28]&IN2[17];
  assign P46[28] = IN1[28]&IN2[18];
  assign P47[28] = IN1[28]&IN2[19];
  assign P48[28] = IN1[28]&IN2[20];
  assign P49[28] = IN1[28]&IN2[21];
  assign P50[28] = IN1[28]&IN2[22];
  assign P51[28] = IN1[28]&IN2[23];
  assign P52[28] = IN1[28]&IN2[24];
  assign P53[28] = IN1[28]&IN2[25];
  assign P54[27] = IN1[28]&IN2[26];
  assign P55[26] = IN1[28]&IN2[27];
  assign P56[25] = IN1[28]&IN2[28];
  assign P57[24] = IN1[28]&IN2[29];
  assign P58[23] = IN1[28]&IN2[30];
  assign P59[22] = IN1[28]&IN2[31];
  assign P60[21] = IN1[28]&IN2[32];
  assign P61[20] = IN1[28]&IN2[33];
  assign P62[19] = IN1[28]&IN2[34];
  assign P63[18] = IN1[28]&IN2[35];
  assign P64[17] = IN1[28]&IN2[36];
  assign P65[16] = IN1[28]&IN2[37];
  assign P66[15] = IN1[28]&IN2[38];
  assign P67[14] = IN1[28]&IN2[39];
  assign P68[13] = IN1[28]&IN2[40];
  assign P69[12] = IN1[28]&IN2[41];
  assign P70[11] = IN1[28]&IN2[42];
  assign P71[10] = IN1[28]&IN2[43];
  assign P72[9] = IN1[28]&IN2[44];
  assign P73[8] = IN1[28]&IN2[45];
  assign P74[7] = IN1[28]&IN2[46];
  assign P75[6] = IN1[28]&IN2[47];
  assign P76[5] = IN1[28]&IN2[48];
  assign P77[4] = IN1[28]&IN2[49];
  assign P78[3] = IN1[28]&IN2[50];
  assign P79[2] = IN1[28]&IN2[51];
  assign P80[1] = IN1[28]&IN2[52];
  assign P81[0] = IN1[28]&IN2[53];
  assign P29[29] = IN1[29]&IN2[0];
  assign P30[29] = IN1[29]&IN2[1];
  assign P31[29] = IN1[29]&IN2[2];
  assign P32[29] = IN1[29]&IN2[3];
  assign P33[29] = IN1[29]&IN2[4];
  assign P34[29] = IN1[29]&IN2[5];
  assign P35[29] = IN1[29]&IN2[6];
  assign P36[29] = IN1[29]&IN2[7];
  assign P37[29] = IN1[29]&IN2[8];
  assign P38[29] = IN1[29]&IN2[9];
  assign P39[29] = IN1[29]&IN2[10];
  assign P40[29] = IN1[29]&IN2[11];
  assign P41[29] = IN1[29]&IN2[12];
  assign P42[29] = IN1[29]&IN2[13];
  assign P43[29] = IN1[29]&IN2[14];
  assign P44[29] = IN1[29]&IN2[15];
  assign P45[29] = IN1[29]&IN2[16];
  assign P46[29] = IN1[29]&IN2[17];
  assign P47[29] = IN1[29]&IN2[18];
  assign P48[29] = IN1[29]&IN2[19];
  assign P49[29] = IN1[29]&IN2[20];
  assign P50[29] = IN1[29]&IN2[21];
  assign P51[29] = IN1[29]&IN2[22];
  assign P52[29] = IN1[29]&IN2[23];
  assign P53[29] = IN1[29]&IN2[24];
  assign P54[28] = IN1[29]&IN2[25];
  assign P55[27] = IN1[29]&IN2[26];
  assign P56[26] = IN1[29]&IN2[27];
  assign P57[25] = IN1[29]&IN2[28];
  assign P58[24] = IN1[29]&IN2[29];
  assign P59[23] = IN1[29]&IN2[30];
  assign P60[22] = IN1[29]&IN2[31];
  assign P61[21] = IN1[29]&IN2[32];
  assign P62[20] = IN1[29]&IN2[33];
  assign P63[19] = IN1[29]&IN2[34];
  assign P64[18] = IN1[29]&IN2[35];
  assign P65[17] = IN1[29]&IN2[36];
  assign P66[16] = IN1[29]&IN2[37];
  assign P67[15] = IN1[29]&IN2[38];
  assign P68[14] = IN1[29]&IN2[39];
  assign P69[13] = IN1[29]&IN2[40];
  assign P70[12] = IN1[29]&IN2[41];
  assign P71[11] = IN1[29]&IN2[42];
  assign P72[10] = IN1[29]&IN2[43];
  assign P73[9] = IN1[29]&IN2[44];
  assign P74[8] = IN1[29]&IN2[45];
  assign P75[7] = IN1[29]&IN2[46];
  assign P76[6] = IN1[29]&IN2[47];
  assign P77[5] = IN1[29]&IN2[48];
  assign P78[4] = IN1[29]&IN2[49];
  assign P79[3] = IN1[29]&IN2[50];
  assign P80[2] = IN1[29]&IN2[51];
  assign P81[1] = IN1[29]&IN2[52];
  assign P82[0] = IN1[29]&IN2[53];
  assign P30[30] = IN1[30]&IN2[0];
  assign P31[30] = IN1[30]&IN2[1];
  assign P32[30] = IN1[30]&IN2[2];
  assign P33[30] = IN1[30]&IN2[3];
  assign P34[30] = IN1[30]&IN2[4];
  assign P35[30] = IN1[30]&IN2[5];
  assign P36[30] = IN1[30]&IN2[6];
  assign P37[30] = IN1[30]&IN2[7];
  assign P38[30] = IN1[30]&IN2[8];
  assign P39[30] = IN1[30]&IN2[9];
  assign P40[30] = IN1[30]&IN2[10];
  assign P41[30] = IN1[30]&IN2[11];
  assign P42[30] = IN1[30]&IN2[12];
  assign P43[30] = IN1[30]&IN2[13];
  assign P44[30] = IN1[30]&IN2[14];
  assign P45[30] = IN1[30]&IN2[15];
  assign P46[30] = IN1[30]&IN2[16];
  assign P47[30] = IN1[30]&IN2[17];
  assign P48[30] = IN1[30]&IN2[18];
  assign P49[30] = IN1[30]&IN2[19];
  assign P50[30] = IN1[30]&IN2[20];
  assign P51[30] = IN1[30]&IN2[21];
  assign P52[30] = IN1[30]&IN2[22];
  assign P53[30] = IN1[30]&IN2[23];
  assign P54[29] = IN1[30]&IN2[24];
  assign P55[28] = IN1[30]&IN2[25];
  assign P56[27] = IN1[30]&IN2[26];
  assign P57[26] = IN1[30]&IN2[27];
  assign P58[25] = IN1[30]&IN2[28];
  assign P59[24] = IN1[30]&IN2[29];
  assign P60[23] = IN1[30]&IN2[30];
  assign P61[22] = IN1[30]&IN2[31];
  assign P62[21] = IN1[30]&IN2[32];
  assign P63[20] = IN1[30]&IN2[33];
  assign P64[19] = IN1[30]&IN2[34];
  assign P65[18] = IN1[30]&IN2[35];
  assign P66[17] = IN1[30]&IN2[36];
  assign P67[16] = IN1[30]&IN2[37];
  assign P68[15] = IN1[30]&IN2[38];
  assign P69[14] = IN1[30]&IN2[39];
  assign P70[13] = IN1[30]&IN2[40];
  assign P71[12] = IN1[30]&IN2[41];
  assign P72[11] = IN1[30]&IN2[42];
  assign P73[10] = IN1[30]&IN2[43];
  assign P74[9] = IN1[30]&IN2[44];
  assign P75[8] = IN1[30]&IN2[45];
  assign P76[7] = IN1[30]&IN2[46];
  assign P77[6] = IN1[30]&IN2[47];
  assign P78[5] = IN1[30]&IN2[48];
  assign P79[4] = IN1[30]&IN2[49];
  assign P80[3] = IN1[30]&IN2[50];
  assign P81[2] = IN1[30]&IN2[51];
  assign P82[1] = IN1[30]&IN2[52];
  assign P83[0] = IN1[30]&IN2[53];
  assign P31[31] = IN1[31]&IN2[0];
  assign P32[31] = IN1[31]&IN2[1];
  assign P33[31] = IN1[31]&IN2[2];
  assign P34[31] = IN1[31]&IN2[3];
  assign P35[31] = IN1[31]&IN2[4];
  assign P36[31] = IN1[31]&IN2[5];
  assign P37[31] = IN1[31]&IN2[6];
  assign P38[31] = IN1[31]&IN2[7];
  assign P39[31] = IN1[31]&IN2[8];
  assign P40[31] = IN1[31]&IN2[9];
  assign P41[31] = IN1[31]&IN2[10];
  assign P42[31] = IN1[31]&IN2[11];
  assign P43[31] = IN1[31]&IN2[12];
  assign P44[31] = IN1[31]&IN2[13];
  assign P45[31] = IN1[31]&IN2[14];
  assign P46[31] = IN1[31]&IN2[15];
  assign P47[31] = IN1[31]&IN2[16];
  assign P48[31] = IN1[31]&IN2[17];
  assign P49[31] = IN1[31]&IN2[18];
  assign P50[31] = IN1[31]&IN2[19];
  assign P51[31] = IN1[31]&IN2[20];
  assign P52[31] = IN1[31]&IN2[21];
  assign P53[31] = IN1[31]&IN2[22];
  assign P54[30] = IN1[31]&IN2[23];
  assign P55[29] = IN1[31]&IN2[24];
  assign P56[28] = IN1[31]&IN2[25];
  assign P57[27] = IN1[31]&IN2[26];
  assign P58[26] = IN1[31]&IN2[27];
  assign P59[25] = IN1[31]&IN2[28];
  assign P60[24] = IN1[31]&IN2[29];
  assign P61[23] = IN1[31]&IN2[30];
  assign P62[22] = IN1[31]&IN2[31];
  assign P63[21] = IN1[31]&IN2[32];
  assign P64[20] = IN1[31]&IN2[33];
  assign P65[19] = IN1[31]&IN2[34];
  assign P66[18] = IN1[31]&IN2[35];
  assign P67[17] = IN1[31]&IN2[36];
  assign P68[16] = IN1[31]&IN2[37];
  assign P69[15] = IN1[31]&IN2[38];
  assign P70[14] = IN1[31]&IN2[39];
  assign P71[13] = IN1[31]&IN2[40];
  assign P72[12] = IN1[31]&IN2[41];
  assign P73[11] = IN1[31]&IN2[42];
  assign P74[10] = IN1[31]&IN2[43];
  assign P75[9] = IN1[31]&IN2[44];
  assign P76[8] = IN1[31]&IN2[45];
  assign P77[7] = IN1[31]&IN2[46];
  assign P78[6] = IN1[31]&IN2[47];
  assign P79[5] = IN1[31]&IN2[48];
  assign P80[4] = IN1[31]&IN2[49];
  assign P81[3] = IN1[31]&IN2[50];
  assign P82[2] = IN1[31]&IN2[51];
  assign P83[1] = IN1[31]&IN2[52];
  assign P84[0] = IN1[31]&IN2[53];
  assign P32[32] = IN1[32]&IN2[0];
  assign P33[32] = IN1[32]&IN2[1];
  assign P34[32] = IN1[32]&IN2[2];
  assign P35[32] = IN1[32]&IN2[3];
  assign P36[32] = IN1[32]&IN2[4];
  assign P37[32] = IN1[32]&IN2[5];
  assign P38[32] = IN1[32]&IN2[6];
  assign P39[32] = IN1[32]&IN2[7];
  assign P40[32] = IN1[32]&IN2[8];
  assign P41[32] = IN1[32]&IN2[9];
  assign P42[32] = IN1[32]&IN2[10];
  assign P43[32] = IN1[32]&IN2[11];
  assign P44[32] = IN1[32]&IN2[12];
  assign P45[32] = IN1[32]&IN2[13];
  assign P46[32] = IN1[32]&IN2[14];
  assign P47[32] = IN1[32]&IN2[15];
  assign P48[32] = IN1[32]&IN2[16];
  assign P49[32] = IN1[32]&IN2[17];
  assign P50[32] = IN1[32]&IN2[18];
  assign P51[32] = IN1[32]&IN2[19];
  assign P52[32] = IN1[32]&IN2[20];
  assign P53[32] = IN1[32]&IN2[21];
  assign P54[31] = IN1[32]&IN2[22];
  assign P55[30] = IN1[32]&IN2[23];
  assign P56[29] = IN1[32]&IN2[24];
  assign P57[28] = IN1[32]&IN2[25];
  assign P58[27] = IN1[32]&IN2[26];
  assign P59[26] = IN1[32]&IN2[27];
  assign P60[25] = IN1[32]&IN2[28];
  assign P61[24] = IN1[32]&IN2[29];
  assign P62[23] = IN1[32]&IN2[30];
  assign P63[22] = IN1[32]&IN2[31];
  assign P64[21] = IN1[32]&IN2[32];
  assign P65[20] = IN1[32]&IN2[33];
  assign P66[19] = IN1[32]&IN2[34];
  assign P67[18] = IN1[32]&IN2[35];
  assign P68[17] = IN1[32]&IN2[36];
  assign P69[16] = IN1[32]&IN2[37];
  assign P70[15] = IN1[32]&IN2[38];
  assign P71[14] = IN1[32]&IN2[39];
  assign P72[13] = IN1[32]&IN2[40];
  assign P73[12] = IN1[32]&IN2[41];
  assign P74[11] = IN1[32]&IN2[42];
  assign P75[10] = IN1[32]&IN2[43];
  assign P76[9] = IN1[32]&IN2[44];
  assign P77[8] = IN1[32]&IN2[45];
  assign P78[7] = IN1[32]&IN2[46];
  assign P79[6] = IN1[32]&IN2[47];
  assign P80[5] = IN1[32]&IN2[48];
  assign P81[4] = IN1[32]&IN2[49];
  assign P82[3] = IN1[32]&IN2[50];
  assign P83[2] = IN1[32]&IN2[51];
  assign P84[1] = IN1[32]&IN2[52];
  assign P85[0] = IN1[32]&IN2[53];
  assign P33[33] = IN1[33]&IN2[0];
  assign P34[33] = IN1[33]&IN2[1];
  assign P35[33] = IN1[33]&IN2[2];
  assign P36[33] = IN1[33]&IN2[3];
  assign P37[33] = IN1[33]&IN2[4];
  assign P38[33] = IN1[33]&IN2[5];
  assign P39[33] = IN1[33]&IN2[6];
  assign P40[33] = IN1[33]&IN2[7];
  assign P41[33] = IN1[33]&IN2[8];
  assign P42[33] = IN1[33]&IN2[9];
  assign P43[33] = IN1[33]&IN2[10];
  assign P44[33] = IN1[33]&IN2[11];
  assign P45[33] = IN1[33]&IN2[12];
  assign P46[33] = IN1[33]&IN2[13];
  assign P47[33] = IN1[33]&IN2[14];
  assign P48[33] = IN1[33]&IN2[15];
  assign P49[33] = IN1[33]&IN2[16];
  assign P50[33] = IN1[33]&IN2[17];
  assign P51[33] = IN1[33]&IN2[18];
  assign P52[33] = IN1[33]&IN2[19];
  assign P53[33] = IN1[33]&IN2[20];
  assign P54[32] = IN1[33]&IN2[21];
  assign P55[31] = IN1[33]&IN2[22];
  assign P56[30] = IN1[33]&IN2[23];
  assign P57[29] = IN1[33]&IN2[24];
  assign P58[28] = IN1[33]&IN2[25];
  assign P59[27] = IN1[33]&IN2[26];
  assign P60[26] = IN1[33]&IN2[27];
  assign P61[25] = IN1[33]&IN2[28];
  assign P62[24] = IN1[33]&IN2[29];
  assign P63[23] = IN1[33]&IN2[30];
  assign P64[22] = IN1[33]&IN2[31];
  assign P65[21] = IN1[33]&IN2[32];
  assign P66[20] = IN1[33]&IN2[33];
  assign P67[19] = IN1[33]&IN2[34];
  assign P68[18] = IN1[33]&IN2[35];
  assign P69[17] = IN1[33]&IN2[36];
  assign P70[16] = IN1[33]&IN2[37];
  assign P71[15] = IN1[33]&IN2[38];
  assign P72[14] = IN1[33]&IN2[39];
  assign P73[13] = IN1[33]&IN2[40];
  assign P74[12] = IN1[33]&IN2[41];
  assign P75[11] = IN1[33]&IN2[42];
  assign P76[10] = IN1[33]&IN2[43];
  assign P77[9] = IN1[33]&IN2[44];
  assign P78[8] = IN1[33]&IN2[45];
  assign P79[7] = IN1[33]&IN2[46];
  assign P80[6] = IN1[33]&IN2[47];
  assign P81[5] = IN1[33]&IN2[48];
  assign P82[4] = IN1[33]&IN2[49];
  assign P83[3] = IN1[33]&IN2[50];
  assign P84[2] = IN1[33]&IN2[51];
  assign P85[1] = IN1[33]&IN2[52];
  assign P86[0] = IN1[33]&IN2[53];
  assign P34[34] = IN1[34]&IN2[0];
  assign P35[34] = IN1[34]&IN2[1];
  assign P36[34] = IN1[34]&IN2[2];
  assign P37[34] = IN1[34]&IN2[3];
  assign P38[34] = IN1[34]&IN2[4];
  assign P39[34] = IN1[34]&IN2[5];
  assign P40[34] = IN1[34]&IN2[6];
  assign P41[34] = IN1[34]&IN2[7];
  assign P42[34] = IN1[34]&IN2[8];
  assign P43[34] = IN1[34]&IN2[9];
  assign P44[34] = IN1[34]&IN2[10];
  assign P45[34] = IN1[34]&IN2[11];
  assign P46[34] = IN1[34]&IN2[12];
  assign P47[34] = IN1[34]&IN2[13];
  assign P48[34] = IN1[34]&IN2[14];
  assign P49[34] = IN1[34]&IN2[15];
  assign P50[34] = IN1[34]&IN2[16];
  assign P51[34] = IN1[34]&IN2[17];
  assign P52[34] = IN1[34]&IN2[18];
  assign P53[34] = IN1[34]&IN2[19];
  assign P54[33] = IN1[34]&IN2[20];
  assign P55[32] = IN1[34]&IN2[21];
  assign P56[31] = IN1[34]&IN2[22];
  assign P57[30] = IN1[34]&IN2[23];
  assign P58[29] = IN1[34]&IN2[24];
  assign P59[28] = IN1[34]&IN2[25];
  assign P60[27] = IN1[34]&IN2[26];
  assign P61[26] = IN1[34]&IN2[27];
  assign P62[25] = IN1[34]&IN2[28];
  assign P63[24] = IN1[34]&IN2[29];
  assign P64[23] = IN1[34]&IN2[30];
  assign P65[22] = IN1[34]&IN2[31];
  assign P66[21] = IN1[34]&IN2[32];
  assign P67[20] = IN1[34]&IN2[33];
  assign P68[19] = IN1[34]&IN2[34];
  assign P69[18] = IN1[34]&IN2[35];
  assign P70[17] = IN1[34]&IN2[36];
  assign P71[16] = IN1[34]&IN2[37];
  assign P72[15] = IN1[34]&IN2[38];
  assign P73[14] = IN1[34]&IN2[39];
  assign P74[13] = IN1[34]&IN2[40];
  assign P75[12] = IN1[34]&IN2[41];
  assign P76[11] = IN1[34]&IN2[42];
  assign P77[10] = IN1[34]&IN2[43];
  assign P78[9] = IN1[34]&IN2[44];
  assign P79[8] = IN1[34]&IN2[45];
  assign P80[7] = IN1[34]&IN2[46];
  assign P81[6] = IN1[34]&IN2[47];
  assign P82[5] = IN1[34]&IN2[48];
  assign P83[4] = IN1[34]&IN2[49];
  assign P84[3] = IN1[34]&IN2[50];
  assign P85[2] = IN1[34]&IN2[51];
  assign P86[1] = IN1[34]&IN2[52];
  assign P87[0] = IN1[34]&IN2[53];
  assign P35[35] = IN1[35]&IN2[0];
  assign P36[35] = IN1[35]&IN2[1];
  assign P37[35] = IN1[35]&IN2[2];
  assign P38[35] = IN1[35]&IN2[3];
  assign P39[35] = IN1[35]&IN2[4];
  assign P40[35] = IN1[35]&IN2[5];
  assign P41[35] = IN1[35]&IN2[6];
  assign P42[35] = IN1[35]&IN2[7];
  assign P43[35] = IN1[35]&IN2[8];
  assign P44[35] = IN1[35]&IN2[9];
  assign P45[35] = IN1[35]&IN2[10];
  assign P46[35] = IN1[35]&IN2[11];
  assign P47[35] = IN1[35]&IN2[12];
  assign P48[35] = IN1[35]&IN2[13];
  assign P49[35] = IN1[35]&IN2[14];
  assign P50[35] = IN1[35]&IN2[15];
  assign P51[35] = IN1[35]&IN2[16];
  assign P52[35] = IN1[35]&IN2[17];
  assign P53[35] = IN1[35]&IN2[18];
  assign P54[34] = IN1[35]&IN2[19];
  assign P55[33] = IN1[35]&IN2[20];
  assign P56[32] = IN1[35]&IN2[21];
  assign P57[31] = IN1[35]&IN2[22];
  assign P58[30] = IN1[35]&IN2[23];
  assign P59[29] = IN1[35]&IN2[24];
  assign P60[28] = IN1[35]&IN2[25];
  assign P61[27] = IN1[35]&IN2[26];
  assign P62[26] = IN1[35]&IN2[27];
  assign P63[25] = IN1[35]&IN2[28];
  assign P64[24] = IN1[35]&IN2[29];
  assign P65[23] = IN1[35]&IN2[30];
  assign P66[22] = IN1[35]&IN2[31];
  assign P67[21] = IN1[35]&IN2[32];
  assign P68[20] = IN1[35]&IN2[33];
  assign P69[19] = IN1[35]&IN2[34];
  assign P70[18] = IN1[35]&IN2[35];
  assign P71[17] = IN1[35]&IN2[36];
  assign P72[16] = IN1[35]&IN2[37];
  assign P73[15] = IN1[35]&IN2[38];
  assign P74[14] = IN1[35]&IN2[39];
  assign P75[13] = IN1[35]&IN2[40];
  assign P76[12] = IN1[35]&IN2[41];
  assign P77[11] = IN1[35]&IN2[42];
  assign P78[10] = IN1[35]&IN2[43];
  assign P79[9] = IN1[35]&IN2[44];
  assign P80[8] = IN1[35]&IN2[45];
  assign P81[7] = IN1[35]&IN2[46];
  assign P82[6] = IN1[35]&IN2[47];
  assign P83[5] = IN1[35]&IN2[48];
  assign P84[4] = IN1[35]&IN2[49];
  assign P85[3] = IN1[35]&IN2[50];
  assign P86[2] = IN1[35]&IN2[51];
  assign P87[1] = IN1[35]&IN2[52];
  assign P88[0] = IN1[35]&IN2[53];
  assign P36[36] = IN1[36]&IN2[0];
  assign P37[36] = IN1[36]&IN2[1];
  assign P38[36] = IN1[36]&IN2[2];
  assign P39[36] = IN1[36]&IN2[3];
  assign P40[36] = IN1[36]&IN2[4];
  assign P41[36] = IN1[36]&IN2[5];
  assign P42[36] = IN1[36]&IN2[6];
  assign P43[36] = IN1[36]&IN2[7];
  assign P44[36] = IN1[36]&IN2[8];
  assign P45[36] = IN1[36]&IN2[9];
  assign P46[36] = IN1[36]&IN2[10];
  assign P47[36] = IN1[36]&IN2[11];
  assign P48[36] = IN1[36]&IN2[12];
  assign P49[36] = IN1[36]&IN2[13];
  assign P50[36] = IN1[36]&IN2[14];
  assign P51[36] = IN1[36]&IN2[15];
  assign P52[36] = IN1[36]&IN2[16];
  assign P53[36] = IN1[36]&IN2[17];
  assign P54[35] = IN1[36]&IN2[18];
  assign P55[34] = IN1[36]&IN2[19];
  assign P56[33] = IN1[36]&IN2[20];
  assign P57[32] = IN1[36]&IN2[21];
  assign P58[31] = IN1[36]&IN2[22];
  assign P59[30] = IN1[36]&IN2[23];
  assign P60[29] = IN1[36]&IN2[24];
  assign P61[28] = IN1[36]&IN2[25];
  assign P62[27] = IN1[36]&IN2[26];
  assign P63[26] = IN1[36]&IN2[27];
  assign P64[25] = IN1[36]&IN2[28];
  assign P65[24] = IN1[36]&IN2[29];
  assign P66[23] = IN1[36]&IN2[30];
  assign P67[22] = IN1[36]&IN2[31];
  assign P68[21] = IN1[36]&IN2[32];
  assign P69[20] = IN1[36]&IN2[33];
  assign P70[19] = IN1[36]&IN2[34];
  assign P71[18] = IN1[36]&IN2[35];
  assign P72[17] = IN1[36]&IN2[36];
  assign P73[16] = IN1[36]&IN2[37];
  assign P74[15] = IN1[36]&IN2[38];
  assign P75[14] = IN1[36]&IN2[39];
  assign P76[13] = IN1[36]&IN2[40];
  assign P77[12] = IN1[36]&IN2[41];
  assign P78[11] = IN1[36]&IN2[42];
  assign P79[10] = IN1[36]&IN2[43];
  assign P80[9] = IN1[36]&IN2[44];
  assign P81[8] = IN1[36]&IN2[45];
  assign P82[7] = IN1[36]&IN2[46];
  assign P83[6] = IN1[36]&IN2[47];
  assign P84[5] = IN1[36]&IN2[48];
  assign P85[4] = IN1[36]&IN2[49];
  assign P86[3] = IN1[36]&IN2[50];
  assign P87[2] = IN1[36]&IN2[51];
  assign P88[1] = IN1[36]&IN2[52];
  assign P89[0] = IN1[36]&IN2[53];
  assign P37[37] = IN1[37]&IN2[0];
  assign P38[37] = IN1[37]&IN2[1];
  assign P39[37] = IN1[37]&IN2[2];
  assign P40[37] = IN1[37]&IN2[3];
  assign P41[37] = IN1[37]&IN2[4];
  assign P42[37] = IN1[37]&IN2[5];
  assign P43[37] = IN1[37]&IN2[6];
  assign P44[37] = IN1[37]&IN2[7];
  assign P45[37] = IN1[37]&IN2[8];
  assign P46[37] = IN1[37]&IN2[9];
  assign P47[37] = IN1[37]&IN2[10];
  assign P48[37] = IN1[37]&IN2[11];
  assign P49[37] = IN1[37]&IN2[12];
  assign P50[37] = IN1[37]&IN2[13];
  assign P51[37] = IN1[37]&IN2[14];
  assign P52[37] = IN1[37]&IN2[15];
  assign P53[37] = IN1[37]&IN2[16];
  assign P54[36] = IN1[37]&IN2[17];
  assign P55[35] = IN1[37]&IN2[18];
  assign P56[34] = IN1[37]&IN2[19];
  assign P57[33] = IN1[37]&IN2[20];
  assign P58[32] = IN1[37]&IN2[21];
  assign P59[31] = IN1[37]&IN2[22];
  assign P60[30] = IN1[37]&IN2[23];
  assign P61[29] = IN1[37]&IN2[24];
  assign P62[28] = IN1[37]&IN2[25];
  assign P63[27] = IN1[37]&IN2[26];
  assign P64[26] = IN1[37]&IN2[27];
  assign P65[25] = IN1[37]&IN2[28];
  assign P66[24] = IN1[37]&IN2[29];
  assign P67[23] = IN1[37]&IN2[30];
  assign P68[22] = IN1[37]&IN2[31];
  assign P69[21] = IN1[37]&IN2[32];
  assign P70[20] = IN1[37]&IN2[33];
  assign P71[19] = IN1[37]&IN2[34];
  assign P72[18] = IN1[37]&IN2[35];
  assign P73[17] = IN1[37]&IN2[36];
  assign P74[16] = IN1[37]&IN2[37];
  assign P75[15] = IN1[37]&IN2[38];
  assign P76[14] = IN1[37]&IN2[39];
  assign P77[13] = IN1[37]&IN2[40];
  assign P78[12] = IN1[37]&IN2[41];
  assign P79[11] = IN1[37]&IN2[42];
  assign P80[10] = IN1[37]&IN2[43];
  assign P81[9] = IN1[37]&IN2[44];
  assign P82[8] = IN1[37]&IN2[45];
  assign P83[7] = IN1[37]&IN2[46];
  assign P84[6] = IN1[37]&IN2[47];
  assign P85[5] = IN1[37]&IN2[48];
  assign P86[4] = IN1[37]&IN2[49];
  assign P87[3] = IN1[37]&IN2[50];
  assign P88[2] = IN1[37]&IN2[51];
  assign P89[1] = IN1[37]&IN2[52];
  assign P90[0] = IN1[37]&IN2[53];
  assign P38[38] = IN1[38]&IN2[0];
  assign P39[38] = IN1[38]&IN2[1];
  assign P40[38] = IN1[38]&IN2[2];
  assign P41[38] = IN1[38]&IN2[3];
  assign P42[38] = IN1[38]&IN2[4];
  assign P43[38] = IN1[38]&IN2[5];
  assign P44[38] = IN1[38]&IN2[6];
  assign P45[38] = IN1[38]&IN2[7];
  assign P46[38] = IN1[38]&IN2[8];
  assign P47[38] = IN1[38]&IN2[9];
  assign P48[38] = IN1[38]&IN2[10];
  assign P49[38] = IN1[38]&IN2[11];
  assign P50[38] = IN1[38]&IN2[12];
  assign P51[38] = IN1[38]&IN2[13];
  assign P52[38] = IN1[38]&IN2[14];
  assign P53[38] = IN1[38]&IN2[15];
  assign P54[37] = IN1[38]&IN2[16];
  assign P55[36] = IN1[38]&IN2[17];
  assign P56[35] = IN1[38]&IN2[18];
  assign P57[34] = IN1[38]&IN2[19];
  assign P58[33] = IN1[38]&IN2[20];
  assign P59[32] = IN1[38]&IN2[21];
  assign P60[31] = IN1[38]&IN2[22];
  assign P61[30] = IN1[38]&IN2[23];
  assign P62[29] = IN1[38]&IN2[24];
  assign P63[28] = IN1[38]&IN2[25];
  assign P64[27] = IN1[38]&IN2[26];
  assign P65[26] = IN1[38]&IN2[27];
  assign P66[25] = IN1[38]&IN2[28];
  assign P67[24] = IN1[38]&IN2[29];
  assign P68[23] = IN1[38]&IN2[30];
  assign P69[22] = IN1[38]&IN2[31];
  assign P70[21] = IN1[38]&IN2[32];
  assign P71[20] = IN1[38]&IN2[33];
  assign P72[19] = IN1[38]&IN2[34];
  assign P73[18] = IN1[38]&IN2[35];
  assign P74[17] = IN1[38]&IN2[36];
  assign P75[16] = IN1[38]&IN2[37];
  assign P76[15] = IN1[38]&IN2[38];
  assign P77[14] = IN1[38]&IN2[39];
  assign P78[13] = IN1[38]&IN2[40];
  assign P79[12] = IN1[38]&IN2[41];
  assign P80[11] = IN1[38]&IN2[42];
  assign P81[10] = IN1[38]&IN2[43];
  assign P82[9] = IN1[38]&IN2[44];
  assign P83[8] = IN1[38]&IN2[45];
  assign P84[7] = IN1[38]&IN2[46];
  assign P85[6] = IN1[38]&IN2[47];
  assign P86[5] = IN1[38]&IN2[48];
  assign P87[4] = IN1[38]&IN2[49];
  assign P88[3] = IN1[38]&IN2[50];
  assign P89[2] = IN1[38]&IN2[51];
  assign P90[1] = IN1[38]&IN2[52];
  assign P91[0] = IN1[38]&IN2[53];
  assign P39[39] = IN1[39]&IN2[0];
  assign P40[39] = IN1[39]&IN2[1];
  assign P41[39] = IN1[39]&IN2[2];
  assign P42[39] = IN1[39]&IN2[3];
  assign P43[39] = IN1[39]&IN2[4];
  assign P44[39] = IN1[39]&IN2[5];
  assign P45[39] = IN1[39]&IN2[6];
  assign P46[39] = IN1[39]&IN2[7];
  assign P47[39] = IN1[39]&IN2[8];
  assign P48[39] = IN1[39]&IN2[9];
  assign P49[39] = IN1[39]&IN2[10];
  assign P50[39] = IN1[39]&IN2[11];
  assign P51[39] = IN1[39]&IN2[12];
  assign P52[39] = IN1[39]&IN2[13];
  assign P53[39] = IN1[39]&IN2[14];
  assign P54[38] = IN1[39]&IN2[15];
  assign P55[37] = IN1[39]&IN2[16];
  assign P56[36] = IN1[39]&IN2[17];
  assign P57[35] = IN1[39]&IN2[18];
  assign P58[34] = IN1[39]&IN2[19];
  assign P59[33] = IN1[39]&IN2[20];
  assign P60[32] = IN1[39]&IN2[21];
  assign P61[31] = IN1[39]&IN2[22];
  assign P62[30] = IN1[39]&IN2[23];
  assign P63[29] = IN1[39]&IN2[24];
  assign P64[28] = IN1[39]&IN2[25];
  assign P65[27] = IN1[39]&IN2[26];
  assign P66[26] = IN1[39]&IN2[27];
  assign P67[25] = IN1[39]&IN2[28];
  assign P68[24] = IN1[39]&IN2[29];
  assign P69[23] = IN1[39]&IN2[30];
  assign P70[22] = IN1[39]&IN2[31];
  assign P71[21] = IN1[39]&IN2[32];
  assign P72[20] = IN1[39]&IN2[33];
  assign P73[19] = IN1[39]&IN2[34];
  assign P74[18] = IN1[39]&IN2[35];
  assign P75[17] = IN1[39]&IN2[36];
  assign P76[16] = IN1[39]&IN2[37];
  assign P77[15] = IN1[39]&IN2[38];
  assign P78[14] = IN1[39]&IN2[39];
  assign P79[13] = IN1[39]&IN2[40];
  assign P80[12] = IN1[39]&IN2[41];
  assign P81[11] = IN1[39]&IN2[42];
  assign P82[10] = IN1[39]&IN2[43];
  assign P83[9] = IN1[39]&IN2[44];
  assign P84[8] = IN1[39]&IN2[45];
  assign P85[7] = IN1[39]&IN2[46];
  assign P86[6] = IN1[39]&IN2[47];
  assign P87[5] = IN1[39]&IN2[48];
  assign P88[4] = IN1[39]&IN2[49];
  assign P89[3] = IN1[39]&IN2[50];
  assign P90[2] = IN1[39]&IN2[51];
  assign P91[1] = IN1[39]&IN2[52];
  assign P92[0] = IN1[39]&IN2[53];
  assign P40[40] = IN1[40]&IN2[0];
  assign P41[40] = IN1[40]&IN2[1];
  assign P42[40] = IN1[40]&IN2[2];
  assign P43[40] = IN1[40]&IN2[3];
  assign P44[40] = IN1[40]&IN2[4];
  assign P45[40] = IN1[40]&IN2[5];
  assign P46[40] = IN1[40]&IN2[6];
  assign P47[40] = IN1[40]&IN2[7];
  assign P48[40] = IN1[40]&IN2[8];
  assign P49[40] = IN1[40]&IN2[9];
  assign P50[40] = IN1[40]&IN2[10];
  assign P51[40] = IN1[40]&IN2[11];
  assign P52[40] = IN1[40]&IN2[12];
  assign P53[40] = IN1[40]&IN2[13];
  assign P54[39] = IN1[40]&IN2[14];
  assign P55[38] = IN1[40]&IN2[15];
  assign P56[37] = IN1[40]&IN2[16];
  assign P57[36] = IN1[40]&IN2[17];
  assign P58[35] = IN1[40]&IN2[18];
  assign P59[34] = IN1[40]&IN2[19];
  assign P60[33] = IN1[40]&IN2[20];
  assign P61[32] = IN1[40]&IN2[21];
  assign P62[31] = IN1[40]&IN2[22];
  assign P63[30] = IN1[40]&IN2[23];
  assign P64[29] = IN1[40]&IN2[24];
  assign P65[28] = IN1[40]&IN2[25];
  assign P66[27] = IN1[40]&IN2[26];
  assign P67[26] = IN1[40]&IN2[27];
  assign P68[25] = IN1[40]&IN2[28];
  assign P69[24] = IN1[40]&IN2[29];
  assign P70[23] = IN1[40]&IN2[30];
  assign P71[22] = IN1[40]&IN2[31];
  assign P72[21] = IN1[40]&IN2[32];
  assign P73[20] = IN1[40]&IN2[33];
  assign P74[19] = IN1[40]&IN2[34];
  assign P75[18] = IN1[40]&IN2[35];
  assign P76[17] = IN1[40]&IN2[36];
  assign P77[16] = IN1[40]&IN2[37];
  assign P78[15] = IN1[40]&IN2[38];
  assign P79[14] = IN1[40]&IN2[39];
  assign P80[13] = IN1[40]&IN2[40];
  assign P81[12] = IN1[40]&IN2[41];
  assign P82[11] = IN1[40]&IN2[42];
  assign P83[10] = IN1[40]&IN2[43];
  assign P84[9] = IN1[40]&IN2[44];
  assign P85[8] = IN1[40]&IN2[45];
  assign P86[7] = IN1[40]&IN2[46];
  assign P87[6] = IN1[40]&IN2[47];
  assign P88[5] = IN1[40]&IN2[48];
  assign P89[4] = IN1[40]&IN2[49];
  assign P90[3] = IN1[40]&IN2[50];
  assign P91[2] = IN1[40]&IN2[51];
  assign P92[1] = IN1[40]&IN2[52];
  assign P93[0] = IN1[40]&IN2[53];

endmodule
module AR(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, IN31, IN32, IN33, IN34, IN35, IN36, IN37, IN38, IN39, IN40, IN41, IN42, IN43, IN44, IN45, IN46, IN47, IN48, IN49, IN50, IN51, IN52, IN53, IN54, IN55, IN56, IN57, IN58, IN59, IN60, IN61, IN62, IN63, IN64, IN65, IN66, IN67, IN68, IN69, IN70, IN71, IN72, IN73, IN74, IN75, IN76, IN77, IN78, IN79, IN80, IN81, IN82, IN83, IN84, IN85, IN86, IN87, IN88, IN89, IN90, IN91, IN92, IN93, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [16:0] IN16;
  input [17:0] IN17;
  input [18:0] IN18;
  input [19:0] IN19;
  input [20:0] IN20;
  input [21:0] IN21;
  input [22:0] IN22;
  input [23:0] IN23;
  input [24:0] IN24;
  input [25:0] IN25;
  input [26:0] IN26;
  input [27:0] IN27;
  input [28:0] IN28;
  input [29:0] IN29;
  input [30:0] IN30;
  input [31:0] IN31;
  input [32:0] IN32;
  input [33:0] IN33;
  input [34:0] IN34;
  input [35:0] IN35;
  input [36:0] IN36;
  input [37:0] IN37;
  input [38:0] IN38;
  input [39:0] IN39;
  input [40:0] IN40;
  input [40:0] IN41;
  input [40:0] IN42;
  input [40:0] IN43;
  input [40:0] IN44;
  input [40:0] IN45;
  input [40:0] IN46;
  input [40:0] IN47;
  input [40:0] IN48;
  input [40:0] IN49;
  input [40:0] IN50;
  input [40:0] IN51;
  input [40:0] IN52;
  input [40:0] IN53;
  input [39:0] IN54;
  input [38:0] IN55;
  input [37:0] IN56;
  input [36:0] IN57;
  input [35:0] IN58;
  input [34:0] IN59;
  input [33:0] IN60;
  input [32:0] IN61;
  input [31:0] IN62;
  input [30:0] IN63;
  input [29:0] IN64;
  input [28:0] IN65;
  input [27:0] IN66;
  input [26:0] IN67;
  input [25:0] IN68;
  input [24:0] IN69;
  input [23:0] IN70;
  input [22:0] IN71;
  input [21:0] IN72;
  input [20:0] IN73;
  input [19:0] IN74;
  input [18:0] IN75;
  input [17:0] IN76;
  input [16:0] IN77;
  input [15:0] IN78;
  input [14:0] IN79;
  input [13:0] IN80;
  input [12:0] IN81;
  input [11:0] IN82;
  input [10:0] IN83;
  input [9:0] IN84;
  input [8:0] IN85;
  input [7:0] IN86;
  input [6:0] IN87;
  input [5:0] IN88;
  input [4:0] IN89;
  input [3:0] IN90;
  input [2:0] IN91;
  input [1:0] IN92;
  input [0:0] IN93;
  output [93:0] Out1;
  output [52:0] Out2;
  wire w2215;
  wire w2216;
  wire w2217;
  wire w2218;
  wire w2219;
  wire w2220;
  wire w2221;
  wire w2222;
  wire w2223;
  wire w2224;
  wire w2225;
  wire w2226;
  wire w2227;
  wire w2228;
  wire w2229;
  wire w2230;
  wire w2231;
  wire w2232;
  wire w2233;
  wire w2234;
  wire w2235;
  wire w2236;
  wire w2237;
  wire w2238;
  wire w2239;
  wire w2240;
  wire w2241;
  wire w2242;
  wire w2243;
  wire w2244;
  wire w2245;
  wire w2246;
  wire w2247;
  wire w2248;
  wire w2249;
  wire w2250;
  wire w2251;
  wire w2252;
  wire w2253;
  wire w2254;
  wire w2255;
  wire w2256;
  wire w2257;
  wire w2258;
  wire w2259;
  wire w2260;
  wire w2261;
  wire w2262;
  wire w2263;
  wire w2264;
  wire w2265;
  wire w2266;
  wire w2267;
  wire w2268;
  wire w2269;
  wire w2270;
  wire w2271;
  wire w2272;
  wire w2273;
  wire w2274;
  wire w2275;
  wire w2276;
  wire w2277;
  wire w2278;
  wire w2279;
  wire w2280;
  wire w2281;
  wire w2282;
  wire w2283;
  wire w2284;
  wire w2285;
  wire w2286;
  wire w2287;
  wire w2288;
  wire w2289;
  wire w2290;
  wire w2291;
  wire w2292;
  wire w2293;
  wire w2295;
  wire w2296;
  wire w2297;
  wire w2298;
  wire w2299;
  wire w2300;
  wire w2301;
  wire w2302;
  wire w2303;
  wire w2304;
  wire w2305;
  wire w2306;
  wire w2307;
  wire w2308;
  wire w2309;
  wire w2310;
  wire w2311;
  wire w2312;
  wire w2313;
  wire w2314;
  wire w2315;
  wire w2316;
  wire w2317;
  wire w2318;
  wire w2319;
  wire w2320;
  wire w2321;
  wire w2322;
  wire w2323;
  wire w2324;
  wire w2325;
  wire w2326;
  wire w2327;
  wire w2328;
  wire w2329;
  wire w2330;
  wire w2331;
  wire w2332;
  wire w2333;
  wire w2334;
  wire w2335;
  wire w2336;
  wire w2337;
  wire w2338;
  wire w2339;
  wire w2340;
  wire w2341;
  wire w2342;
  wire w2343;
  wire w2344;
  wire w2345;
  wire w2346;
  wire w2347;
  wire w2348;
  wire w2349;
  wire w2350;
  wire w2351;
  wire w2352;
  wire w2353;
  wire w2354;
  wire w2355;
  wire w2356;
  wire w2357;
  wire w2358;
  wire w2359;
  wire w2360;
  wire w2361;
  wire w2362;
  wire w2363;
  wire w2364;
  wire w2365;
  wire w2366;
  wire w2367;
  wire w2368;
  wire w2369;
  wire w2370;
  wire w2371;
  wire w2372;
  wire w2373;
  wire w2375;
  wire w2376;
  wire w2377;
  wire w2378;
  wire w2379;
  wire w2380;
  wire w2381;
  wire w2382;
  wire w2383;
  wire w2384;
  wire w2385;
  wire w2386;
  wire w2387;
  wire w2388;
  wire w2389;
  wire w2390;
  wire w2391;
  wire w2392;
  wire w2393;
  wire w2394;
  wire w2395;
  wire w2396;
  wire w2397;
  wire w2398;
  wire w2399;
  wire w2400;
  wire w2401;
  wire w2402;
  wire w2403;
  wire w2404;
  wire w2405;
  wire w2406;
  wire w2407;
  wire w2408;
  wire w2409;
  wire w2410;
  wire w2411;
  wire w2412;
  wire w2413;
  wire w2414;
  wire w2415;
  wire w2416;
  wire w2417;
  wire w2418;
  wire w2419;
  wire w2420;
  wire w2421;
  wire w2422;
  wire w2423;
  wire w2424;
  wire w2425;
  wire w2426;
  wire w2427;
  wire w2428;
  wire w2429;
  wire w2430;
  wire w2431;
  wire w2432;
  wire w2433;
  wire w2434;
  wire w2435;
  wire w2436;
  wire w2437;
  wire w2438;
  wire w2439;
  wire w2440;
  wire w2441;
  wire w2442;
  wire w2443;
  wire w2444;
  wire w2445;
  wire w2446;
  wire w2447;
  wire w2448;
  wire w2449;
  wire w2450;
  wire w2451;
  wire w2452;
  wire w2453;
  wire w2455;
  wire w2456;
  wire w2457;
  wire w2458;
  wire w2459;
  wire w2460;
  wire w2461;
  wire w2462;
  wire w2463;
  wire w2464;
  wire w2465;
  wire w2466;
  wire w2467;
  wire w2468;
  wire w2469;
  wire w2470;
  wire w2471;
  wire w2472;
  wire w2473;
  wire w2474;
  wire w2475;
  wire w2476;
  wire w2477;
  wire w2478;
  wire w2479;
  wire w2480;
  wire w2481;
  wire w2482;
  wire w2483;
  wire w2484;
  wire w2485;
  wire w2486;
  wire w2487;
  wire w2488;
  wire w2489;
  wire w2490;
  wire w2491;
  wire w2492;
  wire w2493;
  wire w2494;
  wire w2495;
  wire w2496;
  wire w2497;
  wire w2498;
  wire w2499;
  wire w2500;
  wire w2501;
  wire w2502;
  wire w2503;
  wire w2504;
  wire w2505;
  wire w2506;
  wire w2507;
  wire w2508;
  wire w2509;
  wire w2510;
  wire w2511;
  wire w2512;
  wire w2513;
  wire w2514;
  wire w2515;
  wire w2516;
  wire w2517;
  wire w2518;
  wire w2519;
  wire w2520;
  wire w2521;
  wire w2522;
  wire w2523;
  wire w2524;
  wire w2525;
  wire w2526;
  wire w2527;
  wire w2528;
  wire w2529;
  wire w2530;
  wire w2531;
  wire w2532;
  wire w2533;
  wire w2535;
  wire w2536;
  wire w2537;
  wire w2538;
  wire w2539;
  wire w2540;
  wire w2541;
  wire w2542;
  wire w2543;
  wire w2544;
  wire w2545;
  wire w2546;
  wire w2547;
  wire w2548;
  wire w2549;
  wire w2550;
  wire w2551;
  wire w2552;
  wire w2553;
  wire w2554;
  wire w2555;
  wire w2556;
  wire w2557;
  wire w2558;
  wire w2559;
  wire w2560;
  wire w2561;
  wire w2562;
  wire w2563;
  wire w2564;
  wire w2565;
  wire w2566;
  wire w2567;
  wire w2568;
  wire w2569;
  wire w2570;
  wire w2571;
  wire w2572;
  wire w2573;
  wire w2574;
  wire w2575;
  wire w2576;
  wire w2577;
  wire w2578;
  wire w2579;
  wire w2580;
  wire w2581;
  wire w2582;
  wire w2583;
  wire w2584;
  wire w2585;
  wire w2586;
  wire w2587;
  wire w2588;
  wire w2589;
  wire w2590;
  wire w2591;
  wire w2592;
  wire w2593;
  wire w2594;
  wire w2595;
  wire w2596;
  wire w2597;
  wire w2598;
  wire w2599;
  wire w2600;
  wire w2601;
  wire w2602;
  wire w2603;
  wire w2604;
  wire w2605;
  wire w2606;
  wire w2607;
  wire w2608;
  wire w2609;
  wire w2610;
  wire w2611;
  wire w2612;
  wire w2613;
  wire w2615;
  wire w2616;
  wire w2617;
  wire w2618;
  wire w2619;
  wire w2620;
  wire w2621;
  wire w2622;
  wire w2623;
  wire w2624;
  wire w2625;
  wire w2626;
  wire w2627;
  wire w2628;
  wire w2629;
  wire w2630;
  wire w2631;
  wire w2632;
  wire w2633;
  wire w2634;
  wire w2635;
  wire w2636;
  wire w2637;
  wire w2638;
  wire w2639;
  wire w2640;
  wire w2641;
  wire w2642;
  wire w2643;
  wire w2644;
  wire w2645;
  wire w2646;
  wire w2647;
  wire w2648;
  wire w2649;
  wire w2650;
  wire w2651;
  wire w2652;
  wire w2653;
  wire w2654;
  wire w2655;
  wire w2656;
  wire w2657;
  wire w2658;
  wire w2659;
  wire w2660;
  wire w2661;
  wire w2662;
  wire w2663;
  wire w2664;
  wire w2665;
  wire w2666;
  wire w2667;
  wire w2668;
  wire w2669;
  wire w2670;
  wire w2671;
  wire w2672;
  wire w2673;
  wire w2674;
  wire w2675;
  wire w2676;
  wire w2677;
  wire w2678;
  wire w2679;
  wire w2680;
  wire w2681;
  wire w2682;
  wire w2683;
  wire w2684;
  wire w2685;
  wire w2686;
  wire w2687;
  wire w2688;
  wire w2689;
  wire w2690;
  wire w2691;
  wire w2692;
  wire w2693;
  wire w2695;
  wire w2696;
  wire w2697;
  wire w2698;
  wire w2699;
  wire w2700;
  wire w2701;
  wire w2702;
  wire w2703;
  wire w2704;
  wire w2705;
  wire w2706;
  wire w2707;
  wire w2708;
  wire w2709;
  wire w2710;
  wire w2711;
  wire w2712;
  wire w2713;
  wire w2714;
  wire w2715;
  wire w2716;
  wire w2717;
  wire w2718;
  wire w2719;
  wire w2720;
  wire w2721;
  wire w2722;
  wire w2723;
  wire w2724;
  wire w2725;
  wire w2726;
  wire w2727;
  wire w2728;
  wire w2729;
  wire w2730;
  wire w2731;
  wire w2732;
  wire w2733;
  wire w2734;
  wire w2735;
  wire w2736;
  wire w2737;
  wire w2738;
  wire w2739;
  wire w2740;
  wire w2741;
  wire w2742;
  wire w2743;
  wire w2744;
  wire w2745;
  wire w2746;
  wire w2747;
  wire w2748;
  wire w2749;
  wire w2750;
  wire w2751;
  wire w2752;
  wire w2753;
  wire w2754;
  wire w2755;
  wire w2756;
  wire w2757;
  wire w2758;
  wire w2759;
  wire w2760;
  wire w2761;
  wire w2762;
  wire w2763;
  wire w2764;
  wire w2765;
  wire w2766;
  wire w2767;
  wire w2768;
  wire w2769;
  wire w2770;
  wire w2771;
  wire w2772;
  wire w2773;
  wire w2775;
  wire w2776;
  wire w2777;
  wire w2778;
  wire w2779;
  wire w2780;
  wire w2781;
  wire w2782;
  wire w2783;
  wire w2784;
  wire w2785;
  wire w2786;
  wire w2787;
  wire w2788;
  wire w2789;
  wire w2790;
  wire w2791;
  wire w2792;
  wire w2793;
  wire w2794;
  wire w2795;
  wire w2796;
  wire w2797;
  wire w2798;
  wire w2799;
  wire w2800;
  wire w2801;
  wire w2802;
  wire w2803;
  wire w2804;
  wire w2805;
  wire w2806;
  wire w2807;
  wire w2808;
  wire w2809;
  wire w2810;
  wire w2811;
  wire w2812;
  wire w2813;
  wire w2814;
  wire w2815;
  wire w2816;
  wire w2817;
  wire w2818;
  wire w2819;
  wire w2820;
  wire w2821;
  wire w2822;
  wire w2823;
  wire w2824;
  wire w2825;
  wire w2826;
  wire w2827;
  wire w2828;
  wire w2829;
  wire w2830;
  wire w2831;
  wire w2832;
  wire w2833;
  wire w2834;
  wire w2835;
  wire w2836;
  wire w2837;
  wire w2838;
  wire w2839;
  wire w2840;
  wire w2841;
  wire w2842;
  wire w2843;
  wire w2844;
  wire w2845;
  wire w2846;
  wire w2847;
  wire w2848;
  wire w2849;
  wire w2850;
  wire w2851;
  wire w2852;
  wire w2853;
  wire w2855;
  wire w2856;
  wire w2857;
  wire w2858;
  wire w2859;
  wire w2860;
  wire w2861;
  wire w2862;
  wire w2863;
  wire w2864;
  wire w2865;
  wire w2866;
  wire w2867;
  wire w2868;
  wire w2869;
  wire w2870;
  wire w2871;
  wire w2872;
  wire w2873;
  wire w2874;
  wire w2875;
  wire w2876;
  wire w2877;
  wire w2878;
  wire w2879;
  wire w2880;
  wire w2881;
  wire w2882;
  wire w2883;
  wire w2884;
  wire w2885;
  wire w2886;
  wire w2887;
  wire w2888;
  wire w2889;
  wire w2890;
  wire w2891;
  wire w2892;
  wire w2893;
  wire w2894;
  wire w2895;
  wire w2896;
  wire w2897;
  wire w2898;
  wire w2899;
  wire w2900;
  wire w2901;
  wire w2902;
  wire w2903;
  wire w2904;
  wire w2905;
  wire w2906;
  wire w2907;
  wire w2908;
  wire w2909;
  wire w2910;
  wire w2911;
  wire w2912;
  wire w2913;
  wire w2914;
  wire w2915;
  wire w2916;
  wire w2917;
  wire w2918;
  wire w2919;
  wire w2920;
  wire w2921;
  wire w2922;
  wire w2923;
  wire w2924;
  wire w2925;
  wire w2926;
  wire w2927;
  wire w2928;
  wire w2929;
  wire w2930;
  wire w2931;
  wire w2932;
  wire w2933;
  wire w2935;
  wire w2936;
  wire w2937;
  wire w2938;
  wire w2939;
  wire w2940;
  wire w2941;
  wire w2942;
  wire w2943;
  wire w2944;
  wire w2945;
  wire w2946;
  wire w2947;
  wire w2948;
  wire w2949;
  wire w2950;
  wire w2951;
  wire w2952;
  wire w2953;
  wire w2954;
  wire w2955;
  wire w2956;
  wire w2957;
  wire w2958;
  wire w2959;
  wire w2960;
  wire w2961;
  wire w2962;
  wire w2963;
  wire w2964;
  wire w2965;
  wire w2966;
  wire w2967;
  wire w2968;
  wire w2969;
  wire w2970;
  wire w2971;
  wire w2972;
  wire w2973;
  wire w2974;
  wire w2975;
  wire w2976;
  wire w2977;
  wire w2978;
  wire w2979;
  wire w2980;
  wire w2981;
  wire w2982;
  wire w2983;
  wire w2984;
  wire w2985;
  wire w2986;
  wire w2987;
  wire w2988;
  wire w2989;
  wire w2990;
  wire w2991;
  wire w2992;
  wire w2993;
  wire w2994;
  wire w2995;
  wire w2996;
  wire w2997;
  wire w2998;
  wire w2999;
  wire w3000;
  wire w3001;
  wire w3002;
  wire w3003;
  wire w3004;
  wire w3005;
  wire w3006;
  wire w3007;
  wire w3008;
  wire w3009;
  wire w3010;
  wire w3011;
  wire w3012;
  wire w3013;
  wire w3015;
  wire w3016;
  wire w3017;
  wire w3018;
  wire w3019;
  wire w3020;
  wire w3021;
  wire w3022;
  wire w3023;
  wire w3024;
  wire w3025;
  wire w3026;
  wire w3027;
  wire w3028;
  wire w3029;
  wire w3030;
  wire w3031;
  wire w3032;
  wire w3033;
  wire w3034;
  wire w3035;
  wire w3036;
  wire w3037;
  wire w3038;
  wire w3039;
  wire w3040;
  wire w3041;
  wire w3042;
  wire w3043;
  wire w3044;
  wire w3045;
  wire w3046;
  wire w3047;
  wire w3048;
  wire w3049;
  wire w3050;
  wire w3051;
  wire w3052;
  wire w3053;
  wire w3054;
  wire w3055;
  wire w3056;
  wire w3057;
  wire w3058;
  wire w3059;
  wire w3060;
  wire w3061;
  wire w3062;
  wire w3063;
  wire w3064;
  wire w3065;
  wire w3066;
  wire w3067;
  wire w3068;
  wire w3069;
  wire w3070;
  wire w3071;
  wire w3072;
  wire w3073;
  wire w3074;
  wire w3075;
  wire w3076;
  wire w3077;
  wire w3078;
  wire w3079;
  wire w3080;
  wire w3081;
  wire w3082;
  wire w3083;
  wire w3084;
  wire w3085;
  wire w3086;
  wire w3087;
  wire w3088;
  wire w3089;
  wire w3090;
  wire w3091;
  wire w3092;
  wire w3093;
  wire w3095;
  wire w3096;
  wire w3097;
  wire w3098;
  wire w3099;
  wire w3100;
  wire w3101;
  wire w3102;
  wire w3103;
  wire w3104;
  wire w3105;
  wire w3106;
  wire w3107;
  wire w3108;
  wire w3109;
  wire w3110;
  wire w3111;
  wire w3112;
  wire w3113;
  wire w3114;
  wire w3115;
  wire w3116;
  wire w3117;
  wire w3118;
  wire w3119;
  wire w3120;
  wire w3121;
  wire w3122;
  wire w3123;
  wire w3124;
  wire w3125;
  wire w3126;
  wire w3127;
  wire w3128;
  wire w3129;
  wire w3130;
  wire w3131;
  wire w3132;
  wire w3133;
  wire w3134;
  wire w3135;
  wire w3136;
  wire w3137;
  wire w3138;
  wire w3139;
  wire w3140;
  wire w3141;
  wire w3142;
  wire w3143;
  wire w3144;
  wire w3145;
  wire w3146;
  wire w3147;
  wire w3148;
  wire w3149;
  wire w3150;
  wire w3151;
  wire w3152;
  wire w3153;
  wire w3154;
  wire w3155;
  wire w3156;
  wire w3157;
  wire w3158;
  wire w3159;
  wire w3160;
  wire w3161;
  wire w3162;
  wire w3163;
  wire w3164;
  wire w3165;
  wire w3166;
  wire w3167;
  wire w3168;
  wire w3169;
  wire w3170;
  wire w3171;
  wire w3172;
  wire w3173;
  wire w3175;
  wire w3176;
  wire w3177;
  wire w3178;
  wire w3179;
  wire w3180;
  wire w3181;
  wire w3182;
  wire w3183;
  wire w3184;
  wire w3185;
  wire w3186;
  wire w3187;
  wire w3188;
  wire w3189;
  wire w3190;
  wire w3191;
  wire w3192;
  wire w3193;
  wire w3194;
  wire w3195;
  wire w3196;
  wire w3197;
  wire w3198;
  wire w3199;
  wire w3200;
  wire w3201;
  wire w3202;
  wire w3203;
  wire w3204;
  wire w3205;
  wire w3206;
  wire w3207;
  wire w3208;
  wire w3209;
  wire w3210;
  wire w3211;
  wire w3212;
  wire w3213;
  wire w3214;
  wire w3215;
  wire w3216;
  wire w3217;
  wire w3218;
  wire w3219;
  wire w3220;
  wire w3221;
  wire w3222;
  wire w3223;
  wire w3224;
  wire w3225;
  wire w3226;
  wire w3227;
  wire w3228;
  wire w3229;
  wire w3230;
  wire w3231;
  wire w3232;
  wire w3233;
  wire w3234;
  wire w3235;
  wire w3236;
  wire w3237;
  wire w3238;
  wire w3239;
  wire w3240;
  wire w3241;
  wire w3242;
  wire w3243;
  wire w3244;
  wire w3245;
  wire w3246;
  wire w3247;
  wire w3248;
  wire w3249;
  wire w3250;
  wire w3251;
  wire w3252;
  wire w3253;
  wire w3255;
  wire w3256;
  wire w3257;
  wire w3258;
  wire w3259;
  wire w3260;
  wire w3261;
  wire w3262;
  wire w3263;
  wire w3264;
  wire w3265;
  wire w3266;
  wire w3267;
  wire w3268;
  wire w3269;
  wire w3270;
  wire w3271;
  wire w3272;
  wire w3273;
  wire w3274;
  wire w3275;
  wire w3276;
  wire w3277;
  wire w3278;
  wire w3279;
  wire w3280;
  wire w3281;
  wire w3282;
  wire w3283;
  wire w3284;
  wire w3285;
  wire w3286;
  wire w3287;
  wire w3288;
  wire w3289;
  wire w3290;
  wire w3291;
  wire w3292;
  wire w3293;
  wire w3294;
  wire w3295;
  wire w3296;
  wire w3297;
  wire w3298;
  wire w3299;
  wire w3300;
  wire w3301;
  wire w3302;
  wire w3303;
  wire w3304;
  wire w3305;
  wire w3306;
  wire w3307;
  wire w3308;
  wire w3309;
  wire w3310;
  wire w3311;
  wire w3312;
  wire w3313;
  wire w3314;
  wire w3315;
  wire w3316;
  wire w3317;
  wire w3318;
  wire w3319;
  wire w3320;
  wire w3321;
  wire w3322;
  wire w3323;
  wire w3324;
  wire w3325;
  wire w3326;
  wire w3327;
  wire w3328;
  wire w3329;
  wire w3330;
  wire w3331;
  wire w3332;
  wire w3333;
  wire w3335;
  wire w3336;
  wire w3337;
  wire w3338;
  wire w3339;
  wire w3340;
  wire w3341;
  wire w3342;
  wire w3343;
  wire w3344;
  wire w3345;
  wire w3346;
  wire w3347;
  wire w3348;
  wire w3349;
  wire w3350;
  wire w3351;
  wire w3352;
  wire w3353;
  wire w3354;
  wire w3355;
  wire w3356;
  wire w3357;
  wire w3358;
  wire w3359;
  wire w3360;
  wire w3361;
  wire w3362;
  wire w3363;
  wire w3364;
  wire w3365;
  wire w3366;
  wire w3367;
  wire w3368;
  wire w3369;
  wire w3370;
  wire w3371;
  wire w3372;
  wire w3373;
  wire w3374;
  wire w3375;
  wire w3376;
  wire w3377;
  wire w3378;
  wire w3379;
  wire w3380;
  wire w3381;
  wire w3382;
  wire w3383;
  wire w3384;
  wire w3385;
  wire w3386;
  wire w3387;
  wire w3388;
  wire w3389;
  wire w3390;
  wire w3391;
  wire w3392;
  wire w3393;
  wire w3394;
  wire w3395;
  wire w3396;
  wire w3397;
  wire w3398;
  wire w3399;
  wire w3400;
  wire w3401;
  wire w3402;
  wire w3403;
  wire w3404;
  wire w3405;
  wire w3406;
  wire w3407;
  wire w3408;
  wire w3409;
  wire w3410;
  wire w3411;
  wire w3412;
  wire w3413;
  wire w3415;
  wire w3416;
  wire w3417;
  wire w3418;
  wire w3419;
  wire w3420;
  wire w3421;
  wire w3422;
  wire w3423;
  wire w3424;
  wire w3425;
  wire w3426;
  wire w3427;
  wire w3428;
  wire w3429;
  wire w3430;
  wire w3431;
  wire w3432;
  wire w3433;
  wire w3434;
  wire w3435;
  wire w3436;
  wire w3437;
  wire w3438;
  wire w3439;
  wire w3440;
  wire w3441;
  wire w3442;
  wire w3443;
  wire w3444;
  wire w3445;
  wire w3446;
  wire w3447;
  wire w3448;
  wire w3449;
  wire w3450;
  wire w3451;
  wire w3452;
  wire w3453;
  wire w3454;
  wire w3455;
  wire w3456;
  wire w3457;
  wire w3458;
  wire w3459;
  wire w3460;
  wire w3461;
  wire w3462;
  wire w3463;
  wire w3464;
  wire w3465;
  wire w3466;
  wire w3467;
  wire w3468;
  wire w3469;
  wire w3470;
  wire w3471;
  wire w3472;
  wire w3473;
  wire w3474;
  wire w3475;
  wire w3476;
  wire w3477;
  wire w3478;
  wire w3479;
  wire w3480;
  wire w3481;
  wire w3482;
  wire w3483;
  wire w3484;
  wire w3485;
  wire w3486;
  wire w3487;
  wire w3488;
  wire w3489;
  wire w3490;
  wire w3491;
  wire w3492;
  wire w3493;
  wire w3495;
  wire w3496;
  wire w3497;
  wire w3498;
  wire w3499;
  wire w3500;
  wire w3501;
  wire w3502;
  wire w3503;
  wire w3504;
  wire w3505;
  wire w3506;
  wire w3507;
  wire w3508;
  wire w3509;
  wire w3510;
  wire w3511;
  wire w3512;
  wire w3513;
  wire w3514;
  wire w3515;
  wire w3516;
  wire w3517;
  wire w3518;
  wire w3519;
  wire w3520;
  wire w3521;
  wire w3522;
  wire w3523;
  wire w3524;
  wire w3525;
  wire w3526;
  wire w3527;
  wire w3528;
  wire w3529;
  wire w3530;
  wire w3531;
  wire w3532;
  wire w3533;
  wire w3534;
  wire w3535;
  wire w3536;
  wire w3537;
  wire w3538;
  wire w3539;
  wire w3540;
  wire w3541;
  wire w3542;
  wire w3543;
  wire w3544;
  wire w3545;
  wire w3546;
  wire w3547;
  wire w3548;
  wire w3549;
  wire w3550;
  wire w3551;
  wire w3552;
  wire w3553;
  wire w3554;
  wire w3555;
  wire w3556;
  wire w3557;
  wire w3558;
  wire w3559;
  wire w3560;
  wire w3561;
  wire w3562;
  wire w3563;
  wire w3564;
  wire w3565;
  wire w3566;
  wire w3567;
  wire w3568;
  wire w3569;
  wire w3570;
  wire w3571;
  wire w3572;
  wire w3573;
  wire w3575;
  wire w3576;
  wire w3577;
  wire w3578;
  wire w3579;
  wire w3580;
  wire w3581;
  wire w3582;
  wire w3583;
  wire w3584;
  wire w3585;
  wire w3586;
  wire w3587;
  wire w3588;
  wire w3589;
  wire w3590;
  wire w3591;
  wire w3592;
  wire w3593;
  wire w3594;
  wire w3595;
  wire w3596;
  wire w3597;
  wire w3598;
  wire w3599;
  wire w3600;
  wire w3601;
  wire w3602;
  wire w3603;
  wire w3604;
  wire w3605;
  wire w3606;
  wire w3607;
  wire w3608;
  wire w3609;
  wire w3610;
  wire w3611;
  wire w3612;
  wire w3613;
  wire w3614;
  wire w3615;
  wire w3616;
  wire w3617;
  wire w3618;
  wire w3619;
  wire w3620;
  wire w3621;
  wire w3622;
  wire w3623;
  wire w3624;
  wire w3625;
  wire w3626;
  wire w3627;
  wire w3628;
  wire w3629;
  wire w3630;
  wire w3631;
  wire w3632;
  wire w3633;
  wire w3634;
  wire w3635;
  wire w3636;
  wire w3637;
  wire w3638;
  wire w3639;
  wire w3640;
  wire w3641;
  wire w3642;
  wire w3643;
  wire w3644;
  wire w3645;
  wire w3646;
  wire w3647;
  wire w3648;
  wire w3649;
  wire w3650;
  wire w3651;
  wire w3652;
  wire w3653;
  wire w3655;
  wire w3656;
  wire w3657;
  wire w3658;
  wire w3659;
  wire w3660;
  wire w3661;
  wire w3662;
  wire w3663;
  wire w3664;
  wire w3665;
  wire w3666;
  wire w3667;
  wire w3668;
  wire w3669;
  wire w3670;
  wire w3671;
  wire w3672;
  wire w3673;
  wire w3674;
  wire w3675;
  wire w3676;
  wire w3677;
  wire w3678;
  wire w3679;
  wire w3680;
  wire w3681;
  wire w3682;
  wire w3683;
  wire w3684;
  wire w3685;
  wire w3686;
  wire w3687;
  wire w3688;
  wire w3689;
  wire w3690;
  wire w3691;
  wire w3692;
  wire w3693;
  wire w3694;
  wire w3695;
  wire w3696;
  wire w3697;
  wire w3698;
  wire w3699;
  wire w3700;
  wire w3701;
  wire w3702;
  wire w3703;
  wire w3704;
  wire w3705;
  wire w3706;
  wire w3707;
  wire w3708;
  wire w3709;
  wire w3710;
  wire w3711;
  wire w3712;
  wire w3713;
  wire w3714;
  wire w3715;
  wire w3716;
  wire w3717;
  wire w3718;
  wire w3719;
  wire w3720;
  wire w3721;
  wire w3722;
  wire w3723;
  wire w3724;
  wire w3725;
  wire w3726;
  wire w3727;
  wire w3728;
  wire w3729;
  wire w3730;
  wire w3731;
  wire w3732;
  wire w3733;
  wire w3735;
  wire w3736;
  wire w3737;
  wire w3738;
  wire w3739;
  wire w3740;
  wire w3741;
  wire w3742;
  wire w3743;
  wire w3744;
  wire w3745;
  wire w3746;
  wire w3747;
  wire w3748;
  wire w3749;
  wire w3750;
  wire w3751;
  wire w3752;
  wire w3753;
  wire w3754;
  wire w3755;
  wire w3756;
  wire w3757;
  wire w3758;
  wire w3759;
  wire w3760;
  wire w3761;
  wire w3762;
  wire w3763;
  wire w3764;
  wire w3765;
  wire w3766;
  wire w3767;
  wire w3768;
  wire w3769;
  wire w3770;
  wire w3771;
  wire w3772;
  wire w3773;
  wire w3774;
  wire w3775;
  wire w3776;
  wire w3777;
  wire w3778;
  wire w3779;
  wire w3780;
  wire w3781;
  wire w3782;
  wire w3783;
  wire w3784;
  wire w3785;
  wire w3786;
  wire w3787;
  wire w3788;
  wire w3789;
  wire w3790;
  wire w3791;
  wire w3792;
  wire w3793;
  wire w3794;
  wire w3795;
  wire w3796;
  wire w3797;
  wire w3798;
  wire w3799;
  wire w3800;
  wire w3801;
  wire w3802;
  wire w3803;
  wire w3804;
  wire w3805;
  wire w3806;
  wire w3807;
  wire w3808;
  wire w3809;
  wire w3810;
  wire w3811;
  wire w3812;
  wire w3813;
  wire w3815;
  wire w3816;
  wire w3817;
  wire w3818;
  wire w3819;
  wire w3820;
  wire w3821;
  wire w3822;
  wire w3823;
  wire w3824;
  wire w3825;
  wire w3826;
  wire w3827;
  wire w3828;
  wire w3829;
  wire w3830;
  wire w3831;
  wire w3832;
  wire w3833;
  wire w3834;
  wire w3835;
  wire w3836;
  wire w3837;
  wire w3838;
  wire w3839;
  wire w3840;
  wire w3841;
  wire w3842;
  wire w3843;
  wire w3844;
  wire w3845;
  wire w3846;
  wire w3847;
  wire w3848;
  wire w3849;
  wire w3850;
  wire w3851;
  wire w3852;
  wire w3853;
  wire w3854;
  wire w3855;
  wire w3856;
  wire w3857;
  wire w3858;
  wire w3859;
  wire w3860;
  wire w3861;
  wire w3862;
  wire w3863;
  wire w3864;
  wire w3865;
  wire w3866;
  wire w3867;
  wire w3868;
  wire w3869;
  wire w3870;
  wire w3871;
  wire w3872;
  wire w3873;
  wire w3874;
  wire w3875;
  wire w3876;
  wire w3877;
  wire w3878;
  wire w3879;
  wire w3880;
  wire w3881;
  wire w3882;
  wire w3883;
  wire w3884;
  wire w3885;
  wire w3886;
  wire w3887;
  wire w3888;
  wire w3889;
  wire w3890;
  wire w3891;
  wire w3892;
  wire w3893;
  wire w3895;
  wire w3896;
  wire w3897;
  wire w3898;
  wire w3899;
  wire w3900;
  wire w3901;
  wire w3902;
  wire w3903;
  wire w3904;
  wire w3905;
  wire w3906;
  wire w3907;
  wire w3908;
  wire w3909;
  wire w3910;
  wire w3911;
  wire w3912;
  wire w3913;
  wire w3914;
  wire w3915;
  wire w3916;
  wire w3917;
  wire w3918;
  wire w3919;
  wire w3920;
  wire w3921;
  wire w3922;
  wire w3923;
  wire w3924;
  wire w3925;
  wire w3926;
  wire w3927;
  wire w3928;
  wire w3929;
  wire w3930;
  wire w3931;
  wire w3932;
  wire w3933;
  wire w3934;
  wire w3935;
  wire w3936;
  wire w3937;
  wire w3938;
  wire w3939;
  wire w3940;
  wire w3941;
  wire w3942;
  wire w3943;
  wire w3944;
  wire w3945;
  wire w3946;
  wire w3947;
  wire w3948;
  wire w3949;
  wire w3950;
  wire w3951;
  wire w3952;
  wire w3953;
  wire w3954;
  wire w3955;
  wire w3956;
  wire w3957;
  wire w3958;
  wire w3959;
  wire w3960;
  wire w3961;
  wire w3962;
  wire w3963;
  wire w3964;
  wire w3965;
  wire w3966;
  wire w3967;
  wire w3968;
  wire w3969;
  wire w3970;
  wire w3971;
  wire w3972;
  wire w3973;
  wire w3975;
  wire w3976;
  wire w3977;
  wire w3978;
  wire w3979;
  wire w3980;
  wire w3981;
  wire w3982;
  wire w3983;
  wire w3984;
  wire w3985;
  wire w3986;
  wire w3987;
  wire w3988;
  wire w3989;
  wire w3990;
  wire w3991;
  wire w3992;
  wire w3993;
  wire w3994;
  wire w3995;
  wire w3996;
  wire w3997;
  wire w3998;
  wire w3999;
  wire w4000;
  wire w4001;
  wire w4002;
  wire w4003;
  wire w4004;
  wire w4005;
  wire w4006;
  wire w4007;
  wire w4008;
  wire w4009;
  wire w4010;
  wire w4011;
  wire w4012;
  wire w4013;
  wire w4014;
  wire w4015;
  wire w4016;
  wire w4017;
  wire w4018;
  wire w4019;
  wire w4020;
  wire w4021;
  wire w4022;
  wire w4023;
  wire w4024;
  wire w4025;
  wire w4026;
  wire w4027;
  wire w4028;
  wire w4029;
  wire w4030;
  wire w4031;
  wire w4032;
  wire w4033;
  wire w4034;
  wire w4035;
  wire w4036;
  wire w4037;
  wire w4038;
  wire w4039;
  wire w4040;
  wire w4041;
  wire w4042;
  wire w4043;
  wire w4044;
  wire w4045;
  wire w4046;
  wire w4047;
  wire w4048;
  wire w4049;
  wire w4050;
  wire w4051;
  wire w4052;
  wire w4053;
  wire w4055;
  wire w4056;
  wire w4057;
  wire w4058;
  wire w4059;
  wire w4060;
  wire w4061;
  wire w4062;
  wire w4063;
  wire w4064;
  wire w4065;
  wire w4066;
  wire w4067;
  wire w4068;
  wire w4069;
  wire w4070;
  wire w4071;
  wire w4072;
  wire w4073;
  wire w4074;
  wire w4075;
  wire w4076;
  wire w4077;
  wire w4078;
  wire w4079;
  wire w4080;
  wire w4081;
  wire w4082;
  wire w4083;
  wire w4084;
  wire w4085;
  wire w4086;
  wire w4087;
  wire w4088;
  wire w4089;
  wire w4090;
  wire w4091;
  wire w4092;
  wire w4093;
  wire w4094;
  wire w4095;
  wire w4096;
  wire w4097;
  wire w4098;
  wire w4099;
  wire w4100;
  wire w4101;
  wire w4102;
  wire w4103;
  wire w4104;
  wire w4105;
  wire w4106;
  wire w4107;
  wire w4108;
  wire w4109;
  wire w4110;
  wire w4111;
  wire w4112;
  wire w4113;
  wire w4114;
  wire w4115;
  wire w4116;
  wire w4117;
  wire w4118;
  wire w4119;
  wire w4120;
  wire w4121;
  wire w4122;
  wire w4123;
  wire w4124;
  wire w4125;
  wire w4126;
  wire w4127;
  wire w4128;
  wire w4129;
  wire w4130;
  wire w4131;
  wire w4132;
  wire w4133;
  wire w4135;
  wire w4136;
  wire w4137;
  wire w4138;
  wire w4139;
  wire w4140;
  wire w4141;
  wire w4142;
  wire w4143;
  wire w4144;
  wire w4145;
  wire w4146;
  wire w4147;
  wire w4148;
  wire w4149;
  wire w4150;
  wire w4151;
  wire w4152;
  wire w4153;
  wire w4154;
  wire w4155;
  wire w4156;
  wire w4157;
  wire w4158;
  wire w4159;
  wire w4160;
  wire w4161;
  wire w4162;
  wire w4163;
  wire w4164;
  wire w4165;
  wire w4166;
  wire w4167;
  wire w4168;
  wire w4169;
  wire w4170;
  wire w4171;
  wire w4172;
  wire w4173;
  wire w4174;
  wire w4175;
  wire w4176;
  wire w4177;
  wire w4178;
  wire w4179;
  wire w4180;
  wire w4181;
  wire w4182;
  wire w4183;
  wire w4184;
  wire w4185;
  wire w4186;
  wire w4187;
  wire w4188;
  wire w4189;
  wire w4190;
  wire w4191;
  wire w4192;
  wire w4193;
  wire w4194;
  wire w4195;
  wire w4196;
  wire w4197;
  wire w4198;
  wire w4199;
  wire w4200;
  wire w4201;
  wire w4202;
  wire w4203;
  wire w4204;
  wire w4205;
  wire w4206;
  wire w4207;
  wire w4208;
  wire w4209;
  wire w4210;
  wire w4211;
  wire w4212;
  wire w4213;
  wire w4215;
  wire w4216;
  wire w4217;
  wire w4218;
  wire w4219;
  wire w4220;
  wire w4221;
  wire w4222;
  wire w4223;
  wire w4224;
  wire w4225;
  wire w4226;
  wire w4227;
  wire w4228;
  wire w4229;
  wire w4230;
  wire w4231;
  wire w4232;
  wire w4233;
  wire w4234;
  wire w4235;
  wire w4236;
  wire w4237;
  wire w4238;
  wire w4239;
  wire w4240;
  wire w4241;
  wire w4242;
  wire w4243;
  wire w4244;
  wire w4245;
  wire w4246;
  wire w4247;
  wire w4248;
  wire w4249;
  wire w4250;
  wire w4251;
  wire w4252;
  wire w4253;
  wire w4254;
  wire w4255;
  wire w4256;
  wire w4257;
  wire w4258;
  wire w4259;
  wire w4260;
  wire w4261;
  wire w4262;
  wire w4263;
  wire w4264;
  wire w4265;
  wire w4266;
  wire w4267;
  wire w4268;
  wire w4269;
  wire w4270;
  wire w4271;
  wire w4272;
  wire w4273;
  wire w4274;
  wire w4275;
  wire w4276;
  wire w4277;
  wire w4278;
  wire w4279;
  wire w4280;
  wire w4281;
  wire w4282;
  wire w4283;
  wire w4284;
  wire w4285;
  wire w4286;
  wire w4287;
  wire w4288;
  wire w4289;
  wire w4290;
  wire w4291;
  wire w4292;
  wire w4293;
  wire w4295;
  wire w4296;
  wire w4297;
  wire w4298;
  wire w4299;
  wire w4300;
  wire w4301;
  wire w4302;
  wire w4303;
  wire w4304;
  wire w4305;
  wire w4306;
  wire w4307;
  wire w4308;
  wire w4309;
  wire w4310;
  wire w4311;
  wire w4312;
  wire w4313;
  wire w4314;
  wire w4315;
  wire w4316;
  wire w4317;
  wire w4318;
  wire w4319;
  wire w4320;
  wire w4321;
  wire w4322;
  wire w4323;
  wire w4324;
  wire w4325;
  wire w4326;
  wire w4327;
  wire w4328;
  wire w4329;
  wire w4330;
  wire w4331;
  wire w4332;
  wire w4333;
  wire w4334;
  wire w4335;
  wire w4336;
  wire w4337;
  wire w4338;
  wire w4339;
  wire w4340;
  wire w4341;
  wire w4342;
  wire w4343;
  wire w4344;
  wire w4345;
  wire w4346;
  wire w4347;
  wire w4348;
  wire w4349;
  wire w4350;
  wire w4351;
  wire w4352;
  wire w4353;
  wire w4354;
  wire w4355;
  wire w4356;
  wire w4357;
  wire w4358;
  wire w4359;
  wire w4360;
  wire w4361;
  wire w4362;
  wire w4363;
  wire w4364;
  wire w4365;
  wire w4366;
  wire w4367;
  wire w4368;
  wire w4369;
  wire w4370;
  wire w4371;
  wire w4372;
  wire w4373;
  wire w4375;
  wire w4376;
  wire w4377;
  wire w4378;
  wire w4379;
  wire w4380;
  wire w4381;
  wire w4382;
  wire w4383;
  wire w4384;
  wire w4385;
  wire w4386;
  wire w4387;
  wire w4388;
  wire w4389;
  wire w4390;
  wire w4391;
  wire w4392;
  wire w4393;
  wire w4394;
  wire w4395;
  wire w4396;
  wire w4397;
  wire w4398;
  wire w4399;
  wire w4400;
  wire w4401;
  wire w4402;
  wire w4403;
  wire w4404;
  wire w4405;
  wire w4406;
  wire w4407;
  wire w4408;
  wire w4409;
  wire w4410;
  wire w4411;
  wire w4412;
  wire w4413;
  wire w4414;
  wire w4415;
  wire w4416;
  wire w4417;
  wire w4418;
  wire w4419;
  wire w4420;
  wire w4421;
  wire w4422;
  wire w4423;
  wire w4424;
  wire w4425;
  wire w4426;
  wire w4427;
  wire w4428;
  wire w4429;
  wire w4430;
  wire w4431;
  wire w4432;
  wire w4433;
  wire w4434;
  wire w4435;
  wire w4436;
  wire w4437;
  wire w4438;
  wire w4439;
  wire w4440;
  wire w4441;
  wire w4442;
  wire w4443;
  wire w4444;
  wire w4445;
  wire w4446;
  wire w4447;
  wire w4448;
  wire w4449;
  wire w4450;
  wire w4451;
  wire w4452;
  wire w4453;
  wire w4455;
  wire w4456;
  wire w4457;
  wire w4458;
  wire w4459;
  wire w4460;
  wire w4461;
  wire w4462;
  wire w4463;
  wire w4464;
  wire w4465;
  wire w4466;
  wire w4467;
  wire w4468;
  wire w4469;
  wire w4470;
  wire w4471;
  wire w4472;
  wire w4473;
  wire w4474;
  wire w4475;
  wire w4476;
  wire w4477;
  wire w4478;
  wire w4479;
  wire w4480;
  wire w4481;
  wire w4482;
  wire w4483;
  wire w4484;
  wire w4485;
  wire w4486;
  wire w4487;
  wire w4488;
  wire w4489;
  wire w4490;
  wire w4491;
  wire w4492;
  wire w4493;
  wire w4494;
  wire w4495;
  wire w4496;
  wire w4497;
  wire w4498;
  wire w4499;
  wire w4500;
  wire w4501;
  wire w4502;
  wire w4503;
  wire w4504;
  wire w4505;
  wire w4506;
  wire w4507;
  wire w4508;
  wire w4509;
  wire w4510;
  wire w4511;
  wire w4512;
  wire w4513;
  wire w4514;
  wire w4515;
  wire w4516;
  wire w4517;
  wire w4518;
  wire w4519;
  wire w4520;
  wire w4521;
  wire w4522;
  wire w4523;
  wire w4524;
  wire w4525;
  wire w4526;
  wire w4527;
  wire w4528;
  wire w4529;
  wire w4530;
  wire w4531;
  wire w4532;
  wire w4533;
  wire w4535;
  wire w4536;
  wire w4537;
  wire w4538;
  wire w4539;
  wire w4540;
  wire w4541;
  wire w4542;
  wire w4543;
  wire w4544;
  wire w4545;
  wire w4546;
  wire w4547;
  wire w4548;
  wire w4549;
  wire w4550;
  wire w4551;
  wire w4552;
  wire w4553;
  wire w4554;
  wire w4555;
  wire w4556;
  wire w4557;
  wire w4558;
  wire w4559;
  wire w4560;
  wire w4561;
  wire w4562;
  wire w4563;
  wire w4564;
  wire w4565;
  wire w4566;
  wire w4567;
  wire w4568;
  wire w4569;
  wire w4570;
  wire w4571;
  wire w4572;
  wire w4573;
  wire w4574;
  wire w4575;
  wire w4576;
  wire w4577;
  wire w4578;
  wire w4579;
  wire w4580;
  wire w4581;
  wire w4582;
  wire w4583;
  wire w4584;
  wire w4585;
  wire w4586;
  wire w4587;
  wire w4588;
  wire w4589;
  wire w4590;
  wire w4591;
  wire w4592;
  wire w4593;
  wire w4594;
  wire w4595;
  wire w4596;
  wire w4597;
  wire w4598;
  wire w4599;
  wire w4600;
  wire w4601;
  wire w4602;
  wire w4603;
  wire w4604;
  wire w4605;
  wire w4606;
  wire w4607;
  wire w4608;
  wire w4609;
  wire w4610;
  wire w4611;
  wire w4612;
  wire w4613;
  wire w4615;
  wire w4616;
  wire w4617;
  wire w4618;
  wire w4619;
  wire w4620;
  wire w4621;
  wire w4622;
  wire w4623;
  wire w4624;
  wire w4625;
  wire w4626;
  wire w4627;
  wire w4628;
  wire w4629;
  wire w4630;
  wire w4631;
  wire w4632;
  wire w4633;
  wire w4634;
  wire w4635;
  wire w4636;
  wire w4637;
  wire w4638;
  wire w4639;
  wire w4640;
  wire w4641;
  wire w4642;
  wire w4643;
  wire w4644;
  wire w4645;
  wire w4646;
  wire w4647;
  wire w4648;
  wire w4649;
  wire w4650;
  wire w4651;
  wire w4652;
  wire w4653;
  wire w4654;
  wire w4655;
  wire w4656;
  wire w4657;
  wire w4658;
  wire w4659;
  wire w4660;
  wire w4661;
  wire w4662;
  wire w4663;
  wire w4664;
  wire w4665;
  wire w4666;
  wire w4667;
  wire w4668;
  wire w4669;
  wire w4670;
  wire w4671;
  wire w4672;
  wire w4673;
  wire w4674;
  wire w4675;
  wire w4676;
  wire w4677;
  wire w4678;
  wire w4679;
  wire w4680;
  wire w4681;
  wire w4682;
  wire w4683;
  wire w4684;
  wire w4685;
  wire w4686;
  wire w4687;
  wire w4688;
  wire w4689;
  wire w4690;
  wire w4691;
  wire w4692;
  wire w4693;
  wire w4695;
  wire w4696;
  wire w4697;
  wire w4698;
  wire w4699;
  wire w4700;
  wire w4701;
  wire w4702;
  wire w4703;
  wire w4704;
  wire w4705;
  wire w4706;
  wire w4707;
  wire w4708;
  wire w4709;
  wire w4710;
  wire w4711;
  wire w4712;
  wire w4713;
  wire w4714;
  wire w4715;
  wire w4716;
  wire w4717;
  wire w4718;
  wire w4719;
  wire w4720;
  wire w4721;
  wire w4722;
  wire w4723;
  wire w4724;
  wire w4725;
  wire w4726;
  wire w4727;
  wire w4728;
  wire w4729;
  wire w4730;
  wire w4731;
  wire w4732;
  wire w4733;
  wire w4734;
  wire w4735;
  wire w4736;
  wire w4737;
  wire w4738;
  wire w4739;
  wire w4740;
  wire w4741;
  wire w4742;
  wire w4743;
  wire w4744;
  wire w4745;
  wire w4746;
  wire w4747;
  wire w4748;
  wire w4749;
  wire w4750;
  wire w4751;
  wire w4752;
  wire w4753;
  wire w4754;
  wire w4755;
  wire w4756;
  wire w4757;
  wire w4758;
  wire w4759;
  wire w4760;
  wire w4761;
  wire w4762;
  wire w4763;
  wire w4764;
  wire w4765;
  wire w4766;
  wire w4767;
  wire w4768;
  wire w4769;
  wire w4770;
  wire w4771;
  wire w4772;
  wire w4773;
  wire w4775;
  wire w4776;
  wire w4777;
  wire w4778;
  wire w4779;
  wire w4780;
  wire w4781;
  wire w4782;
  wire w4783;
  wire w4784;
  wire w4785;
  wire w4786;
  wire w4787;
  wire w4788;
  wire w4789;
  wire w4790;
  wire w4791;
  wire w4792;
  wire w4793;
  wire w4794;
  wire w4795;
  wire w4796;
  wire w4797;
  wire w4798;
  wire w4799;
  wire w4800;
  wire w4801;
  wire w4802;
  wire w4803;
  wire w4804;
  wire w4805;
  wire w4806;
  wire w4807;
  wire w4808;
  wire w4809;
  wire w4810;
  wire w4811;
  wire w4812;
  wire w4813;
  wire w4814;
  wire w4815;
  wire w4816;
  wire w4817;
  wire w4818;
  wire w4819;
  wire w4820;
  wire w4821;
  wire w4822;
  wire w4823;
  wire w4824;
  wire w4825;
  wire w4826;
  wire w4827;
  wire w4828;
  wire w4829;
  wire w4830;
  wire w4831;
  wire w4832;
  wire w4833;
  wire w4834;
  wire w4835;
  wire w4836;
  wire w4837;
  wire w4838;
  wire w4839;
  wire w4840;
  wire w4841;
  wire w4842;
  wire w4843;
  wire w4844;
  wire w4845;
  wire w4846;
  wire w4847;
  wire w4848;
  wire w4849;
  wire w4850;
  wire w4851;
  wire w4852;
  wire w4853;
  wire w4855;
  wire w4856;
  wire w4857;
  wire w4858;
  wire w4859;
  wire w4860;
  wire w4861;
  wire w4862;
  wire w4863;
  wire w4864;
  wire w4865;
  wire w4866;
  wire w4867;
  wire w4868;
  wire w4869;
  wire w4870;
  wire w4871;
  wire w4872;
  wire w4873;
  wire w4874;
  wire w4875;
  wire w4876;
  wire w4877;
  wire w4878;
  wire w4879;
  wire w4880;
  wire w4881;
  wire w4882;
  wire w4883;
  wire w4884;
  wire w4885;
  wire w4886;
  wire w4887;
  wire w4888;
  wire w4889;
  wire w4890;
  wire w4891;
  wire w4892;
  wire w4893;
  wire w4894;
  wire w4895;
  wire w4896;
  wire w4897;
  wire w4898;
  wire w4899;
  wire w4900;
  wire w4901;
  wire w4902;
  wire w4903;
  wire w4904;
  wire w4905;
  wire w4906;
  wire w4907;
  wire w4908;
  wire w4909;
  wire w4910;
  wire w4911;
  wire w4912;
  wire w4913;
  wire w4914;
  wire w4915;
  wire w4916;
  wire w4917;
  wire w4918;
  wire w4919;
  wire w4920;
  wire w4921;
  wire w4922;
  wire w4923;
  wire w4924;
  wire w4925;
  wire w4926;
  wire w4927;
  wire w4928;
  wire w4929;
  wire w4930;
  wire w4931;
  wire w4932;
  wire w4933;
  wire w4935;
  wire w4936;
  wire w4937;
  wire w4938;
  wire w4939;
  wire w4940;
  wire w4941;
  wire w4942;
  wire w4943;
  wire w4944;
  wire w4945;
  wire w4946;
  wire w4947;
  wire w4948;
  wire w4949;
  wire w4950;
  wire w4951;
  wire w4952;
  wire w4953;
  wire w4954;
  wire w4955;
  wire w4956;
  wire w4957;
  wire w4958;
  wire w4959;
  wire w4960;
  wire w4961;
  wire w4962;
  wire w4963;
  wire w4964;
  wire w4965;
  wire w4966;
  wire w4967;
  wire w4968;
  wire w4969;
  wire w4970;
  wire w4971;
  wire w4972;
  wire w4973;
  wire w4974;
  wire w4975;
  wire w4976;
  wire w4977;
  wire w4978;
  wire w4979;
  wire w4980;
  wire w4981;
  wire w4982;
  wire w4983;
  wire w4984;
  wire w4985;
  wire w4986;
  wire w4987;
  wire w4988;
  wire w4989;
  wire w4990;
  wire w4991;
  wire w4992;
  wire w4993;
  wire w4994;
  wire w4995;
  wire w4996;
  wire w4997;
  wire w4998;
  wire w4999;
  wire w5000;
  wire w5001;
  wire w5002;
  wire w5003;
  wire w5004;
  wire w5005;
  wire w5006;
  wire w5007;
  wire w5008;
  wire w5009;
  wire w5010;
  wire w5011;
  wire w5012;
  wire w5013;
  wire w5015;
  wire w5016;
  wire w5017;
  wire w5018;
  wire w5019;
  wire w5020;
  wire w5021;
  wire w5022;
  wire w5023;
  wire w5024;
  wire w5025;
  wire w5026;
  wire w5027;
  wire w5028;
  wire w5029;
  wire w5030;
  wire w5031;
  wire w5032;
  wire w5033;
  wire w5034;
  wire w5035;
  wire w5036;
  wire w5037;
  wire w5038;
  wire w5039;
  wire w5040;
  wire w5041;
  wire w5042;
  wire w5043;
  wire w5044;
  wire w5045;
  wire w5046;
  wire w5047;
  wire w5048;
  wire w5049;
  wire w5050;
  wire w5051;
  wire w5052;
  wire w5053;
  wire w5054;
  wire w5055;
  wire w5056;
  wire w5057;
  wire w5058;
  wire w5059;
  wire w5060;
  wire w5061;
  wire w5062;
  wire w5063;
  wire w5064;
  wire w5065;
  wire w5066;
  wire w5067;
  wire w5068;
  wire w5069;
  wire w5070;
  wire w5071;
  wire w5072;
  wire w5073;
  wire w5074;
  wire w5075;
  wire w5076;
  wire w5077;
  wire w5078;
  wire w5079;
  wire w5080;
  wire w5081;
  wire w5082;
  wire w5083;
  wire w5084;
  wire w5085;
  wire w5086;
  wire w5087;
  wire w5088;
  wire w5089;
  wire w5090;
  wire w5091;
  wire w5092;
  wire w5093;
  wire w5095;
  wire w5096;
  wire w5097;
  wire w5098;
  wire w5099;
  wire w5100;
  wire w5101;
  wire w5102;
  wire w5103;
  wire w5104;
  wire w5105;
  wire w5106;
  wire w5107;
  wire w5108;
  wire w5109;
  wire w5110;
  wire w5111;
  wire w5112;
  wire w5113;
  wire w5114;
  wire w5115;
  wire w5116;
  wire w5117;
  wire w5118;
  wire w5119;
  wire w5120;
  wire w5121;
  wire w5122;
  wire w5123;
  wire w5124;
  wire w5125;
  wire w5126;
  wire w5127;
  wire w5128;
  wire w5129;
  wire w5130;
  wire w5131;
  wire w5132;
  wire w5133;
  wire w5134;
  wire w5135;
  wire w5136;
  wire w5137;
  wire w5138;
  wire w5139;
  wire w5140;
  wire w5141;
  wire w5142;
  wire w5143;
  wire w5144;
  wire w5145;
  wire w5146;
  wire w5147;
  wire w5148;
  wire w5149;
  wire w5150;
  wire w5151;
  wire w5152;
  wire w5153;
  wire w5154;
  wire w5155;
  wire w5156;
  wire w5157;
  wire w5158;
  wire w5159;
  wire w5160;
  wire w5161;
  wire w5162;
  wire w5163;
  wire w5164;
  wire w5165;
  wire w5166;
  wire w5167;
  wire w5168;
  wire w5169;
  wire w5170;
  wire w5171;
  wire w5172;
  wire w5173;
  wire w5175;
  wire w5176;
  wire w5177;
  wire w5178;
  wire w5179;
  wire w5180;
  wire w5181;
  wire w5182;
  wire w5183;
  wire w5184;
  wire w5185;
  wire w5186;
  wire w5187;
  wire w5188;
  wire w5189;
  wire w5190;
  wire w5191;
  wire w5192;
  wire w5193;
  wire w5194;
  wire w5195;
  wire w5196;
  wire w5197;
  wire w5198;
  wire w5199;
  wire w5200;
  wire w5201;
  wire w5202;
  wire w5203;
  wire w5204;
  wire w5205;
  wire w5206;
  wire w5207;
  wire w5208;
  wire w5209;
  wire w5210;
  wire w5211;
  wire w5212;
  wire w5213;
  wire w5214;
  wire w5215;
  wire w5216;
  wire w5217;
  wire w5218;
  wire w5219;
  wire w5220;
  wire w5221;
  wire w5222;
  wire w5223;
  wire w5224;
  wire w5225;
  wire w5226;
  wire w5227;
  wire w5228;
  wire w5229;
  wire w5230;
  wire w5231;
  wire w5232;
  wire w5233;
  wire w5234;
  wire w5235;
  wire w5236;
  wire w5237;
  wire w5238;
  wire w5239;
  wire w5240;
  wire w5241;
  wire w5242;
  wire w5243;
  wire w5244;
  wire w5245;
  wire w5246;
  wire w5247;
  wire w5248;
  wire w5249;
  wire w5250;
  wire w5251;
  wire w5252;
  wire w5253;
  wire w5255;
  wire w5256;
  wire w5257;
  wire w5258;
  wire w5259;
  wire w5260;
  wire w5261;
  wire w5262;
  wire w5263;
  wire w5264;
  wire w5265;
  wire w5266;
  wire w5267;
  wire w5268;
  wire w5269;
  wire w5270;
  wire w5271;
  wire w5272;
  wire w5273;
  wire w5274;
  wire w5275;
  wire w5276;
  wire w5277;
  wire w5278;
  wire w5279;
  wire w5280;
  wire w5281;
  wire w5282;
  wire w5283;
  wire w5284;
  wire w5285;
  wire w5286;
  wire w5287;
  wire w5288;
  wire w5289;
  wire w5290;
  wire w5291;
  wire w5292;
  wire w5293;
  wire w5294;
  wire w5295;
  wire w5296;
  wire w5297;
  wire w5298;
  wire w5299;
  wire w5300;
  wire w5301;
  wire w5302;
  wire w5303;
  wire w5304;
  wire w5305;
  wire w5306;
  wire w5307;
  wire w5308;
  wire w5309;
  wire w5310;
  wire w5311;
  wire w5312;
  wire w5313;
  wire w5314;
  wire w5315;
  wire w5316;
  wire w5317;
  wire w5318;
  wire w5319;
  wire w5320;
  wire w5321;
  wire w5322;
  wire w5323;
  wire w5324;
  wire w5325;
  wire w5326;
  wire w5327;
  wire w5328;
  wire w5329;
  wire w5330;
  wire w5331;
  wire w5332;
  wire w5333;
  wire w5335;
  wire w5336;
  wire w5337;
  wire w5338;
  wire w5339;
  wire w5340;
  wire w5341;
  wire w5342;
  wire w5343;
  wire w5344;
  wire w5345;
  wire w5346;
  wire w5347;
  wire w5348;
  wire w5349;
  wire w5350;
  wire w5351;
  wire w5352;
  wire w5353;
  wire w5354;
  wire w5355;
  wire w5356;
  wire w5357;
  wire w5358;
  wire w5359;
  wire w5360;
  wire w5361;
  wire w5362;
  wire w5363;
  wire w5364;
  wire w5365;
  wire w5366;
  wire w5367;
  wire w5368;
  wire w5369;
  wire w5370;
  wire w5371;
  wire w5372;
  wire w5373;
  wire w5374;
  wire w5375;
  wire w5376;
  wire w5377;
  wire w5378;
  wire w5379;
  wire w5380;
  wire w5381;
  wire w5382;
  wire w5383;
  wire w5384;
  wire w5385;
  wire w5386;
  wire w5387;
  wire w5388;
  wire w5389;
  wire w5390;
  wire w5391;
  wire w5392;
  wire w5393;
  wire w5394;
  wire w5395;
  wire w5396;
  wire w5397;
  wire w5398;
  wire w5399;
  wire w5400;
  wire w5401;
  wire w5402;
  wire w5403;
  wire w5404;
  wire w5405;
  wire w5406;
  wire w5407;
  wire w5408;
  wire w5409;
  wire w5410;
  wire w5411;
  wire w5412;
  wire w5413;
  wire w5415;
  wire w5416;
  wire w5417;
  wire w5418;
  wire w5419;
  wire w5420;
  wire w5421;
  wire w5422;
  wire w5423;
  wire w5424;
  wire w5425;
  wire w5426;
  wire w5427;
  wire w5428;
  wire w5429;
  wire w5430;
  wire w5431;
  wire w5432;
  wire w5433;
  wire w5434;
  wire w5435;
  wire w5436;
  wire w5437;
  wire w5438;
  wire w5439;
  wire w5440;
  wire w5441;
  wire w5442;
  wire w5443;
  wire w5444;
  wire w5445;
  wire w5446;
  wire w5447;
  wire w5448;
  wire w5449;
  wire w5450;
  wire w5451;
  wire w5452;
  wire w5453;
  wire w5454;
  wire w5455;
  wire w5456;
  wire w5457;
  wire w5458;
  wire w5459;
  wire w5460;
  wire w5461;
  wire w5462;
  wire w5463;
  wire w5464;
  wire w5465;
  wire w5466;
  wire w5467;
  wire w5468;
  wire w5469;
  wire w5470;
  wire w5471;
  wire w5472;
  wire w5473;
  wire w5474;
  wire w5475;
  wire w5476;
  wire w5477;
  wire w5478;
  wire w5479;
  wire w5480;
  wire w5481;
  wire w5482;
  wire w5483;
  wire w5484;
  wire w5485;
  wire w5486;
  wire w5487;
  wire w5488;
  wire w5489;
  wire w5490;
  wire w5491;
  wire w5492;
  wire w5493;
  wire w5495;
  wire w5496;
  wire w5497;
  wire w5498;
  wire w5499;
  wire w5500;
  wire w5501;
  wire w5502;
  wire w5503;
  wire w5504;
  wire w5505;
  wire w5506;
  wire w5507;
  wire w5508;
  wire w5509;
  wire w5510;
  wire w5511;
  wire w5512;
  wire w5513;
  wire w5514;
  wire w5515;
  wire w5516;
  wire w5517;
  wire w5518;
  wire w5519;
  wire w5520;
  wire w5521;
  wire w5522;
  wire w5523;
  wire w5524;
  wire w5525;
  wire w5526;
  wire w5527;
  wire w5528;
  wire w5529;
  wire w5530;
  wire w5531;
  wire w5532;
  wire w5533;
  wire w5534;
  wire w5535;
  wire w5536;
  wire w5537;
  wire w5538;
  wire w5539;
  wire w5540;
  wire w5541;
  wire w5542;
  wire w5543;
  wire w5544;
  wire w5545;
  wire w5546;
  wire w5547;
  wire w5548;
  wire w5549;
  wire w5550;
  wire w5551;
  wire w5552;
  wire w5553;
  wire w5554;
  wire w5555;
  wire w5556;
  wire w5557;
  wire w5558;
  wire w5559;
  wire w5560;
  wire w5561;
  wire w5562;
  wire w5563;
  wire w5564;
  wire w5565;
  wire w5566;
  wire w5567;
  wire w5568;
  wire w5569;
  wire w5570;
  wire w5571;
  wire w5572;
  wire w5573;
  wire w5575;
  wire w5576;
  wire w5577;
  wire w5578;
  wire w5579;
  wire w5580;
  wire w5581;
  wire w5582;
  wire w5583;
  wire w5584;
  wire w5585;
  wire w5586;
  wire w5587;
  wire w5588;
  wire w5589;
  wire w5590;
  wire w5591;
  wire w5592;
  wire w5593;
  wire w5594;
  wire w5595;
  wire w5596;
  wire w5597;
  wire w5598;
  wire w5599;
  wire w5600;
  wire w5601;
  wire w5602;
  wire w5603;
  wire w5604;
  wire w5605;
  wire w5606;
  wire w5607;
  wire w5608;
  wire w5609;
  wire w5610;
  wire w5611;
  wire w5612;
  wire w5613;
  wire w5614;
  wire w5615;
  wire w5616;
  wire w5617;
  wire w5618;
  wire w5619;
  wire w5620;
  wire w5621;
  wire w5622;
  wire w5623;
  wire w5624;
  wire w5625;
  wire w5626;
  wire w5627;
  wire w5628;
  wire w5629;
  wire w5630;
  wire w5631;
  wire w5632;
  wire w5633;
  wire w5634;
  wire w5635;
  wire w5636;
  wire w5637;
  wire w5638;
  wire w5639;
  wire w5640;
  wire w5641;
  wire w5642;
  wire w5643;
  wire w5644;
  wire w5645;
  wire w5646;
  wire w5647;
  wire w5648;
  wire w5649;
  wire w5650;
  wire w5651;
  wire w5652;
  wire w5653;
  wire w5655;
  wire w5656;
  wire w5657;
  wire w5658;
  wire w5659;
  wire w5660;
  wire w5661;
  wire w5662;
  wire w5663;
  wire w5664;
  wire w5665;
  wire w5666;
  wire w5667;
  wire w5668;
  wire w5669;
  wire w5670;
  wire w5671;
  wire w5672;
  wire w5673;
  wire w5674;
  wire w5675;
  wire w5676;
  wire w5677;
  wire w5678;
  wire w5679;
  wire w5680;
  wire w5681;
  wire w5682;
  wire w5683;
  wire w5684;
  wire w5685;
  wire w5686;
  wire w5687;
  wire w5688;
  wire w5689;
  wire w5690;
  wire w5691;
  wire w5692;
  wire w5693;
  wire w5694;
  wire w5695;
  wire w5696;
  wire w5697;
  wire w5698;
  wire w5699;
  wire w5700;
  wire w5701;
  wire w5702;
  wire w5703;
  wire w5704;
  wire w5705;
  wire w5706;
  wire w5707;
  wire w5708;
  wire w5709;
  wire w5710;
  wire w5711;
  wire w5712;
  wire w5713;
  wire w5714;
  wire w5715;
  wire w5716;
  wire w5717;
  wire w5718;
  wire w5719;
  wire w5720;
  wire w5721;
  wire w5722;
  wire w5723;
  wire w5724;
  wire w5725;
  wire w5726;
  wire w5727;
  wire w5728;
  wire w5729;
  wire w5730;
  wire w5731;
  wire w5732;
  wire w5733;
  wire w5735;
  wire w5736;
  wire w5737;
  wire w5738;
  wire w5739;
  wire w5740;
  wire w5741;
  wire w5742;
  wire w5743;
  wire w5744;
  wire w5745;
  wire w5746;
  wire w5747;
  wire w5748;
  wire w5749;
  wire w5750;
  wire w5751;
  wire w5752;
  wire w5753;
  wire w5754;
  wire w5755;
  wire w5756;
  wire w5757;
  wire w5758;
  wire w5759;
  wire w5760;
  wire w5761;
  wire w5762;
  wire w5763;
  wire w5764;
  wire w5765;
  wire w5766;
  wire w5767;
  wire w5768;
  wire w5769;
  wire w5770;
  wire w5771;
  wire w5772;
  wire w5773;
  wire w5774;
  wire w5775;
  wire w5776;
  wire w5777;
  wire w5778;
  wire w5779;
  wire w5780;
  wire w5781;
  wire w5782;
  wire w5783;
  wire w5784;
  wire w5785;
  wire w5786;
  wire w5787;
  wire w5788;
  wire w5789;
  wire w5790;
  wire w5791;
  wire w5792;
  wire w5793;
  wire w5794;
  wire w5795;
  wire w5796;
  wire w5797;
  wire w5798;
  wire w5799;
  wire w5800;
  wire w5801;
  wire w5802;
  wire w5803;
  wire w5804;
  wire w5805;
  wire w5806;
  wire w5807;
  wire w5808;
  wire w5809;
  wire w5810;
  wire w5811;
  wire w5812;
  wire w5813;
  wire w5815;
  wire w5816;
  wire w5817;
  wire w5818;
  wire w5819;
  wire w5820;
  wire w5821;
  wire w5822;
  wire w5823;
  wire w5824;
  wire w5825;
  wire w5826;
  wire w5827;
  wire w5828;
  wire w5829;
  wire w5830;
  wire w5831;
  wire w5832;
  wire w5833;
  wire w5834;
  wire w5835;
  wire w5836;
  wire w5837;
  wire w5838;
  wire w5839;
  wire w5840;
  wire w5841;
  wire w5842;
  wire w5843;
  wire w5844;
  wire w5845;
  wire w5846;
  wire w5847;
  wire w5848;
  wire w5849;
  wire w5850;
  wire w5851;
  wire w5852;
  wire w5853;
  wire w5854;
  wire w5855;
  wire w5856;
  wire w5857;
  wire w5858;
  wire w5859;
  wire w5860;
  wire w5861;
  wire w5862;
  wire w5863;
  wire w5864;
  wire w5865;
  wire w5866;
  wire w5867;
  wire w5868;
  wire w5869;
  wire w5870;
  wire w5871;
  wire w5872;
  wire w5873;
  wire w5874;
  wire w5875;
  wire w5876;
  wire w5877;
  wire w5878;
  wire w5879;
  wire w5880;
  wire w5881;
  wire w5882;
  wire w5883;
  wire w5884;
  wire w5885;
  wire w5886;
  wire w5887;
  wire w5888;
  wire w5889;
  wire w5890;
  wire w5891;
  wire w5892;
  wire w5893;
  wire w5895;
  wire w5896;
  wire w5897;
  wire w5898;
  wire w5899;
  wire w5900;
  wire w5901;
  wire w5902;
  wire w5903;
  wire w5904;
  wire w5905;
  wire w5906;
  wire w5907;
  wire w5908;
  wire w5909;
  wire w5910;
  wire w5911;
  wire w5912;
  wire w5913;
  wire w5914;
  wire w5915;
  wire w5916;
  wire w5917;
  wire w5918;
  wire w5919;
  wire w5920;
  wire w5921;
  wire w5922;
  wire w5923;
  wire w5924;
  wire w5925;
  wire w5926;
  wire w5927;
  wire w5928;
  wire w5929;
  wire w5930;
  wire w5931;
  wire w5932;
  wire w5933;
  wire w5934;
  wire w5935;
  wire w5936;
  wire w5937;
  wire w5938;
  wire w5939;
  wire w5940;
  wire w5941;
  wire w5942;
  wire w5943;
  wire w5944;
  wire w5945;
  wire w5946;
  wire w5947;
  wire w5948;
  wire w5949;
  wire w5950;
  wire w5951;
  wire w5952;
  wire w5953;
  wire w5954;
  wire w5955;
  wire w5956;
  wire w5957;
  wire w5958;
  wire w5959;
  wire w5960;
  wire w5961;
  wire w5962;
  wire w5963;
  wire w5964;
  wire w5965;
  wire w5966;
  wire w5967;
  wire w5968;
  wire w5969;
  wire w5970;
  wire w5971;
  wire w5972;
  wire w5973;
  wire w5975;
  wire w5976;
  wire w5977;
  wire w5978;
  wire w5979;
  wire w5980;
  wire w5981;
  wire w5982;
  wire w5983;
  wire w5984;
  wire w5985;
  wire w5986;
  wire w5987;
  wire w5988;
  wire w5989;
  wire w5990;
  wire w5991;
  wire w5992;
  wire w5993;
  wire w5994;
  wire w5995;
  wire w5996;
  wire w5997;
  wire w5998;
  wire w5999;
  wire w6000;
  wire w6001;
  wire w6002;
  wire w6003;
  wire w6004;
  wire w6005;
  wire w6006;
  wire w6007;
  wire w6008;
  wire w6009;
  wire w6010;
  wire w6011;
  wire w6012;
  wire w6013;
  wire w6014;
  wire w6015;
  wire w6016;
  wire w6017;
  wire w6018;
  wire w6019;
  wire w6020;
  wire w6021;
  wire w6022;
  wire w6023;
  wire w6024;
  wire w6025;
  wire w6026;
  wire w6027;
  wire w6028;
  wire w6029;
  wire w6030;
  wire w6031;
  wire w6032;
  wire w6033;
  wire w6034;
  wire w6035;
  wire w6036;
  wire w6037;
  wire w6038;
  wire w6039;
  wire w6040;
  wire w6041;
  wire w6042;
  wire w6043;
  wire w6044;
  wire w6045;
  wire w6046;
  wire w6047;
  wire w6048;
  wire w6049;
  wire w6050;
  wire w6051;
  wire w6052;
  wire w6053;
  wire w6055;
  wire w6056;
  wire w6057;
  wire w6058;
  wire w6059;
  wire w6060;
  wire w6061;
  wire w6062;
  wire w6063;
  wire w6064;
  wire w6065;
  wire w6066;
  wire w6067;
  wire w6068;
  wire w6069;
  wire w6070;
  wire w6071;
  wire w6072;
  wire w6073;
  wire w6074;
  wire w6075;
  wire w6076;
  wire w6077;
  wire w6078;
  wire w6079;
  wire w6080;
  wire w6081;
  wire w6082;
  wire w6083;
  wire w6084;
  wire w6085;
  wire w6086;
  wire w6087;
  wire w6088;
  wire w6089;
  wire w6090;
  wire w6091;
  wire w6092;
  wire w6093;
  wire w6094;
  wire w6095;
  wire w6096;
  wire w6097;
  wire w6098;
  wire w6099;
  wire w6100;
  wire w6101;
  wire w6102;
  wire w6103;
  wire w6104;
  wire w6105;
  wire w6106;
  wire w6107;
  wire w6108;
  wire w6109;
  wire w6110;
  wire w6111;
  wire w6112;
  wire w6113;
  wire w6114;
  wire w6115;
  wire w6116;
  wire w6117;
  wire w6118;
  wire w6119;
  wire w6120;
  wire w6121;
  wire w6122;
  wire w6123;
  wire w6124;
  wire w6125;
  wire w6126;
  wire w6127;
  wire w6128;
  wire w6129;
  wire w6130;
  wire w6131;
  wire w6132;
  wire w6133;
  wire w6135;
  wire w6136;
  wire w6137;
  wire w6138;
  wire w6139;
  wire w6140;
  wire w6141;
  wire w6142;
  wire w6143;
  wire w6144;
  wire w6145;
  wire w6146;
  wire w6147;
  wire w6148;
  wire w6149;
  wire w6150;
  wire w6151;
  wire w6152;
  wire w6153;
  wire w6154;
  wire w6155;
  wire w6156;
  wire w6157;
  wire w6158;
  wire w6159;
  wire w6160;
  wire w6161;
  wire w6162;
  wire w6163;
  wire w6164;
  wire w6165;
  wire w6166;
  wire w6167;
  wire w6168;
  wire w6169;
  wire w6170;
  wire w6171;
  wire w6172;
  wire w6173;
  wire w6174;
  wire w6175;
  wire w6176;
  wire w6177;
  wire w6178;
  wire w6179;
  wire w6180;
  wire w6181;
  wire w6182;
  wire w6183;
  wire w6184;
  wire w6185;
  wire w6186;
  wire w6187;
  wire w6188;
  wire w6189;
  wire w6190;
  wire w6191;
  wire w6192;
  wire w6193;
  wire w6194;
  wire w6195;
  wire w6196;
  wire w6197;
  wire w6198;
  wire w6199;
  wire w6200;
  wire w6201;
  wire w6202;
  wire w6203;
  wire w6204;
  wire w6205;
  wire w6206;
  wire w6207;
  wire w6208;
  wire w6209;
  wire w6210;
  wire w6211;
  wire w6212;
  wire w6213;
  wire w6215;
  wire w6216;
  wire w6217;
  wire w6218;
  wire w6219;
  wire w6220;
  wire w6221;
  wire w6222;
  wire w6223;
  wire w6224;
  wire w6225;
  wire w6226;
  wire w6227;
  wire w6228;
  wire w6229;
  wire w6230;
  wire w6231;
  wire w6232;
  wire w6233;
  wire w6234;
  wire w6235;
  wire w6236;
  wire w6237;
  wire w6238;
  wire w6239;
  wire w6240;
  wire w6241;
  wire w6242;
  wire w6243;
  wire w6244;
  wire w6245;
  wire w6246;
  wire w6247;
  wire w6248;
  wire w6249;
  wire w6250;
  wire w6251;
  wire w6252;
  wire w6253;
  wire w6254;
  wire w6255;
  wire w6256;
  wire w6257;
  wire w6258;
  wire w6259;
  wire w6260;
  wire w6261;
  wire w6262;
  wire w6263;
  wire w6264;
  wire w6265;
  wire w6266;
  wire w6267;
  wire w6268;
  wire w6269;
  wire w6270;
  wire w6271;
  wire w6272;
  wire w6273;
  wire w6274;
  wire w6275;
  wire w6276;
  wire w6277;
  wire w6278;
  wire w6279;
  wire w6280;
  wire w6281;
  wire w6282;
  wire w6283;
  wire w6284;
  wire w6285;
  wire w6286;
  wire w6287;
  wire w6288;
  wire w6289;
  wire w6290;
  wire w6291;
  wire w6292;
  wire w6293;
  wire w6295;
  wire w6296;
  wire w6297;
  wire w6298;
  wire w6299;
  wire w6300;
  wire w6301;
  wire w6302;
  wire w6303;
  wire w6304;
  wire w6305;
  wire w6306;
  wire w6307;
  wire w6308;
  wire w6309;
  wire w6310;
  wire w6311;
  wire w6312;
  wire w6313;
  wire w6314;
  wire w6315;
  wire w6316;
  wire w6317;
  wire w6318;
  wire w6319;
  wire w6320;
  wire w6321;
  wire w6322;
  wire w6323;
  wire w6324;
  wire w6325;
  wire w6326;
  wire w6327;
  wire w6328;
  wire w6329;
  wire w6330;
  wire w6331;
  wire w6332;
  wire w6333;
  wire w6334;
  wire w6335;
  wire w6336;
  wire w6337;
  wire w6338;
  wire w6339;
  wire w6340;
  wire w6341;
  wire w6342;
  wire w6343;
  wire w6344;
  wire w6345;
  wire w6346;
  wire w6347;
  wire w6348;
  wire w6349;
  wire w6350;
  wire w6351;
  wire w6352;
  wire w6353;
  wire w6354;
  wire w6355;
  wire w6356;
  wire w6357;
  wire w6358;
  wire w6359;
  wire w6360;
  wire w6361;
  wire w6362;
  wire w6363;
  wire w6364;
  wire w6365;
  wire w6366;
  wire w6367;
  wire w6368;
  wire w6369;
  wire w6370;
  wire w6371;
  wire w6372;
  wire w6373;
  wire w6375;
  wire w6377;
  wire w6379;
  wire w6381;
  wire w6383;
  wire w6385;
  wire w6387;
  wire w6389;
  wire w6391;
  wire w6393;
  wire w6395;
  wire w6397;
  wire w6399;
  wire w6401;
  wire w6403;
  wire w6405;
  wire w6407;
  wire w6409;
  wire w6411;
  wire w6413;
  wire w6415;
  wire w6417;
  wire w6419;
  wire w6421;
  wire w6423;
  wire w6425;
  wire w6427;
  wire w6429;
  wire w6431;
  wire w6433;
  wire w6435;
  wire w6437;
  wire w6439;
  wire w6441;
  wire w6443;
  wire w6445;
  wire w6447;
  wire w6449;
  wire w6451;
  HalfAdder U0 (IN1[0], IN1[1], Out1[1], w2215);
  FullAdder U1 (w2215, IN2[0], IN2[1], w2216, w2217);
  FullAdder U2 (w2217, IN3[0], IN3[1], w2218, w2219);
  FullAdder U3 (w2219, IN4[0], IN4[1], w2220, w2221);
  FullAdder U4 (w2221, IN5[0], IN5[1], w2222, w2223);
  FullAdder U5 (w2223, IN6[0], IN6[1], w2224, w2225);
  FullAdder U6 (w2225, IN7[0], IN7[1], w2226, w2227);
  FullAdder U7 (w2227, IN8[0], IN8[1], w2228, w2229);
  FullAdder U8 (w2229, IN9[0], IN9[1], w2230, w2231);
  FullAdder U9 (w2231, IN10[0], IN10[1], w2232, w2233);
  FullAdder U10 (w2233, IN11[0], IN11[1], w2234, w2235);
  FullAdder U11 (w2235, IN12[0], IN12[1], w2236, w2237);
  FullAdder U12 (w2237, IN13[0], IN13[1], w2238, w2239);
  FullAdder U13 (w2239, IN14[0], IN14[1], w2240, w2241);
  FullAdder U14 (w2241, IN15[0], IN15[1], w2242, w2243);
  FullAdder U15 (w2243, IN16[0], IN16[1], w2244, w2245);
  FullAdder U16 (w2245, IN17[0], IN17[1], w2246, w2247);
  FullAdder U17 (w2247, IN18[0], IN18[1], w2248, w2249);
  FullAdder U18 (w2249, IN19[0], IN19[1], w2250, w2251);
  FullAdder U19 (w2251, IN20[0], IN20[1], w2252, w2253);
  FullAdder U20 (w2253, IN21[0], IN21[1], w2254, w2255);
  FullAdder U21 (w2255, IN22[0], IN22[1], w2256, w2257);
  FullAdder U22 (w2257, IN23[0], IN23[1], w2258, w2259);
  FullAdder U23 (w2259, IN24[0], IN24[1], w2260, w2261);
  FullAdder U24 (w2261, IN25[0], IN25[1], w2262, w2263);
  FullAdder U25 (w2263, IN26[0], IN26[1], w2264, w2265);
  FullAdder U26 (w2265, IN27[0], IN27[1], w2266, w2267);
  FullAdder U27 (w2267, IN28[0], IN28[1], w2268, w2269);
  FullAdder U28 (w2269, IN29[0], IN29[1], w2270, w2271);
  FullAdder U29 (w2271, IN30[0], IN30[1], w2272, w2273);
  FullAdder U30 (w2273, IN31[0], IN31[1], w2274, w2275);
  FullAdder U31 (w2275, IN32[0], IN32[1], w2276, w2277);
  FullAdder U32 (w2277, IN33[0], IN33[1], w2278, w2279);
  FullAdder U33 (w2279, IN34[0], IN34[1], w2280, w2281);
  FullAdder U34 (w2281, IN35[0], IN35[1], w2282, w2283);
  FullAdder U35 (w2283, IN36[0], IN36[1], w2284, w2285);
  FullAdder U36 (w2285, IN37[0], IN37[1], w2286, w2287);
  FullAdder U37 (w2287, IN38[0], IN38[1], w2288, w2289);
  FullAdder U38 (w2289, IN39[0], IN39[1], w2290, w2291);
  FullAdder U39 (w2291, IN40[0], IN40[1], w2292, w2293);
  HalfAdder U40 (w2216, IN2[2], Out1[2], w2295);
  FullAdder U41 (w2295, w2218, IN3[2], w2296, w2297);
  FullAdder U42 (w2297, w2220, IN4[2], w2298, w2299);
  FullAdder U43 (w2299, w2222, IN5[2], w2300, w2301);
  FullAdder U44 (w2301, w2224, IN6[2], w2302, w2303);
  FullAdder U45 (w2303, w2226, IN7[2], w2304, w2305);
  FullAdder U46 (w2305, w2228, IN8[2], w2306, w2307);
  FullAdder U47 (w2307, w2230, IN9[2], w2308, w2309);
  FullAdder U48 (w2309, w2232, IN10[2], w2310, w2311);
  FullAdder U49 (w2311, w2234, IN11[2], w2312, w2313);
  FullAdder U50 (w2313, w2236, IN12[2], w2314, w2315);
  FullAdder U51 (w2315, w2238, IN13[2], w2316, w2317);
  FullAdder U52 (w2317, w2240, IN14[2], w2318, w2319);
  FullAdder U53 (w2319, w2242, IN15[2], w2320, w2321);
  FullAdder U54 (w2321, w2244, IN16[2], w2322, w2323);
  FullAdder U55 (w2323, w2246, IN17[2], w2324, w2325);
  FullAdder U56 (w2325, w2248, IN18[2], w2326, w2327);
  FullAdder U57 (w2327, w2250, IN19[2], w2328, w2329);
  FullAdder U58 (w2329, w2252, IN20[2], w2330, w2331);
  FullAdder U59 (w2331, w2254, IN21[2], w2332, w2333);
  FullAdder U60 (w2333, w2256, IN22[2], w2334, w2335);
  FullAdder U61 (w2335, w2258, IN23[2], w2336, w2337);
  FullAdder U62 (w2337, w2260, IN24[2], w2338, w2339);
  FullAdder U63 (w2339, w2262, IN25[2], w2340, w2341);
  FullAdder U64 (w2341, w2264, IN26[2], w2342, w2343);
  FullAdder U65 (w2343, w2266, IN27[2], w2344, w2345);
  FullAdder U66 (w2345, w2268, IN28[2], w2346, w2347);
  FullAdder U67 (w2347, w2270, IN29[2], w2348, w2349);
  FullAdder U68 (w2349, w2272, IN30[2], w2350, w2351);
  FullAdder U69 (w2351, w2274, IN31[2], w2352, w2353);
  FullAdder U70 (w2353, w2276, IN32[2], w2354, w2355);
  FullAdder U71 (w2355, w2278, IN33[2], w2356, w2357);
  FullAdder U72 (w2357, w2280, IN34[2], w2358, w2359);
  FullAdder U73 (w2359, w2282, IN35[2], w2360, w2361);
  FullAdder U74 (w2361, w2284, IN36[2], w2362, w2363);
  FullAdder U75 (w2363, w2286, IN37[2], w2364, w2365);
  FullAdder U76 (w2365, w2288, IN38[2], w2366, w2367);
  FullAdder U77 (w2367, w2290, IN39[2], w2368, w2369);
  FullAdder U78 (w2369, w2292, IN40[2], w2370, w2371);
  FullAdder U79 (w2371, w2293, IN41[0], w2372, w2373);
  HalfAdder U80 (w2296, IN3[3], Out1[3], w2375);
  FullAdder U81 (w2375, w2298, IN4[3], w2376, w2377);
  FullAdder U82 (w2377, w2300, IN5[3], w2378, w2379);
  FullAdder U83 (w2379, w2302, IN6[3], w2380, w2381);
  FullAdder U84 (w2381, w2304, IN7[3], w2382, w2383);
  FullAdder U85 (w2383, w2306, IN8[3], w2384, w2385);
  FullAdder U86 (w2385, w2308, IN9[3], w2386, w2387);
  FullAdder U87 (w2387, w2310, IN10[3], w2388, w2389);
  FullAdder U88 (w2389, w2312, IN11[3], w2390, w2391);
  FullAdder U89 (w2391, w2314, IN12[3], w2392, w2393);
  FullAdder U90 (w2393, w2316, IN13[3], w2394, w2395);
  FullAdder U91 (w2395, w2318, IN14[3], w2396, w2397);
  FullAdder U92 (w2397, w2320, IN15[3], w2398, w2399);
  FullAdder U93 (w2399, w2322, IN16[3], w2400, w2401);
  FullAdder U94 (w2401, w2324, IN17[3], w2402, w2403);
  FullAdder U95 (w2403, w2326, IN18[3], w2404, w2405);
  FullAdder U96 (w2405, w2328, IN19[3], w2406, w2407);
  FullAdder U97 (w2407, w2330, IN20[3], w2408, w2409);
  FullAdder U98 (w2409, w2332, IN21[3], w2410, w2411);
  FullAdder U99 (w2411, w2334, IN22[3], w2412, w2413);
  FullAdder U100 (w2413, w2336, IN23[3], w2414, w2415);
  FullAdder U101 (w2415, w2338, IN24[3], w2416, w2417);
  FullAdder U102 (w2417, w2340, IN25[3], w2418, w2419);
  FullAdder U103 (w2419, w2342, IN26[3], w2420, w2421);
  FullAdder U104 (w2421, w2344, IN27[3], w2422, w2423);
  FullAdder U105 (w2423, w2346, IN28[3], w2424, w2425);
  FullAdder U106 (w2425, w2348, IN29[3], w2426, w2427);
  FullAdder U107 (w2427, w2350, IN30[3], w2428, w2429);
  FullAdder U108 (w2429, w2352, IN31[3], w2430, w2431);
  FullAdder U109 (w2431, w2354, IN32[3], w2432, w2433);
  FullAdder U110 (w2433, w2356, IN33[3], w2434, w2435);
  FullAdder U111 (w2435, w2358, IN34[3], w2436, w2437);
  FullAdder U112 (w2437, w2360, IN35[3], w2438, w2439);
  FullAdder U113 (w2439, w2362, IN36[3], w2440, w2441);
  FullAdder U114 (w2441, w2364, IN37[3], w2442, w2443);
  FullAdder U115 (w2443, w2366, IN38[3], w2444, w2445);
  FullAdder U116 (w2445, w2368, IN39[3], w2446, w2447);
  FullAdder U117 (w2447, w2370, IN40[3], w2448, w2449);
  FullAdder U118 (w2449, w2372, IN41[1], w2450, w2451);
  FullAdder U119 (w2451, w2373, IN42[0], w2452, w2453);
  HalfAdder U120 (w2376, IN4[4], Out1[4], w2455);
  FullAdder U121 (w2455, w2378, IN5[4], w2456, w2457);
  FullAdder U122 (w2457, w2380, IN6[4], w2458, w2459);
  FullAdder U123 (w2459, w2382, IN7[4], w2460, w2461);
  FullAdder U124 (w2461, w2384, IN8[4], w2462, w2463);
  FullAdder U125 (w2463, w2386, IN9[4], w2464, w2465);
  FullAdder U126 (w2465, w2388, IN10[4], w2466, w2467);
  FullAdder U127 (w2467, w2390, IN11[4], w2468, w2469);
  FullAdder U128 (w2469, w2392, IN12[4], w2470, w2471);
  FullAdder U129 (w2471, w2394, IN13[4], w2472, w2473);
  FullAdder U130 (w2473, w2396, IN14[4], w2474, w2475);
  FullAdder U131 (w2475, w2398, IN15[4], w2476, w2477);
  FullAdder U132 (w2477, w2400, IN16[4], w2478, w2479);
  FullAdder U133 (w2479, w2402, IN17[4], w2480, w2481);
  FullAdder U134 (w2481, w2404, IN18[4], w2482, w2483);
  FullAdder U135 (w2483, w2406, IN19[4], w2484, w2485);
  FullAdder U136 (w2485, w2408, IN20[4], w2486, w2487);
  FullAdder U137 (w2487, w2410, IN21[4], w2488, w2489);
  FullAdder U138 (w2489, w2412, IN22[4], w2490, w2491);
  FullAdder U139 (w2491, w2414, IN23[4], w2492, w2493);
  FullAdder U140 (w2493, w2416, IN24[4], w2494, w2495);
  FullAdder U141 (w2495, w2418, IN25[4], w2496, w2497);
  FullAdder U142 (w2497, w2420, IN26[4], w2498, w2499);
  FullAdder U143 (w2499, w2422, IN27[4], w2500, w2501);
  FullAdder U144 (w2501, w2424, IN28[4], w2502, w2503);
  FullAdder U145 (w2503, w2426, IN29[4], w2504, w2505);
  FullAdder U146 (w2505, w2428, IN30[4], w2506, w2507);
  FullAdder U147 (w2507, w2430, IN31[4], w2508, w2509);
  FullAdder U148 (w2509, w2432, IN32[4], w2510, w2511);
  FullAdder U149 (w2511, w2434, IN33[4], w2512, w2513);
  FullAdder U150 (w2513, w2436, IN34[4], w2514, w2515);
  FullAdder U151 (w2515, w2438, IN35[4], w2516, w2517);
  FullAdder U152 (w2517, w2440, IN36[4], w2518, w2519);
  FullAdder U153 (w2519, w2442, IN37[4], w2520, w2521);
  FullAdder U154 (w2521, w2444, IN38[4], w2522, w2523);
  FullAdder U155 (w2523, w2446, IN39[4], w2524, w2525);
  FullAdder U156 (w2525, w2448, IN40[4], w2526, w2527);
  FullAdder U157 (w2527, w2450, IN41[2], w2528, w2529);
  FullAdder U158 (w2529, w2452, IN42[1], w2530, w2531);
  FullAdder U159 (w2531, w2453, IN43[0], w2532, w2533);
  HalfAdder U160 (w2456, IN5[5], Out1[5], w2535);
  FullAdder U161 (w2535, w2458, IN6[5], w2536, w2537);
  FullAdder U162 (w2537, w2460, IN7[5], w2538, w2539);
  FullAdder U163 (w2539, w2462, IN8[5], w2540, w2541);
  FullAdder U164 (w2541, w2464, IN9[5], w2542, w2543);
  FullAdder U165 (w2543, w2466, IN10[5], w2544, w2545);
  FullAdder U166 (w2545, w2468, IN11[5], w2546, w2547);
  FullAdder U167 (w2547, w2470, IN12[5], w2548, w2549);
  FullAdder U168 (w2549, w2472, IN13[5], w2550, w2551);
  FullAdder U169 (w2551, w2474, IN14[5], w2552, w2553);
  FullAdder U170 (w2553, w2476, IN15[5], w2554, w2555);
  FullAdder U171 (w2555, w2478, IN16[5], w2556, w2557);
  FullAdder U172 (w2557, w2480, IN17[5], w2558, w2559);
  FullAdder U173 (w2559, w2482, IN18[5], w2560, w2561);
  FullAdder U174 (w2561, w2484, IN19[5], w2562, w2563);
  FullAdder U175 (w2563, w2486, IN20[5], w2564, w2565);
  FullAdder U176 (w2565, w2488, IN21[5], w2566, w2567);
  FullAdder U177 (w2567, w2490, IN22[5], w2568, w2569);
  FullAdder U178 (w2569, w2492, IN23[5], w2570, w2571);
  FullAdder U179 (w2571, w2494, IN24[5], w2572, w2573);
  FullAdder U180 (w2573, w2496, IN25[5], w2574, w2575);
  FullAdder U181 (w2575, w2498, IN26[5], w2576, w2577);
  FullAdder U182 (w2577, w2500, IN27[5], w2578, w2579);
  FullAdder U183 (w2579, w2502, IN28[5], w2580, w2581);
  FullAdder U184 (w2581, w2504, IN29[5], w2582, w2583);
  FullAdder U185 (w2583, w2506, IN30[5], w2584, w2585);
  FullAdder U186 (w2585, w2508, IN31[5], w2586, w2587);
  FullAdder U187 (w2587, w2510, IN32[5], w2588, w2589);
  FullAdder U188 (w2589, w2512, IN33[5], w2590, w2591);
  FullAdder U189 (w2591, w2514, IN34[5], w2592, w2593);
  FullAdder U190 (w2593, w2516, IN35[5], w2594, w2595);
  FullAdder U191 (w2595, w2518, IN36[5], w2596, w2597);
  FullAdder U192 (w2597, w2520, IN37[5], w2598, w2599);
  FullAdder U193 (w2599, w2522, IN38[5], w2600, w2601);
  FullAdder U194 (w2601, w2524, IN39[5], w2602, w2603);
  FullAdder U195 (w2603, w2526, IN40[5], w2604, w2605);
  FullAdder U196 (w2605, w2528, IN41[3], w2606, w2607);
  FullAdder U197 (w2607, w2530, IN42[2], w2608, w2609);
  FullAdder U198 (w2609, w2532, IN43[1], w2610, w2611);
  FullAdder U199 (w2611, w2533, IN44[0], w2612, w2613);
  HalfAdder U200 (w2536, IN6[6], Out1[6], w2615);
  FullAdder U201 (w2615, w2538, IN7[6], w2616, w2617);
  FullAdder U202 (w2617, w2540, IN8[6], w2618, w2619);
  FullAdder U203 (w2619, w2542, IN9[6], w2620, w2621);
  FullAdder U204 (w2621, w2544, IN10[6], w2622, w2623);
  FullAdder U205 (w2623, w2546, IN11[6], w2624, w2625);
  FullAdder U206 (w2625, w2548, IN12[6], w2626, w2627);
  FullAdder U207 (w2627, w2550, IN13[6], w2628, w2629);
  FullAdder U208 (w2629, w2552, IN14[6], w2630, w2631);
  FullAdder U209 (w2631, w2554, IN15[6], w2632, w2633);
  FullAdder U210 (w2633, w2556, IN16[6], w2634, w2635);
  FullAdder U211 (w2635, w2558, IN17[6], w2636, w2637);
  FullAdder U212 (w2637, w2560, IN18[6], w2638, w2639);
  FullAdder U213 (w2639, w2562, IN19[6], w2640, w2641);
  FullAdder U214 (w2641, w2564, IN20[6], w2642, w2643);
  FullAdder U215 (w2643, w2566, IN21[6], w2644, w2645);
  FullAdder U216 (w2645, w2568, IN22[6], w2646, w2647);
  FullAdder U217 (w2647, w2570, IN23[6], w2648, w2649);
  FullAdder U218 (w2649, w2572, IN24[6], w2650, w2651);
  FullAdder U219 (w2651, w2574, IN25[6], w2652, w2653);
  FullAdder U220 (w2653, w2576, IN26[6], w2654, w2655);
  FullAdder U221 (w2655, w2578, IN27[6], w2656, w2657);
  FullAdder U222 (w2657, w2580, IN28[6], w2658, w2659);
  FullAdder U223 (w2659, w2582, IN29[6], w2660, w2661);
  FullAdder U224 (w2661, w2584, IN30[6], w2662, w2663);
  FullAdder U225 (w2663, w2586, IN31[6], w2664, w2665);
  FullAdder U226 (w2665, w2588, IN32[6], w2666, w2667);
  FullAdder U227 (w2667, w2590, IN33[6], w2668, w2669);
  FullAdder U228 (w2669, w2592, IN34[6], w2670, w2671);
  FullAdder U229 (w2671, w2594, IN35[6], w2672, w2673);
  FullAdder U230 (w2673, w2596, IN36[6], w2674, w2675);
  FullAdder U231 (w2675, w2598, IN37[6], w2676, w2677);
  FullAdder U232 (w2677, w2600, IN38[6], w2678, w2679);
  FullAdder U233 (w2679, w2602, IN39[6], w2680, w2681);
  FullAdder U234 (w2681, w2604, IN40[6], w2682, w2683);
  FullAdder U235 (w2683, w2606, IN41[4], w2684, w2685);
  FullAdder U236 (w2685, w2608, IN42[3], w2686, w2687);
  FullAdder U237 (w2687, w2610, IN43[2], w2688, w2689);
  FullAdder U238 (w2689, w2612, IN44[1], w2690, w2691);
  FullAdder U239 (w2691, w2613, IN45[0], w2692, w2693);
  HalfAdder U240 (w2616, IN7[7], Out1[7], w2695);
  FullAdder U241 (w2695, w2618, IN8[7], w2696, w2697);
  FullAdder U242 (w2697, w2620, IN9[7], w2698, w2699);
  FullAdder U243 (w2699, w2622, IN10[7], w2700, w2701);
  FullAdder U244 (w2701, w2624, IN11[7], w2702, w2703);
  FullAdder U245 (w2703, w2626, IN12[7], w2704, w2705);
  FullAdder U246 (w2705, w2628, IN13[7], w2706, w2707);
  FullAdder U247 (w2707, w2630, IN14[7], w2708, w2709);
  FullAdder U248 (w2709, w2632, IN15[7], w2710, w2711);
  FullAdder U249 (w2711, w2634, IN16[7], w2712, w2713);
  FullAdder U250 (w2713, w2636, IN17[7], w2714, w2715);
  FullAdder U251 (w2715, w2638, IN18[7], w2716, w2717);
  FullAdder U252 (w2717, w2640, IN19[7], w2718, w2719);
  FullAdder U253 (w2719, w2642, IN20[7], w2720, w2721);
  FullAdder U254 (w2721, w2644, IN21[7], w2722, w2723);
  FullAdder U255 (w2723, w2646, IN22[7], w2724, w2725);
  FullAdder U256 (w2725, w2648, IN23[7], w2726, w2727);
  FullAdder U257 (w2727, w2650, IN24[7], w2728, w2729);
  FullAdder U258 (w2729, w2652, IN25[7], w2730, w2731);
  FullAdder U259 (w2731, w2654, IN26[7], w2732, w2733);
  FullAdder U260 (w2733, w2656, IN27[7], w2734, w2735);
  FullAdder U261 (w2735, w2658, IN28[7], w2736, w2737);
  FullAdder U262 (w2737, w2660, IN29[7], w2738, w2739);
  FullAdder U263 (w2739, w2662, IN30[7], w2740, w2741);
  FullAdder U264 (w2741, w2664, IN31[7], w2742, w2743);
  FullAdder U265 (w2743, w2666, IN32[7], w2744, w2745);
  FullAdder U266 (w2745, w2668, IN33[7], w2746, w2747);
  FullAdder U267 (w2747, w2670, IN34[7], w2748, w2749);
  FullAdder U268 (w2749, w2672, IN35[7], w2750, w2751);
  FullAdder U269 (w2751, w2674, IN36[7], w2752, w2753);
  FullAdder U270 (w2753, w2676, IN37[7], w2754, w2755);
  FullAdder U271 (w2755, w2678, IN38[7], w2756, w2757);
  FullAdder U272 (w2757, w2680, IN39[7], w2758, w2759);
  FullAdder U273 (w2759, w2682, IN40[7], w2760, w2761);
  FullAdder U274 (w2761, w2684, IN41[5], w2762, w2763);
  FullAdder U275 (w2763, w2686, IN42[4], w2764, w2765);
  FullAdder U276 (w2765, w2688, IN43[3], w2766, w2767);
  FullAdder U277 (w2767, w2690, IN44[2], w2768, w2769);
  FullAdder U278 (w2769, w2692, IN45[1], w2770, w2771);
  FullAdder U279 (w2771, w2693, IN46[0], w2772, w2773);
  HalfAdder U280 (w2696, IN8[8], Out1[8], w2775);
  FullAdder U281 (w2775, w2698, IN9[8], w2776, w2777);
  FullAdder U282 (w2777, w2700, IN10[8], w2778, w2779);
  FullAdder U283 (w2779, w2702, IN11[8], w2780, w2781);
  FullAdder U284 (w2781, w2704, IN12[8], w2782, w2783);
  FullAdder U285 (w2783, w2706, IN13[8], w2784, w2785);
  FullAdder U286 (w2785, w2708, IN14[8], w2786, w2787);
  FullAdder U287 (w2787, w2710, IN15[8], w2788, w2789);
  FullAdder U288 (w2789, w2712, IN16[8], w2790, w2791);
  FullAdder U289 (w2791, w2714, IN17[8], w2792, w2793);
  FullAdder U290 (w2793, w2716, IN18[8], w2794, w2795);
  FullAdder U291 (w2795, w2718, IN19[8], w2796, w2797);
  FullAdder U292 (w2797, w2720, IN20[8], w2798, w2799);
  FullAdder U293 (w2799, w2722, IN21[8], w2800, w2801);
  FullAdder U294 (w2801, w2724, IN22[8], w2802, w2803);
  FullAdder U295 (w2803, w2726, IN23[8], w2804, w2805);
  FullAdder U296 (w2805, w2728, IN24[8], w2806, w2807);
  FullAdder U297 (w2807, w2730, IN25[8], w2808, w2809);
  FullAdder U298 (w2809, w2732, IN26[8], w2810, w2811);
  FullAdder U299 (w2811, w2734, IN27[8], w2812, w2813);
  FullAdder U300 (w2813, w2736, IN28[8], w2814, w2815);
  FullAdder U301 (w2815, w2738, IN29[8], w2816, w2817);
  FullAdder U302 (w2817, w2740, IN30[8], w2818, w2819);
  FullAdder U303 (w2819, w2742, IN31[8], w2820, w2821);
  FullAdder U304 (w2821, w2744, IN32[8], w2822, w2823);
  FullAdder U305 (w2823, w2746, IN33[8], w2824, w2825);
  FullAdder U306 (w2825, w2748, IN34[8], w2826, w2827);
  FullAdder U307 (w2827, w2750, IN35[8], w2828, w2829);
  FullAdder U308 (w2829, w2752, IN36[8], w2830, w2831);
  FullAdder U309 (w2831, w2754, IN37[8], w2832, w2833);
  FullAdder U310 (w2833, w2756, IN38[8], w2834, w2835);
  FullAdder U311 (w2835, w2758, IN39[8], w2836, w2837);
  FullAdder U312 (w2837, w2760, IN40[8], w2838, w2839);
  FullAdder U313 (w2839, w2762, IN41[6], w2840, w2841);
  FullAdder U314 (w2841, w2764, IN42[5], w2842, w2843);
  FullAdder U315 (w2843, w2766, IN43[4], w2844, w2845);
  FullAdder U316 (w2845, w2768, IN44[3], w2846, w2847);
  FullAdder U317 (w2847, w2770, IN45[2], w2848, w2849);
  FullAdder U318 (w2849, w2772, IN46[1], w2850, w2851);
  FullAdder U319 (w2851, w2773, IN47[0], w2852, w2853);
  HalfAdder U320 (w2776, IN9[9], Out1[9], w2855);
  FullAdder U321 (w2855, w2778, IN10[9], w2856, w2857);
  FullAdder U322 (w2857, w2780, IN11[9], w2858, w2859);
  FullAdder U323 (w2859, w2782, IN12[9], w2860, w2861);
  FullAdder U324 (w2861, w2784, IN13[9], w2862, w2863);
  FullAdder U325 (w2863, w2786, IN14[9], w2864, w2865);
  FullAdder U326 (w2865, w2788, IN15[9], w2866, w2867);
  FullAdder U327 (w2867, w2790, IN16[9], w2868, w2869);
  FullAdder U328 (w2869, w2792, IN17[9], w2870, w2871);
  FullAdder U329 (w2871, w2794, IN18[9], w2872, w2873);
  FullAdder U330 (w2873, w2796, IN19[9], w2874, w2875);
  FullAdder U331 (w2875, w2798, IN20[9], w2876, w2877);
  FullAdder U332 (w2877, w2800, IN21[9], w2878, w2879);
  FullAdder U333 (w2879, w2802, IN22[9], w2880, w2881);
  FullAdder U334 (w2881, w2804, IN23[9], w2882, w2883);
  FullAdder U335 (w2883, w2806, IN24[9], w2884, w2885);
  FullAdder U336 (w2885, w2808, IN25[9], w2886, w2887);
  FullAdder U337 (w2887, w2810, IN26[9], w2888, w2889);
  FullAdder U338 (w2889, w2812, IN27[9], w2890, w2891);
  FullAdder U339 (w2891, w2814, IN28[9], w2892, w2893);
  FullAdder U340 (w2893, w2816, IN29[9], w2894, w2895);
  FullAdder U341 (w2895, w2818, IN30[9], w2896, w2897);
  FullAdder U342 (w2897, w2820, IN31[9], w2898, w2899);
  FullAdder U343 (w2899, w2822, IN32[9], w2900, w2901);
  FullAdder U344 (w2901, w2824, IN33[9], w2902, w2903);
  FullAdder U345 (w2903, w2826, IN34[9], w2904, w2905);
  FullAdder U346 (w2905, w2828, IN35[9], w2906, w2907);
  FullAdder U347 (w2907, w2830, IN36[9], w2908, w2909);
  FullAdder U348 (w2909, w2832, IN37[9], w2910, w2911);
  FullAdder U349 (w2911, w2834, IN38[9], w2912, w2913);
  FullAdder U350 (w2913, w2836, IN39[9], w2914, w2915);
  FullAdder U351 (w2915, w2838, IN40[9], w2916, w2917);
  FullAdder U352 (w2917, w2840, IN41[7], w2918, w2919);
  FullAdder U353 (w2919, w2842, IN42[6], w2920, w2921);
  FullAdder U354 (w2921, w2844, IN43[5], w2922, w2923);
  FullAdder U355 (w2923, w2846, IN44[4], w2924, w2925);
  FullAdder U356 (w2925, w2848, IN45[3], w2926, w2927);
  FullAdder U357 (w2927, w2850, IN46[2], w2928, w2929);
  FullAdder U358 (w2929, w2852, IN47[1], w2930, w2931);
  FullAdder U359 (w2931, w2853, IN48[0], w2932, w2933);
  HalfAdder U360 (w2856, IN10[10], Out1[10], w2935);
  FullAdder U361 (w2935, w2858, IN11[10], w2936, w2937);
  FullAdder U362 (w2937, w2860, IN12[10], w2938, w2939);
  FullAdder U363 (w2939, w2862, IN13[10], w2940, w2941);
  FullAdder U364 (w2941, w2864, IN14[10], w2942, w2943);
  FullAdder U365 (w2943, w2866, IN15[10], w2944, w2945);
  FullAdder U366 (w2945, w2868, IN16[10], w2946, w2947);
  FullAdder U367 (w2947, w2870, IN17[10], w2948, w2949);
  FullAdder U368 (w2949, w2872, IN18[10], w2950, w2951);
  FullAdder U369 (w2951, w2874, IN19[10], w2952, w2953);
  FullAdder U370 (w2953, w2876, IN20[10], w2954, w2955);
  FullAdder U371 (w2955, w2878, IN21[10], w2956, w2957);
  FullAdder U372 (w2957, w2880, IN22[10], w2958, w2959);
  FullAdder U373 (w2959, w2882, IN23[10], w2960, w2961);
  FullAdder U374 (w2961, w2884, IN24[10], w2962, w2963);
  FullAdder U375 (w2963, w2886, IN25[10], w2964, w2965);
  FullAdder U376 (w2965, w2888, IN26[10], w2966, w2967);
  FullAdder U377 (w2967, w2890, IN27[10], w2968, w2969);
  FullAdder U378 (w2969, w2892, IN28[10], w2970, w2971);
  FullAdder U379 (w2971, w2894, IN29[10], w2972, w2973);
  FullAdder U380 (w2973, w2896, IN30[10], w2974, w2975);
  FullAdder U381 (w2975, w2898, IN31[10], w2976, w2977);
  FullAdder U382 (w2977, w2900, IN32[10], w2978, w2979);
  FullAdder U383 (w2979, w2902, IN33[10], w2980, w2981);
  FullAdder U384 (w2981, w2904, IN34[10], w2982, w2983);
  FullAdder U385 (w2983, w2906, IN35[10], w2984, w2985);
  FullAdder U386 (w2985, w2908, IN36[10], w2986, w2987);
  FullAdder U387 (w2987, w2910, IN37[10], w2988, w2989);
  FullAdder U388 (w2989, w2912, IN38[10], w2990, w2991);
  FullAdder U389 (w2991, w2914, IN39[10], w2992, w2993);
  FullAdder U390 (w2993, w2916, IN40[10], w2994, w2995);
  FullAdder U391 (w2995, w2918, IN41[8], w2996, w2997);
  FullAdder U392 (w2997, w2920, IN42[7], w2998, w2999);
  FullAdder U393 (w2999, w2922, IN43[6], w3000, w3001);
  FullAdder U394 (w3001, w2924, IN44[5], w3002, w3003);
  FullAdder U395 (w3003, w2926, IN45[4], w3004, w3005);
  FullAdder U396 (w3005, w2928, IN46[3], w3006, w3007);
  FullAdder U397 (w3007, w2930, IN47[2], w3008, w3009);
  FullAdder U398 (w3009, w2932, IN48[1], w3010, w3011);
  FullAdder U399 (w3011, w2933, IN49[0], w3012, w3013);
  HalfAdder U400 (w2936, IN11[11], Out1[11], w3015);
  FullAdder U401 (w3015, w2938, IN12[11], w3016, w3017);
  FullAdder U402 (w3017, w2940, IN13[11], w3018, w3019);
  FullAdder U403 (w3019, w2942, IN14[11], w3020, w3021);
  FullAdder U404 (w3021, w2944, IN15[11], w3022, w3023);
  FullAdder U405 (w3023, w2946, IN16[11], w3024, w3025);
  FullAdder U406 (w3025, w2948, IN17[11], w3026, w3027);
  FullAdder U407 (w3027, w2950, IN18[11], w3028, w3029);
  FullAdder U408 (w3029, w2952, IN19[11], w3030, w3031);
  FullAdder U409 (w3031, w2954, IN20[11], w3032, w3033);
  FullAdder U410 (w3033, w2956, IN21[11], w3034, w3035);
  FullAdder U411 (w3035, w2958, IN22[11], w3036, w3037);
  FullAdder U412 (w3037, w2960, IN23[11], w3038, w3039);
  FullAdder U413 (w3039, w2962, IN24[11], w3040, w3041);
  FullAdder U414 (w3041, w2964, IN25[11], w3042, w3043);
  FullAdder U415 (w3043, w2966, IN26[11], w3044, w3045);
  FullAdder U416 (w3045, w2968, IN27[11], w3046, w3047);
  FullAdder U417 (w3047, w2970, IN28[11], w3048, w3049);
  FullAdder U418 (w3049, w2972, IN29[11], w3050, w3051);
  FullAdder U419 (w3051, w2974, IN30[11], w3052, w3053);
  FullAdder U420 (w3053, w2976, IN31[11], w3054, w3055);
  FullAdder U421 (w3055, w2978, IN32[11], w3056, w3057);
  FullAdder U422 (w3057, w2980, IN33[11], w3058, w3059);
  FullAdder U423 (w3059, w2982, IN34[11], w3060, w3061);
  FullAdder U424 (w3061, w2984, IN35[11], w3062, w3063);
  FullAdder U425 (w3063, w2986, IN36[11], w3064, w3065);
  FullAdder U426 (w3065, w2988, IN37[11], w3066, w3067);
  FullAdder U427 (w3067, w2990, IN38[11], w3068, w3069);
  FullAdder U428 (w3069, w2992, IN39[11], w3070, w3071);
  FullAdder U429 (w3071, w2994, IN40[11], w3072, w3073);
  FullAdder U430 (w3073, w2996, IN41[9], w3074, w3075);
  FullAdder U431 (w3075, w2998, IN42[8], w3076, w3077);
  FullAdder U432 (w3077, w3000, IN43[7], w3078, w3079);
  FullAdder U433 (w3079, w3002, IN44[6], w3080, w3081);
  FullAdder U434 (w3081, w3004, IN45[5], w3082, w3083);
  FullAdder U435 (w3083, w3006, IN46[4], w3084, w3085);
  FullAdder U436 (w3085, w3008, IN47[3], w3086, w3087);
  FullAdder U437 (w3087, w3010, IN48[2], w3088, w3089);
  FullAdder U438 (w3089, w3012, IN49[1], w3090, w3091);
  FullAdder U439 (w3091, w3013, IN50[0], w3092, w3093);
  HalfAdder U440 (w3016, IN12[12], Out1[12], w3095);
  FullAdder U441 (w3095, w3018, IN13[12], w3096, w3097);
  FullAdder U442 (w3097, w3020, IN14[12], w3098, w3099);
  FullAdder U443 (w3099, w3022, IN15[12], w3100, w3101);
  FullAdder U444 (w3101, w3024, IN16[12], w3102, w3103);
  FullAdder U445 (w3103, w3026, IN17[12], w3104, w3105);
  FullAdder U446 (w3105, w3028, IN18[12], w3106, w3107);
  FullAdder U447 (w3107, w3030, IN19[12], w3108, w3109);
  FullAdder U448 (w3109, w3032, IN20[12], w3110, w3111);
  FullAdder U449 (w3111, w3034, IN21[12], w3112, w3113);
  FullAdder U450 (w3113, w3036, IN22[12], w3114, w3115);
  FullAdder U451 (w3115, w3038, IN23[12], w3116, w3117);
  FullAdder U452 (w3117, w3040, IN24[12], w3118, w3119);
  FullAdder U453 (w3119, w3042, IN25[12], w3120, w3121);
  FullAdder U454 (w3121, w3044, IN26[12], w3122, w3123);
  FullAdder U455 (w3123, w3046, IN27[12], w3124, w3125);
  FullAdder U456 (w3125, w3048, IN28[12], w3126, w3127);
  FullAdder U457 (w3127, w3050, IN29[12], w3128, w3129);
  FullAdder U458 (w3129, w3052, IN30[12], w3130, w3131);
  FullAdder U459 (w3131, w3054, IN31[12], w3132, w3133);
  FullAdder U460 (w3133, w3056, IN32[12], w3134, w3135);
  FullAdder U461 (w3135, w3058, IN33[12], w3136, w3137);
  FullAdder U462 (w3137, w3060, IN34[12], w3138, w3139);
  FullAdder U463 (w3139, w3062, IN35[12], w3140, w3141);
  FullAdder U464 (w3141, w3064, IN36[12], w3142, w3143);
  FullAdder U465 (w3143, w3066, IN37[12], w3144, w3145);
  FullAdder U466 (w3145, w3068, IN38[12], w3146, w3147);
  FullAdder U467 (w3147, w3070, IN39[12], w3148, w3149);
  FullAdder U468 (w3149, w3072, IN40[12], w3150, w3151);
  FullAdder U469 (w3151, w3074, IN41[10], w3152, w3153);
  FullAdder U470 (w3153, w3076, IN42[9], w3154, w3155);
  FullAdder U471 (w3155, w3078, IN43[8], w3156, w3157);
  FullAdder U472 (w3157, w3080, IN44[7], w3158, w3159);
  FullAdder U473 (w3159, w3082, IN45[6], w3160, w3161);
  FullAdder U474 (w3161, w3084, IN46[5], w3162, w3163);
  FullAdder U475 (w3163, w3086, IN47[4], w3164, w3165);
  FullAdder U476 (w3165, w3088, IN48[3], w3166, w3167);
  FullAdder U477 (w3167, w3090, IN49[2], w3168, w3169);
  FullAdder U478 (w3169, w3092, IN50[1], w3170, w3171);
  FullAdder U479 (w3171, w3093, IN51[0], w3172, w3173);
  HalfAdder U480 (w3096, IN13[13], Out1[13], w3175);
  FullAdder U481 (w3175, w3098, IN14[13], w3176, w3177);
  FullAdder U482 (w3177, w3100, IN15[13], w3178, w3179);
  FullAdder U483 (w3179, w3102, IN16[13], w3180, w3181);
  FullAdder U484 (w3181, w3104, IN17[13], w3182, w3183);
  FullAdder U485 (w3183, w3106, IN18[13], w3184, w3185);
  FullAdder U486 (w3185, w3108, IN19[13], w3186, w3187);
  FullAdder U487 (w3187, w3110, IN20[13], w3188, w3189);
  FullAdder U488 (w3189, w3112, IN21[13], w3190, w3191);
  FullAdder U489 (w3191, w3114, IN22[13], w3192, w3193);
  FullAdder U490 (w3193, w3116, IN23[13], w3194, w3195);
  FullAdder U491 (w3195, w3118, IN24[13], w3196, w3197);
  FullAdder U492 (w3197, w3120, IN25[13], w3198, w3199);
  FullAdder U493 (w3199, w3122, IN26[13], w3200, w3201);
  FullAdder U494 (w3201, w3124, IN27[13], w3202, w3203);
  FullAdder U495 (w3203, w3126, IN28[13], w3204, w3205);
  FullAdder U496 (w3205, w3128, IN29[13], w3206, w3207);
  FullAdder U497 (w3207, w3130, IN30[13], w3208, w3209);
  FullAdder U498 (w3209, w3132, IN31[13], w3210, w3211);
  FullAdder U499 (w3211, w3134, IN32[13], w3212, w3213);
  FullAdder U500 (w3213, w3136, IN33[13], w3214, w3215);
  FullAdder U501 (w3215, w3138, IN34[13], w3216, w3217);
  FullAdder U502 (w3217, w3140, IN35[13], w3218, w3219);
  FullAdder U503 (w3219, w3142, IN36[13], w3220, w3221);
  FullAdder U504 (w3221, w3144, IN37[13], w3222, w3223);
  FullAdder U505 (w3223, w3146, IN38[13], w3224, w3225);
  FullAdder U506 (w3225, w3148, IN39[13], w3226, w3227);
  FullAdder U507 (w3227, w3150, IN40[13], w3228, w3229);
  FullAdder U508 (w3229, w3152, IN41[11], w3230, w3231);
  FullAdder U509 (w3231, w3154, IN42[10], w3232, w3233);
  FullAdder U510 (w3233, w3156, IN43[9], w3234, w3235);
  FullAdder U511 (w3235, w3158, IN44[8], w3236, w3237);
  FullAdder U512 (w3237, w3160, IN45[7], w3238, w3239);
  FullAdder U513 (w3239, w3162, IN46[6], w3240, w3241);
  FullAdder U514 (w3241, w3164, IN47[5], w3242, w3243);
  FullAdder U515 (w3243, w3166, IN48[4], w3244, w3245);
  FullAdder U516 (w3245, w3168, IN49[3], w3246, w3247);
  FullAdder U517 (w3247, w3170, IN50[2], w3248, w3249);
  FullAdder U518 (w3249, w3172, IN51[1], w3250, w3251);
  FullAdder U519 (w3251, w3173, IN52[0], w3252, w3253);
  HalfAdder U520 (w3176, IN14[14], Out1[14], w3255);
  FullAdder U521 (w3255, w3178, IN15[14], w3256, w3257);
  FullAdder U522 (w3257, w3180, IN16[14], w3258, w3259);
  FullAdder U523 (w3259, w3182, IN17[14], w3260, w3261);
  FullAdder U524 (w3261, w3184, IN18[14], w3262, w3263);
  FullAdder U525 (w3263, w3186, IN19[14], w3264, w3265);
  FullAdder U526 (w3265, w3188, IN20[14], w3266, w3267);
  FullAdder U527 (w3267, w3190, IN21[14], w3268, w3269);
  FullAdder U528 (w3269, w3192, IN22[14], w3270, w3271);
  FullAdder U529 (w3271, w3194, IN23[14], w3272, w3273);
  FullAdder U530 (w3273, w3196, IN24[14], w3274, w3275);
  FullAdder U531 (w3275, w3198, IN25[14], w3276, w3277);
  FullAdder U532 (w3277, w3200, IN26[14], w3278, w3279);
  FullAdder U533 (w3279, w3202, IN27[14], w3280, w3281);
  FullAdder U534 (w3281, w3204, IN28[14], w3282, w3283);
  FullAdder U535 (w3283, w3206, IN29[14], w3284, w3285);
  FullAdder U536 (w3285, w3208, IN30[14], w3286, w3287);
  FullAdder U537 (w3287, w3210, IN31[14], w3288, w3289);
  FullAdder U538 (w3289, w3212, IN32[14], w3290, w3291);
  FullAdder U539 (w3291, w3214, IN33[14], w3292, w3293);
  FullAdder U540 (w3293, w3216, IN34[14], w3294, w3295);
  FullAdder U541 (w3295, w3218, IN35[14], w3296, w3297);
  FullAdder U542 (w3297, w3220, IN36[14], w3298, w3299);
  FullAdder U543 (w3299, w3222, IN37[14], w3300, w3301);
  FullAdder U544 (w3301, w3224, IN38[14], w3302, w3303);
  FullAdder U545 (w3303, w3226, IN39[14], w3304, w3305);
  FullAdder U546 (w3305, w3228, IN40[14], w3306, w3307);
  FullAdder U547 (w3307, w3230, IN41[12], w3308, w3309);
  FullAdder U548 (w3309, w3232, IN42[11], w3310, w3311);
  FullAdder U549 (w3311, w3234, IN43[10], w3312, w3313);
  FullAdder U550 (w3313, w3236, IN44[9], w3314, w3315);
  FullAdder U551 (w3315, w3238, IN45[8], w3316, w3317);
  FullAdder U552 (w3317, w3240, IN46[7], w3318, w3319);
  FullAdder U553 (w3319, w3242, IN47[6], w3320, w3321);
  FullAdder U554 (w3321, w3244, IN48[5], w3322, w3323);
  FullAdder U555 (w3323, w3246, IN49[4], w3324, w3325);
  FullAdder U556 (w3325, w3248, IN50[3], w3326, w3327);
  FullAdder U557 (w3327, w3250, IN51[2], w3328, w3329);
  FullAdder U558 (w3329, w3252, IN52[1], w3330, w3331);
  FullAdder U559 (w3331, w3253, IN53[0], w3332, w3333);
  HalfAdder U560 (w3256, IN15[15], Out1[15], w3335);
  FullAdder U561 (w3335, w3258, IN16[15], w3336, w3337);
  FullAdder U562 (w3337, w3260, IN17[15], w3338, w3339);
  FullAdder U563 (w3339, w3262, IN18[15], w3340, w3341);
  FullAdder U564 (w3341, w3264, IN19[15], w3342, w3343);
  FullAdder U565 (w3343, w3266, IN20[15], w3344, w3345);
  FullAdder U566 (w3345, w3268, IN21[15], w3346, w3347);
  FullAdder U567 (w3347, w3270, IN22[15], w3348, w3349);
  FullAdder U568 (w3349, w3272, IN23[15], w3350, w3351);
  FullAdder U569 (w3351, w3274, IN24[15], w3352, w3353);
  FullAdder U570 (w3353, w3276, IN25[15], w3354, w3355);
  FullAdder U571 (w3355, w3278, IN26[15], w3356, w3357);
  FullAdder U572 (w3357, w3280, IN27[15], w3358, w3359);
  FullAdder U573 (w3359, w3282, IN28[15], w3360, w3361);
  FullAdder U574 (w3361, w3284, IN29[15], w3362, w3363);
  FullAdder U575 (w3363, w3286, IN30[15], w3364, w3365);
  FullAdder U576 (w3365, w3288, IN31[15], w3366, w3367);
  FullAdder U577 (w3367, w3290, IN32[15], w3368, w3369);
  FullAdder U578 (w3369, w3292, IN33[15], w3370, w3371);
  FullAdder U579 (w3371, w3294, IN34[15], w3372, w3373);
  FullAdder U580 (w3373, w3296, IN35[15], w3374, w3375);
  FullAdder U581 (w3375, w3298, IN36[15], w3376, w3377);
  FullAdder U582 (w3377, w3300, IN37[15], w3378, w3379);
  FullAdder U583 (w3379, w3302, IN38[15], w3380, w3381);
  FullAdder U584 (w3381, w3304, IN39[15], w3382, w3383);
  FullAdder U585 (w3383, w3306, IN40[15], w3384, w3385);
  FullAdder U586 (w3385, w3308, IN41[13], w3386, w3387);
  FullAdder U587 (w3387, w3310, IN42[12], w3388, w3389);
  FullAdder U588 (w3389, w3312, IN43[11], w3390, w3391);
  FullAdder U589 (w3391, w3314, IN44[10], w3392, w3393);
  FullAdder U590 (w3393, w3316, IN45[9], w3394, w3395);
  FullAdder U591 (w3395, w3318, IN46[8], w3396, w3397);
  FullAdder U592 (w3397, w3320, IN47[7], w3398, w3399);
  FullAdder U593 (w3399, w3322, IN48[6], w3400, w3401);
  FullAdder U594 (w3401, w3324, IN49[5], w3402, w3403);
  FullAdder U595 (w3403, w3326, IN50[4], w3404, w3405);
  FullAdder U596 (w3405, w3328, IN51[3], w3406, w3407);
  FullAdder U597 (w3407, w3330, IN52[2], w3408, w3409);
  FullAdder U598 (w3409, w3332, IN53[1], w3410, w3411);
  FullAdder U599 (w3411, w3333, IN54[0], w3412, w3413);
  HalfAdder U600 (w3336, IN16[16], Out1[16], w3415);
  FullAdder U601 (w3415, w3338, IN17[16], w3416, w3417);
  FullAdder U602 (w3417, w3340, IN18[16], w3418, w3419);
  FullAdder U603 (w3419, w3342, IN19[16], w3420, w3421);
  FullAdder U604 (w3421, w3344, IN20[16], w3422, w3423);
  FullAdder U605 (w3423, w3346, IN21[16], w3424, w3425);
  FullAdder U606 (w3425, w3348, IN22[16], w3426, w3427);
  FullAdder U607 (w3427, w3350, IN23[16], w3428, w3429);
  FullAdder U608 (w3429, w3352, IN24[16], w3430, w3431);
  FullAdder U609 (w3431, w3354, IN25[16], w3432, w3433);
  FullAdder U610 (w3433, w3356, IN26[16], w3434, w3435);
  FullAdder U611 (w3435, w3358, IN27[16], w3436, w3437);
  FullAdder U612 (w3437, w3360, IN28[16], w3438, w3439);
  FullAdder U613 (w3439, w3362, IN29[16], w3440, w3441);
  FullAdder U614 (w3441, w3364, IN30[16], w3442, w3443);
  FullAdder U615 (w3443, w3366, IN31[16], w3444, w3445);
  FullAdder U616 (w3445, w3368, IN32[16], w3446, w3447);
  FullAdder U617 (w3447, w3370, IN33[16], w3448, w3449);
  FullAdder U618 (w3449, w3372, IN34[16], w3450, w3451);
  FullAdder U619 (w3451, w3374, IN35[16], w3452, w3453);
  FullAdder U620 (w3453, w3376, IN36[16], w3454, w3455);
  FullAdder U621 (w3455, w3378, IN37[16], w3456, w3457);
  FullAdder U622 (w3457, w3380, IN38[16], w3458, w3459);
  FullAdder U623 (w3459, w3382, IN39[16], w3460, w3461);
  FullAdder U624 (w3461, w3384, IN40[16], w3462, w3463);
  FullAdder U625 (w3463, w3386, IN41[14], w3464, w3465);
  FullAdder U626 (w3465, w3388, IN42[13], w3466, w3467);
  FullAdder U627 (w3467, w3390, IN43[12], w3468, w3469);
  FullAdder U628 (w3469, w3392, IN44[11], w3470, w3471);
  FullAdder U629 (w3471, w3394, IN45[10], w3472, w3473);
  FullAdder U630 (w3473, w3396, IN46[9], w3474, w3475);
  FullAdder U631 (w3475, w3398, IN47[8], w3476, w3477);
  FullAdder U632 (w3477, w3400, IN48[7], w3478, w3479);
  FullAdder U633 (w3479, w3402, IN49[6], w3480, w3481);
  FullAdder U634 (w3481, w3404, IN50[5], w3482, w3483);
  FullAdder U635 (w3483, w3406, IN51[4], w3484, w3485);
  FullAdder U636 (w3485, w3408, IN52[3], w3486, w3487);
  FullAdder U637 (w3487, w3410, IN53[2], w3488, w3489);
  FullAdder U638 (w3489, w3412, IN54[1], w3490, w3491);
  FullAdder U639 (w3491, w3413, IN55[0], w3492, w3493);
  HalfAdder U640 (w3416, IN17[17], Out1[17], w3495);
  FullAdder U641 (w3495, w3418, IN18[17], w3496, w3497);
  FullAdder U642 (w3497, w3420, IN19[17], w3498, w3499);
  FullAdder U643 (w3499, w3422, IN20[17], w3500, w3501);
  FullAdder U644 (w3501, w3424, IN21[17], w3502, w3503);
  FullAdder U645 (w3503, w3426, IN22[17], w3504, w3505);
  FullAdder U646 (w3505, w3428, IN23[17], w3506, w3507);
  FullAdder U647 (w3507, w3430, IN24[17], w3508, w3509);
  FullAdder U648 (w3509, w3432, IN25[17], w3510, w3511);
  FullAdder U649 (w3511, w3434, IN26[17], w3512, w3513);
  FullAdder U650 (w3513, w3436, IN27[17], w3514, w3515);
  FullAdder U651 (w3515, w3438, IN28[17], w3516, w3517);
  FullAdder U652 (w3517, w3440, IN29[17], w3518, w3519);
  FullAdder U653 (w3519, w3442, IN30[17], w3520, w3521);
  FullAdder U654 (w3521, w3444, IN31[17], w3522, w3523);
  FullAdder U655 (w3523, w3446, IN32[17], w3524, w3525);
  FullAdder U656 (w3525, w3448, IN33[17], w3526, w3527);
  FullAdder U657 (w3527, w3450, IN34[17], w3528, w3529);
  FullAdder U658 (w3529, w3452, IN35[17], w3530, w3531);
  FullAdder U659 (w3531, w3454, IN36[17], w3532, w3533);
  FullAdder U660 (w3533, w3456, IN37[17], w3534, w3535);
  FullAdder U661 (w3535, w3458, IN38[17], w3536, w3537);
  FullAdder U662 (w3537, w3460, IN39[17], w3538, w3539);
  FullAdder U663 (w3539, w3462, IN40[17], w3540, w3541);
  FullAdder U664 (w3541, w3464, IN41[15], w3542, w3543);
  FullAdder U665 (w3543, w3466, IN42[14], w3544, w3545);
  FullAdder U666 (w3545, w3468, IN43[13], w3546, w3547);
  FullAdder U667 (w3547, w3470, IN44[12], w3548, w3549);
  FullAdder U668 (w3549, w3472, IN45[11], w3550, w3551);
  FullAdder U669 (w3551, w3474, IN46[10], w3552, w3553);
  FullAdder U670 (w3553, w3476, IN47[9], w3554, w3555);
  FullAdder U671 (w3555, w3478, IN48[8], w3556, w3557);
  FullAdder U672 (w3557, w3480, IN49[7], w3558, w3559);
  FullAdder U673 (w3559, w3482, IN50[6], w3560, w3561);
  FullAdder U674 (w3561, w3484, IN51[5], w3562, w3563);
  FullAdder U675 (w3563, w3486, IN52[4], w3564, w3565);
  FullAdder U676 (w3565, w3488, IN53[3], w3566, w3567);
  FullAdder U677 (w3567, w3490, IN54[2], w3568, w3569);
  FullAdder U678 (w3569, w3492, IN55[1], w3570, w3571);
  FullAdder U679 (w3571, w3493, IN56[0], w3572, w3573);
  HalfAdder U680 (w3496, IN18[18], Out1[18], w3575);
  FullAdder U681 (w3575, w3498, IN19[18], w3576, w3577);
  FullAdder U682 (w3577, w3500, IN20[18], w3578, w3579);
  FullAdder U683 (w3579, w3502, IN21[18], w3580, w3581);
  FullAdder U684 (w3581, w3504, IN22[18], w3582, w3583);
  FullAdder U685 (w3583, w3506, IN23[18], w3584, w3585);
  FullAdder U686 (w3585, w3508, IN24[18], w3586, w3587);
  FullAdder U687 (w3587, w3510, IN25[18], w3588, w3589);
  FullAdder U688 (w3589, w3512, IN26[18], w3590, w3591);
  FullAdder U689 (w3591, w3514, IN27[18], w3592, w3593);
  FullAdder U690 (w3593, w3516, IN28[18], w3594, w3595);
  FullAdder U691 (w3595, w3518, IN29[18], w3596, w3597);
  FullAdder U692 (w3597, w3520, IN30[18], w3598, w3599);
  FullAdder U693 (w3599, w3522, IN31[18], w3600, w3601);
  FullAdder U694 (w3601, w3524, IN32[18], w3602, w3603);
  FullAdder U695 (w3603, w3526, IN33[18], w3604, w3605);
  FullAdder U696 (w3605, w3528, IN34[18], w3606, w3607);
  FullAdder U697 (w3607, w3530, IN35[18], w3608, w3609);
  FullAdder U698 (w3609, w3532, IN36[18], w3610, w3611);
  FullAdder U699 (w3611, w3534, IN37[18], w3612, w3613);
  FullAdder U700 (w3613, w3536, IN38[18], w3614, w3615);
  FullAdder U701 (w3615, w3538, IN39[18], w3616, w3617);
  FullAdder U702 (w3617, w3540, IN40[18], w3618, w3619);
  FullAdder U703 (w3619, w3542, IN41[16], w3620, w3621);
  FullAdder U704 (w3621, w3544, IN42[15], w3622, w3623);
  FullAdder U705 (w3623, w3546, IN43[14], w3624, w3625);
  FullAdder U706 (w3625, w3548, IN44[13], w3626, w3627);
  FullAdder U707 (w3627, w3550, IN45[12], w3628, w3629);
  FullAdder U708 (w3629, w3552, IN46[11], w3630, w3631);
  FullAdder U709 (w3631, w3554, IN47[10], w3632, w3633);
  FullAdder U710 (w3633, w3556, IN48[9], w3634, w3635);
  FullAdder U711 (w3635, w3558, IN49[8], w3636, w3637);
  FullAdder U712 (w3637, w3560, IN50[7], w3638, w3639);
  FullAdder U713 (w3639, w3562, IN51[6], w3640, w3641);
  FullAdder U714 (w3641, w3564, IN52[5], w3642, w3643);
  FullAdder U715 (w3643, w3566, IN53[4], w3644, w3645);
  FullAdder U716 (w3645, w3568, IN54[3], w3646, w3647);
  FullAdder U717 (w3647, w3570, IN55[2], w3648, w3649);
  FullAdder U718 (w3649, w3572, IN56[1], w3650, w3651);
  FullAdder U719 (w3651, w3573, IN57[0], w3652, w3653);
  HalfAdder U720 (w3576, IN19[19], Out1[19], w3655);
  FullAdder U721 (w3655, w3578, IN20[19], w3656, w3657);
  FullAdder U722 (w3657, w3580, IN21[19], w3658, w3659);
  FullAdder U723 (w3659, w3582, IN22[19], w3660, w3661);
  FullAdder U724 (w3661, w3584, IN23[19], w3662, w3663);
  FullAdder U725 (w3663, w3586, IN24[19], w3664, w3665);
  FullAdder U726 (w3665, w3588, IN25[19], w3666, w3667);
  FullAdder U727 (w3667, w3590, IN26[19], w3668, w3669);
  FullAdder U728 (w3669, w3592, IN27[19], w3670, w3671);
  FullAdder U729 (w3671, w3594, IN28[19], w3672, w3673);
  FullAdder U730 (w3673, w3596, IN29[19], w3674, w3675);
  FullAdder U731 (w3675, w3598, IN30[19], w3676, w3677);
  FullAdder U732 (w3677, w3600, IN31[19], w3678, w3679);
  FullAdder U733 (w3679, w3602, IN32[19], w3680, w3681);
  FullAdder U734 (w3681, w3604, IN33[19], w3682, w3683);
  FullAdder U735 (w3683, w3606, IN34[19], w3684, w3685);
  FullAdder U736 (w3685, w3608, IN35[19], w3686, w3687);
  FullAdder U737 (w3687, w3610, IN36[19], w3688, w3689);
  FullAdder U738 (w3689, w3612, IN37[19], w3690, w3691);
  FullAdder U739 (w3691, w3614, IN38[19], w3692, w3693);
  FullAdder U740 (w3693, w3616, IN39[19], w3694, w3695);
  FullAdder U741 (w3695, w3618, IN40[19], w3696, w3697);
  FullAdder U742 (w3697, w3620, IN41[17], w3698, w3699);
  FullAdder U743 (w3699, w3622, IN42[16], w3700, w3701);
  FullAdder U744 (w3701, w3624, IN43[15], w3702, w3703);
  FullAdder U745 (w3703, w3626, IN44[14], w3704, w3705);
  FullAdder U746 (w3705, w3628, IN45[13], w3706, w3707);
  FullAdder U747 (w3707, w3630, IN46[12], w3708, w3709);
  FullAdder U748 (w3709, w3632, IN47[11], w3710, w3711);
  FullAdder U749 (w3711, w3634, IN48[10], w3712, w3713);
  FullAdder U750 (w3713, w3636, IN49[9], w3714, w3715);
  FullAdder U751 (w3715, w3638, IN50[8], w3716, w3717);
  FullAdder U752 (w3717, w3640, IN51[7], w3718, w3719);
  FullAdder U753 (w3719, w3642, IN52[6], w3720, w3721);
  FullAdder U754 (w3721, w3644, IN53[5], w3722, w3723);
  FullAdder U755 (w3723, w3646, IN54[4], w3724, w3725);
  FullAdder U756 (w3725, w3648, IN55[3], w3726, w3727);
  FullAdder U757 (w3727, w3650, IN56[2], w3728, w3729);
  FullAdder U758 (w3729, w3652, IN57[1], w3730, w3731);
  FullAdder U759 (w3731, w3653, IN58[0], w3732, w3733);
  HalfAdder U760 (w3656, IN20[20], Out1[20], w3735);
  FullAdder U761 (w3735, w3658, IN21[20], w3736, w3737);
  FullAdder U762 (w3737, w3660, IN22[20], w3738, w3739);
  FullAdder U763 (w3739, w3662, IN23[20], w3740, w3741);
  FullAdder U764 (w3741, w3664, IN24[20], w3742, w3743);
  FullAdder U765 (w3743, w3666, IN25[20], w3744, w3745);
  FullAdder U766 (w3745, w3668, IN26[20], w3746, w3747);
  FullAdder U767 (w3747, w3670, IN27[20], w3748, w3749);
  FullAdder U768 (w3749, w3672, IN28[20], w3750, w3751);
  FullAdder U769 (w3751, w3674, IN29[20], w3752, w3753);
  FullAdder U770 (w3753, w3676, IN30[20], w3754, w3755);
  FullAdder U771 (w3755, w3678, IN31[20], w3756, w3757);
  FullAdder U772 (w3757, w3680, IN32[20], w3758, w3759);
  FullAdder U773 (w3759, w3682, IN33[20], w3760, w3761);
  FullAdder U774 (w3761, w3684, IN34[20], w3762, w3763);
  FullAdder U775 (w3763, w3686, IN35[20], w3764, w3765);
  FullAdder U776 (w3765, w3688, IN36[20], w3766, w3767);
  FullAdder U777 (w3767, w3690, IN37[20], w3768, w3769);
  FullAdder U778 (w3769, w3692, IN38[20], w3770, w3771);
  FullAdder U779 (w3771, w3694, IN39[20], w3772, w3773);
  FullAdder U780 (w3773, w3696, IN40[20], w3774, w3775);
  FullAdder U781 (w3775, w3698, IN41[18], w3776, w3777);
  FullAdder U782 (w3777, w3700, IN42[17], w3778, w3779);
  FullAdder U783 (w3779, w3702, IN43[16], w3780, w3781);
  FullAdder U784 (w3781, w3704, IN44[15], w3782, w3783);
  FullAdder U785 (w3783, w3706, IN45[14], w3784, w3785);
  FullAdder U786 (w3785, w3708, IN46[13], w3786, w3787);
  FullAdder U787 (w3787, w3710, IN47[12], w3788, w3789);
  FullAdder U788 (w3789, w3712, IN48[11], w3790, w3791);
  FullAdder U789 (w3791, w3714, IN49[10], w3792, w3793);
  FullAdder U790 (w3793, w3716, IN50[9], w3794, w3795);
  FullAdder U791 (w3795, w3718, IN51[8], w3796, w3797);
  FullAdder U792 (w3797, w3720, IN52[7], w3798, w3799);
  FullAdder U793 (w3799, w3722, IN53[6], w3800, w3801);
  FullAdder U794 (w3801, w3724, IN54[5], w3802, w3803);
  FullAdder U795 (w3803, w3726, IN55[4], w3804, w3805);
  FullAdder U796 (w3805, w3728, IN56[3], w3806, w3807);
  FullAdder U797 (w3807, w3730, IN57[2], w3808, w3809);
  FullAdder U798 (w3809, w3732, IN58[1], w3810, w3811);
  FullAdder U799 (w3811, w3733, IN59[0], w3812, w3813);
  HalfAdder U800 (w3736, IN21[21], Out1[21], w3815);
  FullAdder U801 (w3815, w3738, IN22[21], w3816, w3817);
  FullAdder U802 (w3817, w3740, IN23[21], w3818, w3819);
  FullAdder U803 (w3819, w3742, IN24[21], w3820, w3821);
  FullAdder U804 (w3821, w3744, IN25[21], w3822, w3823);
  FullAdder U805 (w3823, w3746, IN26[21], w3824, w3825);
  FullAdder U806 (w3825, w3748, IN27[21], w3826, w3827);
  FullAdder U807 (w3827, w3750, IN28[21], w3828, w3829);
  FullAdder U808 (w3829, w3752, IN29[21], w3830, w3831);
  FullAdder U809 (w3831, w3754, IN30[21], w3832, w3833);
  FullAdder U810 (w3833, w3756, IN31[21], w3834, w3835);
  FullAdder U811 (w3835, w3758, IN32[21], w3836, w3837);
  FullAdder U812 (w3837, w3760, IN33[21], w3838, w3839);
  FullAdder U813 (w3839, w3762, IN34[21], w3840, w3841);
  FullAdder U814 (w3841, w3764, IN35[21], w3842, w3843);
  FullAdder U815 (w3843, w3766, IN36[21], w3844, w3845);
  FullAdder U816 (w3845, w3768, IN37[21], w3846, w3847);
  FullAdder U817 (w3847, w3770, IN38[21], w3848, w3849);
  FullAdder U818 (w3849, w3772, IN39[21], w3850, w3851);
  FullAdder U819 (w3851, w3774, IN40[21], w3852, w3853);
  FullAdder U820 (w3853, w3776, IN41[19], w3854, w3855);
  FullAdder U821 (w3855, w3778, IN42[18], w3856, w3857);
  FullAdder U822 (w3857, w3780, IN43[17], w3858, w3859);
  FullAdder U823 (w3859, w3782, IN44[16], w3860, w3861);
  FullAdder U824 (w3861, w3784, IN45[15], w3862, w3863);
  FullAdder U825 (w3863, w3786, IN46[14], w3864, w3865);
  FullAdder U826 (w3865, w3788, IN47[13], w3866, w3867);
  FullAdder U827 (w3867, w3790, IN48[12], w3868, w3869);
  FullAdder U828 (w3869, w3792, IN49[11], w3870, w3871);
  FullAdder U829 (w3871, w3794, IN50[10], w3872, w3873);
  FullAdder U830 (w3873, w3796, IN51[9], w3874, w3875);
  FullAdder U831 (w3875, w3798, IN52[8], w3876, w3877);
  FullAdder U832 (w3877, w3800, IN53[7], w3878, w3879);
  FullAdder U833 (w3879, w3802, IN54[6], w3880, w3881);
  FullAdder U834 (w3881, w3804, IN55[5], w3882, w3883);
  FullAdder U835 (w3883, w3806, IN56[4], w3884, w3885);
  FullAdder U836 (w3885, w3808, IN57[3], w3886, w3887);
  FullAdder U837 (w3887, w3810, IN58[2], w3888, w3889);
  FullAdder U838 (w3889, w3812, IN59[1], w3890, w3891);
  FullAdder U839 (w3891, w3813, IN60[0], w3892, w3893);
  HalfAdder U840 (w3816, IN22[22], Out1[22], w3895);
  FullAdder U841 (w3895, w3818, IN23[22], w3896, w3897);
  FullAdder U842 (w3897, w3820, IN24[22], w3898, w3899);
  FullAdder U843 (w3899, w3822, IN25[22], w3900, w3901);
  FullAdder U844 (w3901, w3824, IN26[22], w3902, w3903);
  FullAdder U845 (w3903, w3826, IN27[22], w3904, w3905);
  FullAdder U846 (w3905, w3828, IN28[22], w3906, w3907);
  FullAdder U847 (w3907, w3830, IN29[22], w3908, w3909);
  FullAdder U848 (w3909, w3832, IN30[22], w3910, w3911);
  FullAdder U849 (w3911, w3834, IN31[22], w3912, w3913);
  FullAdder U850 (w3913, w3836, IN32[22], w3914, w3915);
  FullAdder U851 (w3915, w3838, IN33[22], w3916, w3917);
  FullAdder U852 (w3917, w3840, IN34[22], w3918, w3919);
  FullAdder U853 (w3919, w3842, IN35[22], w3920, w3921);
  FullAdder U854 (w3921, w3844, IN36[22], w3922, w3923);
  FullAdder U855 (w3923, w3846, IN37[22], w3924, w3925);
  FullAdder U856 (w3925, w3848, IN38[22], w3926, w3927);
  FullAdder U857 (w3927, w3850, IN39[22], w3928, w3929);
  FullAdder U858 (w3929, w3852, IN40[22], w3930, w3931);
  FullAdder U859 (w3931, w3854, IN41[20], w3932, w3933);
  FullAdder U860 (w3933, w3856, IN42[19], w3934, w3935);
  FullAdder U861 (w3935, w3858, IN43[18], w3936, w3937);
  FullAdder U862 (w3937, w3860, IN44[17], w3938, w3939);
  FullAdder U863 (w3939, w3862, IN45[16], w3940, w3941);
  FullAdder U864 (w3941, w3864, IN46[15], w3942, w3943);
  FullAdder U865 (w3943, w3866, IN47[14], w3944, w3945);
  FullAdder U866 (w3945, w3868, IN48[13], w3946, w3947);
  FullAdder U867 (w3947, w3870, IN49[12], w3948, w3949);
  FullAdder U868 (w3949, w3872, IN50[11], w3950, w3951);
  FullAdder U869 (w3951, w3874, IN51[10], w3952, w3953);
  FullAdder U870 (w3953, w3876, IN52[9], w3954, w3955);
  FullAdder U871 (w3955, w3878, IN53[8], w3956, w3957);
  FullAdder U872 (w3957, w3880, IN54[7], w3958, w3959);
  FullAdder U873 (w3959, w3882, IN55[6], w3960, w3961);
  FullAdder U874 (w3961, w3884, IN56[5], w3962, w3963);
  FullAdder U875 (w3963, w3886, IN57[4], w3964, w3965);
  FullAdder U876 (w3965, w3888, IN58[3], w3966, w3967);
  FullAdder U877 (w3967, w3890, IN59[2], w3968, w3969);
  FullAdder U878 (w3969, w3892, IN60[1], w3970, w3971);
  FullAdder U879 (w3971, w3893, IN61[0], w3972, w3973);
  HalfAdder U880 (w3896, IN23[23], Out1[23], w3975);
  FullAdder U881 (w3975, w3898, IN24[23], w3976, w3977);
  FullAdder U882 (w3977, w3900, IN25[23], w3978, w3979);
  FullAdder U883 (w3979, w3902, IN26[23], w3980, w3981);
  FullAdder U884 (w3981, w3904, IN27[23], w3982, w3983);
  FullAdder U885 (w3983, w3906, IN28[23], w3984, w3985);
  FullAdder U886 (w3985, w3908, IN29[23], w3986, w3987);
  FullAdder U887 (w3987, w3910, IN30[23], w3988, w3989);
  FullAdder U888 (w3989, w3912, IN31[23], w3990, w3991);
  FullAdder U889 (w3991, w3914, IN32[23], w3992, w3993);
  FullAdder U890 (w3993, w3916, IN33[23], w3994, w3995);
  FullAdder U891 (w3995, w3918, IN34[23], w3996, w3997);
  FullAdder U892 (w3997, w3920, IN35[23], w3998, w3999);
  FullAdder U893 (w3999, w3922, IN36[23], w4000, w4001);
  FullAdder U894 (w4001, w3924, IN37[23], w4002, w4003);
  FullAdder U895 (w4003, w3926, IN38[23], w4004, w4005);
  FullAdder U896 (w4005, w3928, IN39[23], w4006, w4007);
  FullAdder U897 (w4007, w3930, IN40[23], w4008, w4009);
  FullAdder U898 (w4009, w3932, IN41[21], w4010, w4011);
  FullAdder U899 (w4011, w3934, IN42[20], w4012, w4013);
  FullAdder U900 (w4013, w3936, IN43[19], w4014, w4015);
  FullAdder U901 (w4015, w3938, IN44[18], w4016, w4017);
  FullAdder U902 (w4017, w3940, IN45[17], w4018, w4019);
  FullAdder U903 (w4019, w3942, IN46[16], w4020, w4021);
  FullAdder U904 (w4021, w3944, IN47[15], w4022, w4023);
  FullAdder U905 (w4023, w3946, IN48[14], w4024, w4025);
  FullAdder U906 (w4025, w3948, IN49[13], w4026, w4027);
  FullAdder U907 (w4027, w3950, IN50[12], w4028, w4029);
  FullAdder U908 (w4029, w3952, IN51[11], w4030, w4031);
  FullAdder U909 (w4031, w3954, IN52[10], w4032, w4033);
  FullAdder U910 (w4033, w3956, IN53[9], w4034, w4035);
  FullAdder U911 (w4035, w3958, IN54[8], w4036, w4037);
  FullAdder U912 (w4037, w3960, IN55[7], w4038, w4039);
  FullAdder U913 (w4039, w3962, IN56[6], w4040, w4041);
  FullAdder U914 (w4041, w3964, IN57[5], w4042, w4043);
  FullAdder U915 (w4043, w3966, IN58[4], w4044, w4045);
  FullAdder U916 (w4045, w3968, IN59[3], w4046, w4047);
  FullAdder U917 (w4047, w3970, IN60[2], w4048, w4049);
  FullAdder U918 (w4049, w3972, IN61[1], w4050, w4051);
  FullAdder U919 (w4051, w3973, IN62[0], w4052, w4053);
  HalfAdder U920 (w3976, IN24[24], Out1[24], w4055);
  FullAdder U921 (w4055, w3978, IN25[24], w4056, w4057);
  FullAdder U922 (w4057, w3980, IN26[24], w4058, w4059);
  FullAdder U923 (w4059, w3982, IN27[24], w4060, w4061);
  FullAdder U924 (w4061, w3984, IN28[24], w4062, w4063);
  FullAdder U925 (w4063, w3986, IN29[24], w4064, w4065);
  FullAdder U926 (w4065, w3988, IN30[24], w4066, w4067);
  FullAdder U927 (w4067, w3990, IN31[24], w4068, w4069);
  FullAdder U928 (w4069, w3992, IN32[24], w4070, w4071);
  FullAdder U929 (w4071, w3994, IN33[24], w4072, w4073);
  FullAdder U930 (w4073, w3996, IN34[24], w4074, w4075);
  FullAdder U931 (w4075, w3998, IN35[24], w4076, w4077);
  FullAdder U932 (w4077, w4000, IN36[24], w4078, w4079);
  FullAdder U933 (w4079, w4002, IN37[24], w4080, w4081);
  FullAdder U934 (w4081, w4004, IN38[24], w4082, w4083);
  FullAdder U935 (w4083, w4006, IN39[24], w4084, w4085);
  FullAdder U936 (w4085, w4008, IN40[24], w4086, w4087);
  FullAdder U937 (w4087, w4010, IN41[22], w4088, w4089);
  FullAdder U938 (w4089, w4012, IN42[21], w4090, w4091);
  FullAdder U939 (w4091, w4014, IN43[20], w4092, w4093);
  FullAdder U940 (w4093, w4016, IN44[19], w4094, w4095);
  FullAdder U941 (w4095, w4018, IN45[18], w4096, w4097);
  FullAdder U942 (w4097, w4020, IN46[17], w4098, w4099);
  FullAdder U943 (w4099, w4022, IN47[16], w4100, w4101);
  FullAdder U944 (w4101, w4024, IN48[15], w4102, w4103);
  FullAdder U945 (w4103, w4026, IN49[14], w4104, w4105);
  FullAdder U946 (w4105, w4028, IN50[13], w4106, w4107);
  FullAdder U947 (w4107, w4030, IN51[12], w4108, w4109);
  FullAdder U948 (w4109, w4032, IN52[11], w4110, w4111);
  FullAdder U949 (w4111, w4034, IN53[10], w4112, w4113);
  FullAdder U950 (w4113, w4036, IN54[9], w4114, w4115);
  FullAdder U951 (w4115, w4038, IN55[8], w4116, w4117);
  FullAdder U952 (w4117, w4040, IN56[7], w4118, w4119);
  FullAdder U953 (w4119, w4042, IN57[6], w4120, w4121);
  FullAdder U954 (w4121, w4044, IN58[5], w4122, w4123);
  FullAdder U955 (w4123, w4046, IN59[4], w4124, w4125);
  FullAdder U956 (w4125, w4048, IN60[3], w4126, w4127);
  FullAdder U957 (w4127, w4050, IN61[2], w4128, w4129);
  FullAdder U958 (w4129, w4052, IN62[1], w4130, w4131);
  FullAdder U959 (w4131, w4053, IN63[0], w4132, w4133);
  HalfAdder U960 (w4056, IN25[25], Out1[25], w4135);
  FullAdder U961 (w4135, w4058, IN26[25], w4136, w4137);
  FullAdder U962 (w4137, w4060, IN27[25], w4138, w4139);
  FullAdder U963 (w4139, w4062, IN28[25], w4140, w4141);
  FullAdder U964 (w4141, w4064, IN29[25], w4142, w4143);
  FullAdder U965 (w4143, w4066, IN30[25], w4144, w4145);
  FullAdder U966 (w4145, w4068, IN31[25], w4146, w4147);
  FullAdder U967 (w4147, w4070, IN32[25], w4148, w4149);
  FullAdder U968 (w4149, w4072, IN33[25], w4150, w4151);
  FullAdder U969 (w4151, w4074, IN34[25], w4152, w4153);
  FullAdder U970 (w4153, w4076, IN35[25], w4154, w4155);
  FullAdder U971 (w4155, w4078, IN36[25], w4156, w4157);
  FullAdder U972 (w4157, w4080, IN37[25], w4158, w4159);
  FullAdder U973 (w4159, w4082, IN38[25], w4160, w4161);
  FullAdder U974 (w4161, w4084, IN39[25], w4162, w4163);
  FullAdder U975 (w4163, w4086, IN40[25], w4164, w4165);
  FullAdder U976 (w4165, w4088, IN41[23], w4166, w4167);
  FullAdder U977 (w4167, w4090, IN42[22], w4168, w4169);
  FullAdder U978 (w4169, w4092, IN43[21], w4170, w4171);
  FullAdder U979 (w4171, w4094, IN44[20], w4172, w4173);
  FullAdder U980 (w4173, w4096, IN45[19], w4174, w4175);
  FullAdder U981 (w4175, w4098, IN46[18], w4176, w4177);
  FullAdder U982 (w4177, w4100, IN47[17], w4178, w4179);
  FullAdder U983 (w4179, w4102, IN48[16], w4180, w4181);
  FullAdder U984 (w4181, w4104, IN49[15], w4182, w4183);
  FullAdder U985 (w4183, w4106, IN50[14], w4184, w4185);
  FullAdder U986 (w4185, w4108, IN51[13], w4186, w4187);
  FullAdder U987 (w4187, w4110, IN52[12], w4188, w4189);
  FullAdder U988 (w4189, w4112, IN53[11], w4190, w4191);
  FullAdder U989 (w4191, w4114, IN54[10], w4192, w4193);
  FullAdder U990 (w4193, w4116, IN55[9], w4194, w4195);
  FullAdder U991 (w4195, w4118, IN56[8], w4196, w4197);
  FullAdder U992 (w4197, w4120, IN57[7], w4198, w4199);
  FullAdder U993 (w4199, w4122, IN58[6], w4200, w4201);
  FullAdder U994 (w4201, w4124, IN59[5], w4202, w4203);
  FullAdder U995 (w4203, w4126, IN60[4], w4204, w4205);
  FullAdder U996 (w4205, w4128, IN61[3], w4206, w4207);
  FullAdder U997 (w4207, w4130, IN62[2], w4208, w4209);
  FullAdder U998 (w4209, w4132, IN63[1], w4210, w4211);
  FullAdder U999 (w4211, w4133, IN64[0], w4212, w4213);
  HalfAdder U1000 (w4136, IN26[26], Out1[26], w4215);
  FullAdder U1001 (w4215, w4138, IN27[26], w4216, w4217);
  FullAdder U1002 (w4217, w4140, IN28[26], w4218, w4219);
  FullAdder U1003 (w4219, w4142, IN29[26], w4220, w4221);
  FullAdder U1004 (w4221, w4144, IN30[26], w4222, w4223);
  FullAdder U1005 (w4223, w4146, IN31[26], w4224, w4225);
  FullAdder U1006 (w4225, w4148, IN32[26], w4226, w4227);
  FullAdder U1007 (w4227, w4150, IN33[26], w4228, w4229);
  FullAdder U1008 (w4229, w4152, IN34[26], w4230, w4231);
  FullAdder U1009 (w4231, w4154, IN35[26], w4232, w4233);
  FullAdder U1010 (w4233, w4156, IN36[26], w4234, w4235);
  FullAdder U1011 (w4235, w4158, IN37[26], w4236, w4237);
  FullAdder U1012 (w4237, w4160, IN38[26], w4238, w4239);
  FullAdder U1013 (w4239, w4162, IN39[26], w4240, w4241);
  FullAdder U1014 (w4241, w4164, IN40[26], w4242, w4243);
  FullAdder U1015 (w4243, w4166, IN41[24], w4244, w4245);
  FullAdder U1016 (w4245, w4168, IN42[23], w4246, w4247);
  FullAdder U1017 (w4247, w4170, IN43[22], w4248, w4249);
  FullAdder U1018 (w4249, w4172, IN44[21], w4250, w4251);
  FullAdder U1019 (w4251, w4174, IN45[20], w4252, w4253);
  FullAdder U1020 (w4253, w4176, IN46[19], w4254, w4255);
  FullAdder U1021 (w4255, w4178, IN47[18], w4256, w4257);
  FullAdder U1022 (w4257, w4180, IN48[17], w4258, w4259);
  FullAdder U1023 (w4259, w4182, IN49[16], w4260, w4261);
  FullAdder U1024 (w4261, w4184, IN50[15], w4262, w4263);
  FullAdder U1025 (w4263, w4186, IN51[14], w4264, w4265);
  FullAdder U1026 (w4265, w4188, IN52[13], w4266, w4267);
  FullAdder U1027 (w4267, w4190, IN53[12], w4268, w4269);
  FullAdder U1028 (w4269, w4192, IN54[11], w4270, w4271);
  FullAdder U1029 (w4271, w4194, IN55[10], w4272, w4273);
  FullAdder U1030 (w4273, w4196, IN56[9], w4274, w4275);
  FullAdder U1031 (w4275, w4198, IN57[8], w4276, w4277);
  FullAdder U1032 (w4277, w4200, IN58[7], w4278, w4279);
  FullAdder U1033 (w4279, w4202, IN59[6], w4280, w4281);
  FullAdder U1034 (w4281, w4204, IN60[5], w4282, w4283);
  FullAdder U1035 (w4283, w4206, IN61[4], w4284, w4285);
  FullAdder U1036 (w4285, w4208, IN62[3], w4286, w4287);
  FullAdder U1037 (w4287, w4210, IN63[2], w4288, w4289);
  FullAdder U1038 (w4289, w4212, IN64[1], w4290, w4291);
  FullAdder U1039 (w4291, w4213, IN65[0], w4292, w4293);
  HalfAdder U1040 (w4216, IN27[27], Out1[27], w4295);
  FullAdder U1041 (w4295, w4218, IN28[27], w4296, w4297);
  FullAdder U1042 (w4297, w4220, IN29[27], w4298, w4299);
  FullAdder U1043 (w4299, w4222, IN30[27], w4300, w4301);
  FullAdder U1044 (w4301, w4224, IN31[27], w4302, w4303);
  FullAdder U1045 (w4303, w4226, IN32[27], w4304, w4305);
  FullAdder U1046 (w4305, w4228, IN33[27], w4306, w4307);
  FullAdder U1047 (w4307, w4230, IN34[27], w4308, w4309);
  FullAdder U1048 (w4309, w4232, IN35[27], w4310, w4311);
  FullAdder U1049 (w4311, w4234, IN36[27], w4312, w4313);
  FullAdder U1050 (w4313, w4236, IN37[27], w4314, w4315);
  FullAdder U1051 (w4315, w4238, IN38[27], w4316, w4317);
  FullAdder U1052 (w4317, w4240, IN39[27], w4318, w4319);
  FullAdder U1053 (w4319, w4242, IN40[27], w4320, w4321);
  FullAdder U1054 (w4321, w4244, IN41[25], w4322, w4323);
  FullAdder U1055 (w4323, w4246, IN42[24], w4324, w4325);
  FullAdder U1056 (w4325, w4248, IN43[23], w4326, w4327);
  FullAdder U1057 (w4327, w4250, IN44[22], w4328, w4329);
  FullAdder U1058 (w4329, w4252, IN45[21], w4330, w4331);
  FullAdder U1059 (w4331, w4254, IN46[20], w4332, w4333);
  FullAdder U1060 (w4333, w4256, IN47[19], w4334, w4335);
  FullAdder U1061 (w4335, w4258, IN48[18], w4336, w4337);
  FullAdder U1062 (w4337, w4260, IN49[17], w4338, w4339);
  FullAdder U1063 (w4339, w4262, IN50[16], w4340, w4341);
  FullAdder U1064 (w4341, w4264, IN51[15], w4342, w4343);
  FullAdder U1065 (w4343, w4266, IN52[14], w4344, w4345);
  FullAdder U1066 (w4345, w4268, IN53[13], w4346, w4347);
  FullAdder U1067 (w4347, w4270, IN54[12], w4348, w4349);
  FullAdder U1068 (w4349, w4272, IN55[11], w4350, w4351);
  FullAdder U1069 (w4351, w4274, IN56[10], w4352, w4353);
  FullAdder U1070 (w4353, w4276, IN57[9], w4354, w4355);
  FullAdder U1071 (w4355, w4278, IN58[8], w4356, w4357);
  FullAdder U1072 (w4357, w4280, IN59[7], w4358, w4359);
  FullAdder U1073 (w4359, w4282, IN60[6], w4360, w4361);
  FullAdder U1074 (w4361, w4284, IN61[5], w4362, w4363);
  FullAdder U1075 (w4363, w4286, IN62[4], w4364, w4365);
  FullAdder U1076 (w4365, w4288, IN63[3], w4366, w4367);
  FullAdder U1077 (w4367, w4290, IN64[2], w4368, w4369);
  FullAdder U1078 (w4369, w4292, IN65[1], w4370, w4371);
  FullAdder U1079 (w4371, w4293, IN66[0], w4372, w4373);
  HalfAdder U1080 (w4296, IN28[28], Out1[28], w4375);
  FullAdder U1081 (w4375, w4298, IN29[28], w4376, w4377);
  FullAdder U1082 (w4377, w4300, IN30[28], w4378, w4379);
  FullAdder U1083 (w4379, w4302, IN31[28], w4380, w4381);
  FullAdder U1084 (w4381, w4304, IN32[28], w4382, w4383);
  FullAdder U1085 (w4383, w4306, IN33[28], w4384, w4385);
  FullAdder U1086 (w4385, w4308, IN34[28], w4386, w4387);
  FullAdder U1087 (w4387, w4310, IN35[28], w4388, w4389);
  FullAdder U1088 (w4389, w4312, IN36[28], w4390, w4391);
  FullAdder U1089 (w4391, w4314, IN37[28], w4392, w4393);
  FullAdder U1090 (w4393, w4316, IN38[28], w4394, w4395);
  FullAdder U1091 (w4395, w4318, IN39[28], w4396, w4397);
  FullAdder U1092 (w4397, w4320, IN40[28], w4398, w4399);
  FullAdder U1093 (w4399, w4322, IN41[26], w4400, w4401);
  FullAdder U1094 (w4401, w4324, IN42[25], w4402, w4403);
  FullAdder U1095 (w4403, w4326, IN43[24], w4404, w4405);
  FullAdder U1096 (w4405, w4328, IN44[23], w4406, w4407);
  FullAdder U1097 (w4407, w4330, IN45[22], w4408, w4409);
  FullAdder U1098 (w4409, w4332, IN46[21], w4410, w4411);
  FullAdder U1099 (w4411, w4334, IN47[20], w4412, w4413);
  FullAdder U1100 (w4413, w4336, IN48[19], w4414, w4415);
  FullAdder U1101 (w4415, w4338, IN49[18], w4416, w4417);
  FullAdder U1102 (w4417, w4340, IN50[17], w4418, w4419);
  FullAdder U1103 (w4419, w4342, IN51[16], w4420, w4421);
  FullAdder U1104 (w4421, w4344, IN52[15], w4422, w4423);
  FullAdder U1105 (w4423, w4346, IN53[14], w4424, w4425);
  FullAdder U1106 (w4425, w4348, IN54[13], w4426, w4427);
  FullAdder U1107 (w4427, w4350, IN55[12], w4428, w4429);
  FullAdder U1108 (w4429, w4352, IN56[11], w4430, w4431);
  FullAdder U1109 (w4431, w4354, IN57[10], w4432, w4433);
  FullAdder U1110 (w4433, w4356, IN58[9], w4434, w4435);
  FullAdder U1111 (w4435, w4358, IN59[8], w4436, w4437);
  FullAdder U1112 (w4437, w4360, IN60[7], w4438, w4439);
  FullAdder U1113 (w4439, w4362, IN61[6], w4440, w4441);
  FullAdder U1114 (w4441, w4364, IN62[5], w4442, w4443);
  FullAdder U1115 (w4443, w4366, IN63[4], w4444, w4445);
  FullAdder U1116 (w4445, w4368, IN64[3], w4446, w4447);
  FullAdder U1117 (w4447, w4370, IN65[2], w4448, w4449);
  FullAdder U1118 (w4449, w4372, IN66[1], w4450, w4451);
  FullAdder U1119 (w4451, w4373, IN67[0], w4452, w4453);
  HalfAdder U1120 (w4376, IN29[29], Out1[29], w4455);
  FullAdder U1121 (w4455, w4378, IN30[29], w4456, w4457);
  FullAdder U1122 (w4457, w4380, IN31[29], w4458, w4459);
  FullAdder U1123 (w4459, w4382, IN32[29], w4460, w4461);
  FullAdder U1124 (w4461, w4384, IN33[29], w4462, w4463);
  FullAdder U1125 (w4463, w4386, IN34[29], w4464, w4465);
  FullAdder U1126 (w4465, w4388, IN35[29], w4466, w4467);
  FullAdder U1127 (w4467, w4390, IN36[29], w4468, w4469);
  FullAdder U1128 (w4469, w4392, IN37[29], w4470, w4471);
  FullAdder U1129 (w4471, w4394, IN38[29], w4472, w4473);
  FullAdder U1130 (w4473, w4396, IN39[29], w4474, w4475);
  FullAdder U1131 (w4475, w4398, IN40[29], w4476, w4477);
  FullAdder U1132 (w4477, w4400, IN41[27], w4478, w4479);
  FullAdder U1133 (w4479, w4402, IN42[26], w4480, w4481);
  FullAdder U1134 (w4481, w4404, IN43[25], w4482, w4483);
  FullAdder U1135 (w4483, w4406, IN44[24], w4484, w4485);
  FullAdder U1136 (w4485, w4408, IN45[23], w4486, w4487);
  FullAdder U1137 (w4487, w4410, IN46[22], w4488, w4489);
  FullAdder U1138 (w4489, w4412, IN47[21], w4490, w4491);
  FullAdder U1139 (w4491, w4414, IN48[20], w4492, w4493);
  FullAdder U1140 (w4493, w4416, IN49[19], w4494, w4495);
  FullAdder U1141 (w4495, w4418, IN50[18], w4496, w4497);
  FullAdder U1142 (w4497, w4420, IN51[17], w4498, w4499);
  FullAdder U1143 (w4499, w4422, IN52[16], w4500, w4501);
  FullAdder U1144 (w4501, w4424, IN53[15], w4502, w4503);
  FullAdder U1145 (w4503, w4426, IN54[14], w4504, w4505);
  FullAdder U1146 (w4505, w4428, IN55[13], w4506, w4507);
  FullAdder U1147 (w4507, w4430, IN56[12], w4508, w4509);
  FullAdder U1148 (w4509, w4432, IN57[11], w4510, w4511);
  FullAdder U1149 (w4511, w4434, IN58[10], w4512, w4513);
  FullAdder U1150 (w4513, w4436, IN59[9], w4514, w4515);
  FullAdder U1151 (w4515, w4438, IN60[8], w4516, w4517);
  FullAdder U1152 (w4517, w4440, IN61[7], w4518, w4519);
  FullAdder U1153 (w4519, w4442, IN62[6], w4520, w4521);
  FullAdder U1154 (w4521, w4444, IN63[5], w4522, w4523);
  FullAdder U1155 (w4523, w4446, IN64[4], w4524, w4525);
  FullAdder U1156 (w4525, w4448, IN65[3], w4526, w4527);
  FullAdder U1157 (w4527, w4450, IN66[2], w4528, w4529);
  FullAdder U1158 (w4529, w4452, IN67[1], w4530, w4531);
  FullAdder U1159 (w4531, w4453, IN68[0], w4532, w4533);
  HalfAdder U1160 (w4456, IN30[30], Out1[30], w4535);
  FullAdder U1161 (w4535, w4458, IN31[30], w4536, w4537);
  FullAdder U1162 (w4537, w4460, IN32[30], w4538, w4539);
  FullAdder U1163 (w4539, w4462, IN33[30], w4540, w4541);
  FullAdder U1164 (w4541, w4464, IN34[30], w4542, w4543);
  FullAdder U1165 (w4543, w4466, IN35[30], w4544, w4545);
  FullAdder U1166 (w4545, w4468, IN36[30], w4546, w4547);
  FullAdder U1167 (w4547, w4470, IN37[30], w4548, w4549);
  FullAdder U1168 (w4549, w4472, IN38[30], w4550, w4551);
  FullAdder U1169 (w4551, w4474, IN39[30], w4552, w4553);
  FullAdder U1170 (w4553, w4476, IN40[30], w4554, w4555);
  FullAdder U1171 (w4555, w4478, IN41[28], w4556, w4557);
  FullAdder U1172 (w4557, w4480, IN42[27], w4558, w4559);
  FullAdder U1173 (w4559, w4482, IN43[26], w4560, w4561);
  FullAdder U1174 (w4561, w4484, IN44[25], w4562, w4563);
  FullAdder U1175 (w4563, w4486, IN45[24], w4564, w4565);
  FullAdder U1176 (w4565, w4488, IN46[23], w4566, w4567);
  FullAdder U1177 (w4567, w4490, IN47[22], w4568, w4569);
  FullAdder U1178 (w4569, w4492, IN48[21], w4570, w4571);
  FullAdder U1179 (w4571, w4494, IN49[20], w4572, w4573);
  FullAdder U1180 (w4573, w4496, IN50[19], w4574, w4575);
  FullAdder U1181 (w4575, w4498, IN51[18], w4576, w4577);
  FullAdder U1182 (w4577, w4500, IN52[17], w4578, w4579);
  FullAdder U1183 (w4579, w4502, IN53[16], w4580, w4581);
  FullAdder U1184 (w4581, w4504, IN54[15], w4582, w4583);
  FullAdder U1185 (w4583, w4506, IN55[14], w4584, w4585);
  FullAdder U1186 (w4585, w4508, IN56[13], w4586, w4587);
  FullAdder U1187 (w4587, w4510, IN57[12], w4588, w4589);
  FullAdder U1188 (w4589, w4512, IN58[11], w4590, w4591);
  FullAdder U1189 (w4591, w4514, IN59[10], w4592, w4593);
  FullAdder U1190 (w4593, w4516, IN60[9], w4594, w4595);
  FullAdder U1191 (w4595, w4518, IN61[8], w4596, w4597);
  FullAdder U1192 (w4597, w4520, IN62[7], w4598, w4599);
  FullAdder U1193 (w4599, w4522, IN63[6], w4600, w4601);
  FullAdder U1194 (w4601, w4524, IN64[5], w4602, w4603);
  FullAdder U1195 (w4603, w4526, IN65[4], w4604, w4605);
  FullAdder U1196 (w4605, w4528, IN66[3], w4606, w4607);
  FullAdder U1197 (w4607, w4530, IN67[2], w4608, w4609);
  FullAdder U1198 (w4609, w4532, IN68[1], w4610, w4611);
  FullAdder U1199 (w4611, w4533, IN69[0], w4612, w4613);
  HalfAdder U1200 (w4536, IN31[31], Out1[31], w4615);
  FullAdder U1201 (w4615, w4538, IN32[31], w4616, w4617);
  FullAdder U1202 (w4617, w4540, IN33[31], w4618, w4619);
  FullAdder U1203 (w4619, w4542, IN34[31], w4620, w4621);
  FullAdder U1204 (w4621, w4544, IN35[31], w4622, w4623);
  FullAdder U1205 (w4623, w4546, IN36[31], w4624, w4625);
  FullAdder U1206 (w4625, w4548, IN37[31], w4626, w4627);
  FullAdder U1207 (w4627, w4550, IN38[31], w4628, w4629);
  FullAdder U1208 (w4629, w4552, IN39[31], w4630, w4631);
  FullAdder U1209 (w4631, w4554, IN40[31], w4632, w4633);
  FullAdder U1210 (w4633, w4556, IN41[29], w4634, w4635);
  FullAdder U1211 (w4635, w4558, IN42[28], w4636, w4637);
  FullAdder U1212 (w4637, w4560, IN43[27], w4638, w4639);
  FullAdder U1213 (w4639, w4562, IN44[26], w4640, w4641);
  FullAdder U1214 (w4641, w4564, IN45[25], w4642, w4643);
  FullAdder U1215 (w4643, w4566, IN46[24], w4644, w4645);
  FullAdder U1216 (w4645, w4568, IN47[23], w4646, w4647);
  FullAdder U1217 (w4647, w4570, IN48[22], w4648, w4649);
  FullAdder U1218 (w4649, w4572, IN49[21], w4650, w4651);
  FullAdder U1219 (w4651, w4574, IN50[20], w4652, w4653);
  FullAdder U1220 (w4653, w4576, IN51[19], w4654, w4655);
  FullAdder U1221 (w4655, w4578, IN52[18], w4656, w4657);
  FullAdder U1222 (w4657, w4580, IN53[17], w4658, w4659);
  FullAdder U1223 (w4659, w4582, IN54[16], w4660, w4661);
  FullAdder U1224 (w4661, w4584, IN55[15], w4662, w4663);
  FullAdder U1225 (w4663, w4586, IN56[14], w4664, w4665);
  FullAdder U1226 (w4665, w4588, IN57[13], w4666, w4667);
  FullAdder U1227 (w4667, w4590, IN58[12], w4668, w4669);
  FullAdder U1228 (w4669, w4592, IN59[11], w4670, w4671);
  FullAdder U1229 (w4671, w4594, IN60[10], w4672, w4673);
  FullAdder U1230 (w4673, w4596, IN61[9], w4674, w4675);
  FullAdder U1231 (w4675, w4598, IN62[8], w4676, w4677);
  FullAdder U1232 (w4677, w4600, IN63[7], w4678, w4679);
  FullAdder U1233 (w4679, w4602, IN64[6], w4680, w4681);
  FullAdder U1234 (w4681, w4604, IN65[5], w4682, w4683);
  FullAdder U1235 (w4683, w4606, IN66[4], w4684, w4685);
  FullAdder U1236 (w4685, w4608, IN67[3], w4686, w4687);
  FullAdder U1237 (w4687, w4610, IN68[2], w4688, w4689);
  FullAdder U1238 (w4689, w4612, IN69[1], w4690, w4691);
  FullAdder U1239 (w4691, w4613, IN70[0], w4692, w4693);
  HalfAdder U1240 (w4616, IN32[32], Out1[32], w4695);
  FullAdder U1241 (w4695, w4618, IN33[32], w4696, w4697);
  FullAdder U1242 (w4697, w4620, IN34[32], w4698, w4699);
  FullAdder U1243 (w4699, w4622, IN35[32], w4700, w4701);
  FullAdder U1244 (w4701, w4624, IN36[32], w4702, w4703);
  FullAdder U1245 (w4703, w4626, IN37[32], w4704, w4705);
  FullAdder U1246 (w4705, w4628, IN38[32], w4706, w4707);
  FullAdder U1247 (w4707, w4630, IN39[32], w4708, w4709);
  FullAdder U1248 (w4709, w4632, IN40[32], w4710, w4711);
  FullAdder U1249 (w4711, w4634, IN41[30], w4712, w4713);
  FullAdder U1250 (w4713, w4636, IN42[29], w4714, w4715);
  FullAdder U1251 (w4715, w4638, IN43[28], w4716, w4717);
  FullAdder U1252 (w4717, w4640, IN44[27], w4718, w4719);
  FullAdder U1253 (w4719, w4642, IN45[26], w4720, w4721);
  FullAdder U1254 (w4721, w4644, IN46[25], w4722, w4723);
  FullAdder U1255 (w4723, w4646, IN47[24], w4724, w4725);
  FullAdder U1256 (w4725, w4648, IN48[23], w4726, w4727);
  FullAdder U1257 (w4727, w4650, IN49[22], w4728, w4729);
  FullAdder U1258 (w4729, w4652, IN50[21], w4730, w4731);
  FullAdder U1259 (w4731, w4654, IN51[20], w4732, w4733);
  FullAdder U1260 (w4733, w4656, IN52[19], w4734, w4735);
  FullAdder U1261 (w4735, w4658, IN53[18], w4736, w4737);
  FullAdder U1262 (w4737, w4660, IN54[17], w4738, w4739);
  FullAdder U1263 (w4739, w4662, IN55[16], w4740, w4741);
  FullAdder U1264 (w4741, w4664, IN56[15], w4742, w4743);
  FullAdder U1265 (w4743, w4666, IN57[14], w4744, w4745);
  FullAdder U1266 (w4745, w4668, IN58[13], w4746, w4747);
  FullAdder U1267 (w4747, w4670, IN59[12], w4748, w4749);
  FullAdder U1268 (w4749, w4672, IN60[11], w4750, w4751);
  FullAdder U1269 (w4751, w4674, IN61[10], w4752, w4753);
  FullAdder U1270 (w4753, w4676, IN62[9], w4754, w4755);
  FullAdder U1271 (w4755, w4678, IN63[8], w4756, w4757);
  FullAdder U1272 (w4757, w4680, IN64[7], w4758, w4759);
  FullAdder U1273 (w4759, w4682, IN65[6], w4760, w4761);
  FullAdder U1274 (w4761, w4684, IN66[5], w4762, w4763);
  FullAdder U1275 (w4763, w4686, IN67[4], w4764, w4765);
  FullAdder U1276 (w4765, w4688, IN68[3], w4766, w4767);
  FullAdder U1277 (w4767, w4690, IN69[2], w4768, w4769);
  FullAdder U1278 (w4769, w4692, IN70[1], w4770, w4771);
  FullAdder U1279 (w4771, w4693, IN71[0], w4772, w4773);
  HalfAdder U1280 (w4696, IN33[33], Out1[33], w4775);
  FullAdder U1281 (w4775, w4698, IN34[33], w4776, w4777);
  FullAdder U1282 (w4777, w4700, IN35[33], w4778, w4779);
  FullAdder U1283 (w4779, w4702, IN36[33], w4780, w4781);
  FullAdder U1284 (w4781, w4704, IN37[33], w4782, w4783);
  FullAdder U1285 (w4783, w4706, IN38[33], w4784, w4785);
  FullAdder U1286 (w4785, w4708, IN39[33], w4786, w4787);
  FullAdder U1287 (w4787, w4710, IN40[33], w4788, w4789);
  FullAdder U1288 (w4789, w4712, IN41[31], w4790, w4791);
  FullAdder U1289 (w4791, w4714, IN42[30], w4792, w4793);
  FullAdder U1290 (w4793, w4716, IN43[29], w4794, w4795);
  FullAdder U1291 (w4795, w4718, IN44[28], w4796, w4797);
  FullAdder U1292 (w4797, w4720, IN45[27], w4798, w4799);
  FullAdder U1293 (w4799, w4722, IN46[26], w4800, w4801);
  FullAdder U1294 (w4801, w4724, IN47[25], w4802, w4803);
  FullAdder U1295 (w4803, w4726, IN48[24], w4804, w4805);
  FullAdder U1296 (w4805, w4728, IN49[23], w4806, w4807);
  FullAdder U1297 (w4807, w4730, IN50[22], w4808, w4809);
  FullAdder U1298 (w4809, w4732, IN51[21], w4810, w4811);
  FullAdder U1299 (w4811, w4734, IN52[20], w4812, w4813);
  FullAdder U1300 (w4813, w4736, IN53[19], w4814, w4815);
  FullAdder U1301 (w4815, w4738, IN54[18], w4816, w4817);
  FullAdder U1302 (w4817, w4740, IN55[17], w4818, w4819);
  FullAdder U1303 (w4819, w4742, IN56[16], w4820, w4821);
  FullAdder U1304 (w4821, w4744, IN57[15], w4822, w4823);
  FullAdder U1305 (w4823, w4746, IN58[14], w4824, w4825);
  FullAdder U1306 (w4825, w4748, IN59[13], w4826, w4827);
  FullAdder U1307 (w4827, w4750, IN60[12], w4828, w4829);
  FullAdder U1308 (w4829, w4752, IN61[11], w4830, w4831);
  FullAdder U1309 (w4831, w4754, IN62[10], w4832, w4833);
  FullAdder U1310 (w4833, w4756, IN63[9], w4834, w4835);
  FullAdder U1311 (w4835, w4758, IN64[8], w4836, w4837);
  FullAdder U1312 (w4837, w4760, IN65[7], w4838, w4839);
  FullAdder U1313 (w4839, w4762, IN66[6], w4840, w4841);
  FullAdder U1314 (w4841, w4764, IN67[5], w4842, w4843);
  FullAdder U1315 (w4843, w4766, IN68[4], w4844, w4845);
  FullAdder U1316 (w4845, w4768, IN69[3], w4846, w4847);
  FullAdder U1317 (w4847, w4770, IN70[2], w4848, w4849);
  FullAdder U1318 (w4849, w4772, IN71[1], w4850, w4851);
  FullAdder U1319 (w4851, w4773, IN72[0], w4852, w4853);
  HalfAdder U1320 (w4776, IN34[34], Out1[34], w4855);
  FullAdder U1321 (w4855, w4778, IN35[34], w4856, w4857);
  FullAdder U1322 (w4857, w4780, IN36[34], w4858, w4859);
  FullAdder U1323 (w4859, w4782, IN37[34], w4860, w4861);
  FullAdder U1324 (w4861, w4784, IN38[34], w4862, w4863);
  FullAdder U1325 (w4863, w4786, IN39[34], w4864, w4865);
  FullAdder U1326 (w4865, w4788, IN40[34], w4866, w4867);
  FullAdder U1327 (w4867, w4790, IN41[32], w4868, w4869);
  FullAdder U1328 (w4869, w4792, IN42[31], w4870, w4871);
  FullAdder U1329 (w4871, w4794, IN43[30], w4872, w4873);
  FullAdder U1330 (w4873, w4796, IN44[29], w4874, w4875);
  FullAdder U1331 (w4875, w4798, IN45[28], w4876, w4877);
  FullAdder U1332 (w4877, w4800, IN46[27], w4878, w4879);
  FullAdder U1333 (w4879, w4802, IN47[26], w4880, w4881);
  FullAdder U1334 (w4881, w4804, IN48[25], w4882, w4883);
  FullAdder U1335 (w4883, w4806, IN49[24], w4884, w4885);
  FullAdder U1336 (w4885, w4808, IN50[23], w4886, w4887);
  FullAdder U1337 (w4887, w4810, IN51[22], w4888, w4889);
  FullAdder U1338 (w4889, w4812, IN52[21], w4890, w4891);
  FullAdder U1339 (w4891, w4814, IN53[20], w4892, w4893);
  FullAdder U1340 (w4893, w4816, IN54[19], w4894, w4895);
  FullAdder U1341 (w4895, w4818, IN55[18], w4896, w4897);
  FullAdder U1342 (w4897, w4820, IN56[17], w4898, w4899);
  FullAdder U1343 (w4899, w4822, IN57[16], w4900, w4901);
  FullAdder U1344 (w4901, w4824, IN58[15], w4902, w4903);
  FullAdder U1345 (w4903, w4826, IN59[14], w4904, w4905);
  FullAdder U1346 (w4905, w4828, IN60[13], w4906, w4907);
  FullAdder U1347 (w4907, w4830, IN61[12], w4908, w4909);
  FullAdder U1348 (w4909, w4832, IN62[11], w4910, w4911);
  FullAdder U1349 (w4911, w4834, IN63[10], w4912, w4913);
  FullAdder U1350 (w4913, w4836, IN64[9], w4914, w4915);
  FullAdder U1351 (w4915, w4838, IN65[8], w4916, w4917);
  FullAdder U1352 (w4917, w4840, IN66[7], w4918, w4919);
  FullAdder U1353 (w4919, w4842, IN67[6], w4920, w4921);
  FullAdder U1354 (w4921, w4844, IN68[5], w4922, w4923);
  FullAdder U1355 (w4923, w4846, IN69[4], w4924, w4925);
  FullAdder U1356 (w4925, w4848, IN70[3], w4926, w4927);
  FullAdder U1357 (w4927, w4850, IN71[2], w4928, w4929);
  FullAdder U1358 (w4929, w4852, IN72[1], w4930, w4931);
  FullAdder U1359 (w4931, w4853, IN73[0], w4932, w4933);
  HalfAdder U1360 (w4856, IN35[35], Out1[35], w4935);
  FullAdder U1361 (w4935, w4858, IN36[35], w4936, w4937);
  FullAdder U1362 (w4937, w4860, IN37[35], w4938, w4939);
  FullAdder U1363 (w4939, w4862, IN38[35], w4940, w4941);
  FullAdder U1364 (w4941, w4864, IN39[35], w4942, w4943);
  FullAdder U1365 (w4943, w4866, IN40[35], w4944, w4945);
  FullAdder U1366 (w4945, w4868, IN41[33], w4946, w4947);
  FullAdder U1367 (w4947, w4870, IN42[32], w4948, w4949);
  FullAdder U1368 (w4949, w4872, IN43[31], w4950, w4951);
  FullAdder U1369 (w4951, w4874, IN44[30], w4952, w4953);
  FullAdder U1370 (w4953, w4876, IN45[29], w4954, w4955);
  FullAdder U1371 (w4955, w4878, IN46[28], w4956, w4957);
  FullAdder U1372 (w4957, w4880, IN47[27], w4958, w4959);
  FullAdder U1373 (w4959, w4882, IN48[26], w4960, w4961);
  FullAdder U1374 (w4961, w4884, IN49[25], w4962, w4963);
  FullAdder U1375 (w4963, w4886, IN50[24], w4964, w4965);
  FullAdder U1376 (w4965, w4888, IN51[23], w4966, w4967);
  FullAdder U1377 (w4967, w4890, IN52[22], w4968, w4969);
  FullAdder U1378 (w4969, w4892, IN53[21], w4970, w4971);
  FullAdder U1379 (w4971, w4894, IN54[20], w4972, w4973);
  FullAdder U1380 (w4973, w4896, IN55[19], w4974, w4975);
  FullAdder U1381 (w4975, w4898, IN56[18], w4976, w4977);
  FullAdder U1382 (w4977, w4900, IN57[17], w4978, w4979);
  FullAdder U1383 (w4979, w4902, IN58[16], w4980, w4981);
  FullAdder U1384 (w4981, w4904, IN59[15], w4982, w4983);
  FullAdder U1385 (w4983, w4906, IN60[14], w4984, w4985);
  FullAdder U1386 (w4985, w4908, IN61[13], w4986, w4987);
  FullAdder U1387 (w4987, w4910, IN62[12], w4988, w4989);
  FullAdder U1388 (w4989, w4912, IN63[11], w4990, w4991);
  FullAdder U1389 (w4991, w4914, IN64[10], w4992, w4993);
  FullAdder U1390 (w4993, w4916, IN65[9], w4994, w4995);
  FullAdder U1391 (w4995, w4918, IN66[8], w4996, w4997);
  FullAdder U1392 (w4997, w4920, IN67[7], w4998, w4999);
  FullAdder U1393 (w4999, w4922, IN68[6], w5000, w5001);
  FullAdder U1394 (w5001, w4924, IN69[5], w5002, w5003);
  FullAdder U1395 (w5003, w4926, IN70[4], w5004, w5005);
  FullAdder U1396 (w5005, w4928, IN71[3], w5006, w5007);
  FullAdder U1397 (w5007, w4930, IN72[2], w5008, w5009);
  FullAdder U1398 (w5009, w4932, IN73[1], w5010, w5011);
  FullAdder U1399 (w5011, w4933, IN74[0], w5012, w5013);
  HalfAdder U1400 (w4936, IN36[36], Out1[36], w5015);
  FullAdder U1401 (w5015, w4938, IN37[36], w5016, w5017);
  FullAdder U1402 (w5017, w4940, IN38[36], w5018, w5019);
  FullAdder U1403 (w5019, w4942, IN39[36], w5020, w5021);
  FullAdder U1404 (w5021, w4944, IN40[36], w5022, w5023);
  FullAdder U1405 (w5023, w4946, IN41[34], w5024, w5025);
  FullAdder U1406 (w5025, w4948, IN42[33], w5026, w5027);
  FullAdder U1407 (w5027, w4950, IN43[32], w5028, w5029);
  FullAdder U1408 (w5029, w4952, IN44[31], w5030, w5031);
  FullAdder U1409 (w5031, w4954, IN45[30], w5032, w5033);
  FullAdder U1410 (w5033, w4956, IN46[29], w5034, w5035);
  FullAdder U1411 (w5035, w4958, IN47[28], w5036, w5037);
  FullAdder U1412 (w5037, w4960, IN48[27], w5038, w5039);
  FullAdder U1413 (w5039, w4962, IN49[26], w5040, w5041);
  FullAdder U1414 (w5041, w4964, IN50[25], w5042, w5043);
  FullAdder U1415 (w5043, w4966, IN51[24], w5044, w5045);
  FullAdder U1416 (w5045, w4968, IN52[23], w5046, w5047);
  FullAdder U1417 (w5047, w4970, IN53[22], w5048, w5049);
  FullAdder U1418 (w5049, w4972, IN54[21], w5050, w5051);
  FullAdder U1419 (w5051, w4974, IN55[20], w5052, w5053);
  FullAdder U1420 (w5053, w4976, IN56[19], w5054, w5055);
  FullAdder U1421 (w5055, w4978, IN57[18], w5056, w5057);
  FullAdder U1422 (w5057, w4980, IN58[17], w5058, w5059);
  FullAdder U1423 (w5059, w4982, IN59[16], w5060, w5061);
  FullAdder U1424 (w5061, w4984, IN60[15], w5062, w5063);
  FullAdder U1425 (w5063, w4986, IN61[14], w5064, w5065);
  FullAdder U1426 (w5065, w4988, IN62[13], w5066, w5067);
  FullAdder U1427 (w5067, w4990, IN63[12], w5068, w5069);
  FullAdder U1428 (w5069, w4992, IN64[11], w5070, w5071);
  FullAdder U1429 (w5071, w4994, IN65[10], w5072, w5073);
  FullAdder U1430 (w5073, w4996, IN66[9], w5074, w5075);
  FullAdder U1431 (w5075, w4998, IN67[8], w5076, w5077);
  FullAdder U1432 (w5077, w5000, IN68[7], w5078, w5079);
  FullAdder U1433 (w5079, w5002, IN69[6], w5080, w5081);
  FullAdder U1434 (w5081, w5004, IN70[5], w5082, w5083);
  FullAdder U1435 (w5083, w5006, IN71[4], w5084, w5085);
  FullAdder U1436 (w5085, w5008, IN72[3], w5086, w5087);
  FullAdder U1437 (w5087, w5010, IN73[2], w5088, w5089);
  FullAdder U1438 (w5089, w5012, IN74[1], w5090, w5091);
  FullAdder U1439 (w5091, w5013, IN75[0], w5092, w5093);
  HalfAdder U1440 (w5016, IN37[37], Out1[37], w5095);
  FullAdder U1441 (w5095, w5018, IN38[37], w5096, w5097);
  FullAdder U1442 (w5097, w5020, IN39[37], w5098, w5099);
  FullAdder U1443 (w5099, w5022, IN40[37], w5100, w5101);
  FullAdder U1444 (w5101, w5024, IN41[35], w5102, w5103);
  FullAdder U1445 (w5103, w5026, IN42[34], w5104, w5105);
  FullAdder U1446 (w5105, w5028, IN43[33], w5106, w5107);
  FullAdder U1447 (w5107, w5030, IN44[32], w5108, w5109);
  FullAdder U1448 (w5109, w5032, IN45[31], w5110, w5111);
  FullAdder U1449 (w5111, w5034, IN46[30], w5112, w5113);
  FullAdder U1450 (w5113, w5036, IN47[29], w5114, w5115);
  FullAdder U1451 (w5115, w5038, IN48[28], w5116, w5117);
  FullAdder U1452 (w5117, w5040, IN49[27], w5118, w5119);
  FullAdder U1453 (w5119, w5042, IN50[26], w5120, w5121);
  FullAdder U1454 (w5121, w5044, IN51[25], w5122, w5123);
  FullAdder U1455 (w5123, w5046, IN52[24], w5124, w5125);
  FullAdder U1456 (w5125, w5048, IN53[23], w5126, w5127);
  FullAdder U1457 (w5127, w5050, IN54[22], w5128, w5129);
  FullAdder U1458 (w5129, w5052, IN55[21], w5130, w5131);
  FullAdder U1459 (w5131, w5054, IN56[20], w5132, w5133);
  FullAdder U1460 (w5133, w5056, IN57[19], w5134, w5135);
  FullAdder U1461 (w5135, w5058, IN58[18], w5136, w5137);
  FullAdder U1462 (w5137, w5060, IN59[17], w5138, w5139);
  FullAdder U1463 (w5139, w5062, IN60[16], w5140, w5141);
  FullAdder U1464 (w5141, w5064, IN61[15], w5142, w5143);
  FullAdder U1465 (w5143, w5066, IN62[14], w5144, w5145);
  FullAdder U1466 (w5145, w5068, IN63[13], w5146, w5147);
  FullAdder U1467 (w5147, w5070, IN64[12], w5148, w5149);
  FullAdder U1468 (w5149, w5072, IN65[11], w5150, w5151);
  FullAdder U1469 (w5151, w5074, IN66[10], w5152, w5153);
  FullAdder U1470 (w5153, w5076, IN67[9], w5154, w5155);
  FullAdder U1471 (w5155, w5078, IN68[8], w5156, w5157);
  FullAdder U1472 (w5157, w5080, IN69[7], w5158, w5159);
  FullAdder U1473 (w5159, w5082, IN70[6], w5160, w5161);
  FullAdder U1474 (w5161, w5084, IN71[5], w5162, w5163);
  FullAdder U1475 (w5163, w5086, IN72[4], w5164, w5165);
  FullAdder U1476 (w5165, w5088, IN73[3], w5166, w5167);
  FullAdder U1477 (w5167, w5090, IN74[2], w5168, w5169);
  FullAdder U1478 (w5169, w5092, IN75[1], w5170, w5171);
  FullAdder U1479 (w5171, w5093, IN76[0], w5172, w5173);
  HalfAdder U1480 (w5096, IN38[38], Out1[38], w5175);
  FullAdder U1481 (w5175, w5098, IN39[38], w5176, w5177);
  FullAdder U1482 (w5177, w5100, IN40[38], w5178, w5179);
  FullAdder U1483 (w5179, w5102, IN41[36], w5180, w5181);
  FullAdder U1484 (w5181, w5104, IN42[35], w5182, w5183);
  FullAdder U1485 (w5183, w5106, IN43[34], w5184, w5185);
  FullAdder U1486 (w5185, w5108, IN44[33], w5186, w5187);
  FullAdder U1487 (w5187, w5110, IN45[32], w5188, w5189);
  FullAdder U1488 (w5189, w5112, IN46[31], w5190, w5191);
  FullAdder U1489 (w5191, w5114, IN47[30], w5192, w5193);
  FullAdder U1490 (w5193, w5116, IN48[29], w5194, w5195);
  FullAdder U1491 (w5195, w5118, IN49[28], w5196, w5197);
  FullAdder U1492 (w5197, w5120, IN50[27], w5198, w5199);
  FullAdder U1493 (w5199, w5122, IN51[26], w5200, w5201);
  FullAdder U1494 (w5201, w5124, IN52[25], w5202, w5203);
  FullAdder U1495 (w5203, w5126, IN53[24], w5204, w5205);
  FullAdder U1496 (w5205, w5128, IN54[23], w5206, w5207);
  FullAdder U1497 (w5207, w5130, IN55[22], w5208, w5209);
  FullAdder U1498 (w5209, w5132, IN56[21], w5210, w5211);
  FullAdder U1499 (w5211, w5134, IN57[20], w5212, w5213);
  FullAdder U1500 (w5213, w5136, IN58[19], w5214, w5215);
  FullAdder U1501 (w5215, w5138, IN59[18], w5216, w5217);
  FullAdder U1502 (w5217, w5140, IN60[17], w5218, w5219);
  FullAdder U1503 (w5219, w5142, IN61[16], w5220, w5221);
  FullAdder U1504 (w5221, w5144, IN62[15], w5222, w5223);
  FullAdder U1505 (w5223, w5146, IN63[14], w5224, w5225);
  FullAdder U1506 (w5225, w5148, IN64[13], w5226, w5227);
  FullAdder U1507 (w5227, w5150, IN65[12], w5228, w5229);
  FullAdder U1508 (w5229, w5152, IN66[11], w5230, w5231);
  FullAdder U1509 (w5231, w5154, IN67[10], w5232, w5233);
  FullAdder U1510 (w5233, w5156, IN68[9], w5234, w5235);
  FullAdder U1511 (w5235, w5158, IN69[8], w5236, w5237);
  FullAdder U1512 (w5237, w5160, IN70[7], w5238, w5239);
  FullAdder U1513 (w5239, w5162, IN71[6], w5240, w5241);
  FullAdder U1514 (w5241, w5164, IN72[5], w5242, w5243);
  FullAdder U1515 (w5243, w5166, IN73[4], w5244, w5245);
  FullAdder U1516 (w5245, w5168, IN74[3], w5246, w5247);
  FullAdder U1517 (w5247, w5170, IN75[2], w5248, w5249);
  FullAdder U1518 (w5249, w5172, IN76[1], w5250, w5251);
  FullAdder U1519 (w5251, w5173, IN77[0], w5252, w5253);
  HalfAdder U1520 (w5176, IN39[39], Out1[39], w5255);
  FullAdder U1521 (w5255, w5178, IN40[39], w5256, w5257);
  FullAdder U1522 (w5257, w5180, IN41[37], w5258, w5259);
  FullAdder U1523 (w5259, w5182, IN42[36], w5260, w5261);
  FullAdder U1524 (w5261, w5184, IN43[35], w5262, w5263);
  FullAdder U1525 (w5263, w5186, IN44[34], w5264, w5265);
  FullAdder U1526 (w5265, w5188, IN45[33], w5266, w5267);
  FullAdder U1527 (w5267, w5190, IN46[32], w5268, w5269);
  FullAdder U1528 (w5269, w5192, IN47[31], w5270, w5271);
  FullAdder U1529 (w5271, w5194, IN48[30], w5272, w5273);
  FullAdder U1530 (w5273, w5196, IN49[29], w5274, w5275);
  FullAdder U1531 (w5275, w5198, IN50[28], w5276, w5277);
  FullAdder U1532 (w5277, w5200, IN51[27], w5278, w5279);
  FullAdder U1533 (w5279, w5202, IN52[26], w5280, w5281);
  FullAdder U1534 (w5281, w5204, IN53[25], w5282, w5283);
  FullAdder U1535 (w5283, w5206, IN54[24], w5284, w5285);
  FullAdder U1536 (w5285, w5208, IN55[23], w5286, w5287);
  FullAdder U1537 (w5287, w5210, IN56[22], w5288, w5289);
  FullAdder U1538 (w5289, w5212, IN57[21], w5290, w5291);
  FullAdder U1539 (w5291, w5214, IN58[20], w5292, w5293);
  FullAdder U1540 (w5293, w5216, IN59[19], w5294, w5295);
  FullAdder U1541 (w5295, w5218, IN60[18], w5296, w5297);
  FullAdder U1542 (w5297, w5220, IN61[17], w5298, w5299);
  FullAdder U1543 (w5299, w5222, IN62[16], w5300, w5301);
  FullAdder U1544 (w5301, w5224, IN63[15], w5302, w5303);
  FullAdder U1545 (w5303, w5226, IN64[14], w5304, w5305);
  FullAdder U1546 (w5305, w5228, IN65[13], w5306, w5307);
  FullAdder U1547 (w5307, w5230, IN66[12], w5308, w5309);
  FullAdder U1548 (w5309, w5232, IN67[11], w5310, w5311);
  FullAdder U1549 (w5311, w5234, IN68[10], w5312, w5313);
  FullAdder U1550 (w5313, w5236, IN69[9], w5314, w5315);
  FullAdder U1551 (w5315, w5238, IN70[8], w5316, w5317);
  FullAdder U1552 (w5317, w5240, IN71[7], w5318, w5319);
  FullAdder U1553 (w5319, w5242, IN72[6], w5320, w5321);
  FullAdder U1554 (w5321, w5244, IN73[5], w5322, w5323);
  FullAdder U1555 (w5323, w5246, IN74[4], w5324, w5325);
  FullAdder U1556 (w5325, w5248, IN75[3], w5326, w5327);
  FullAdder U1557 (w5327, w5250, IN76[2], w5328, w5329);
  FullAdder U1558 (w5329, w5252, IN77[1], w5330, w5331);
  FullAdder U1559 (w5331, w5253, IN78[0], w5332, w5333);
  HalfAdder U1560 (w5256, IN40[40], Out1[40], w5335);
  FullAdder U1561 (w5335, w5258, IN41[38], w5336, w5337);
  FullAdder U1562 (w5337, w5260, IN42[37], w5338, w5339);
  FullAdder U1563 (w5339, w5262, IN43[36], w5340, w5341);
  FullAdder U1564 (w5341, w5264, IN44[35], w5342, w5343);
  FullAdder U1565 (w5343, w5266, IN45[34], w5344, w5345);
  FullAdder U1566 (w5345, w5268, IN46[33], w5346, w5347);
  FullAdder U1567 (w5347, w5270, IN47[32], w5348, w5349);
  FullAdder U1568 (w5349, w5272, IN48[31], w5350, w5351);
  FullAdder U1569 (w5351, w5274, IN49[30], w5352, w5353);
  FullAdder U1570 (w5353, w5276, IN50[29], w5354, w5355);
  FullAdder U1571 (w5355, w5278, IN51[28], w5356, w5357);
  FullAdder U1572 (w5357, w5280, IN52[27], w5358, w5359);
  FullAdder U1573 (w5359, w5282, IN53[26], w5360, w5361);
  FullAdder U1574 (w5361, w5284, IN54[25], w5362, w5363);
  FullAdder U1575 (w5363, w5286, IN55[24], w5364, w5365);
  FullAdder U1576 (w5365, w5288, IN56[23], w5366, w5367);
  FullAdder U1577 (w5367, w5290, IN57[22], w5368, w5369);
  FullAdder U1578 (w5369, w5292, IN58[21], w5370, w5371);
  FullAdder U1579 (w5371, w5294, IN59[20], w5372, w5373);
  FullAdder U1580 (w5373, w5296, IN60[19], w5374, w5375);
  FullAdder U1581 (w5375, w5298, IN61[18], w5376, w5377);
  FullAdder U1582 (w5377, w5300, IN62[17], w5378, w5379);
  FullAdder U1583 (w5379, w5302, IN63[16], w5380, w5381);
  FullAdder U1584 (w5381, w5304, IN64[15], w5382, w5383);
  FullAdder U1585 (w5383, w5306, IN65[14], w5384, w5385);
  FullAdder U1586 (w5385, w5308, IN66[13], w5386, w5387);
  FullAdder U1587 (w5387, w5310, IN67[12], w5388, w5389);
  FullAdder U1588 (w5389, w5312, IN68[11], w5390, w5391);
  FullAdder U1589 (w5391, w5314, IN69[10], w5392, w5393);
  FullAdder U1590 (w5393, w5316, IN70[9], w5394, w5395);
  FullAdder U1591 (w5395, w5318, IN71[8], w5396, w5397);
  FullAdder U1592 (w5397, w5320, IN72[7], w5398, w5399);
  FullAdder U1593 (w5399, w5322, IN73[6], w5400, w5401);
  FullAdder U1594 (w5401, w5324, IN74[5], w5402, w5403);
  FullAdder U1595 (w5403, w5326, IN75[4], w5404, w5405);
  FullAdder U1596 (w5405, w5328, IN76[3], w5406, w5407);
  FullAdder U1597 (w5407, w5330, IN77[2], w5408, w5409);
  FullAdder U1598 (w5409, w5332, IN78[1], w5410, w5411);
  FullAdder U1599 (w5411, w5333, IN79[0], w5412, w5413);
  HalfAdder U1600 (w5336, IN41[39], Out1[41], w5415);
  FullAdder U1601 (w5415, w5338, IN42[38], w5416, w5417);
  FullAdder U1602 (w5417, w5340, IN43[37], w5418, w5419);
  FullAdder U1603 (w5419, w5342, IN44[36], w5420, w5421);
  FullAdder U1604 (w5421, w5344, IN45[35], w5422, w5423);
  FullAdder U1605 (w5423, w5346, IN46[34], w5424, w5425);
  FullAdder U1606 (w5425, w5348, IN47[33], w5426, w5427);
  FullAdder U1607 (w5427, w5350, IN48[32], w5428, w5429);
  FullAdder U1608 (w5429, w5352, IN49[31], w5430, w5431);
  FullAdder U1609 (w5431, w5354, IN50[30], w5432, w5433);
  FullAdder U1610 (w5433, w5356, IN51[29], w5434, w5435);
  FullAdder U1611 (w5435, w5358, IN52[28], w5436, w5437);
  FullAdder U1612 (w5437, w5360, IN53[27], w5438, w5439);
  FullAdder U1613 (w5439, w5362, IN54[26], w5440, w5441);
  FullAdder U1614 (w5441, w5364, IN55[25], w5442, w5443);
  FullAdder U1615 (w5443, w5366, IN56[24], w5444, w5445);
  FullAdder U1616 (w5445, w5368, IN57[23], w5446, w5447);
  FullAdder U1617 (w5447, w5370, IN58[22], w5448, w5449);
  FullAdder U1618 (w5449, w5372, IN59[21], w5450, w5451);
  FullAdder U1619 (w5451, w5374, IN60[20], w5452, w5453);
  FullAdder U1620 (w5453, w5376, IN61[19], w5454, w5455);
  FullAdder U1621 (w5455, w5378, IN62[18], w5456, w5457);
  FullAdder U1622 (w5457, w5380, IN63[17], w5458, w5459);
  FullAdder U1623 (w5459, w5382, IN64[16], w5460, w5461);
  FullAdder U1624 (w5461, w5384, IN65[15], w5462, w5463);
  FullAdder U1625 (w5463, w5386, IN66[14], w5464, w5465);
  FullAdder U1626 (w5465, w5388, IN67[13], w5466, w5467);
  FullAdder U1627 (w5467, w5390, IN68[12], w5468, w5469);
  FullAdder U1628 (w5469, w5392, IN69[11], w5470, w5471);
  FullAdder U1629 (w5471, w5394, IN70[10], w5472, w5473);
  FullAdder U1630 (w5473, w5396, IN71[9], w5474, w5475);
  FullAdder U1631 (w5475, w5398, IN72[8], w5476, w5477);
  FullAdder U1632 (w5477, w5400, IN73[7], w5478, w5479);
  FullAdder U1633 (w5479, w5402, IN74[6], w5480, w5481);
  FullAdder U1634 (w5481, w5404, IN75[5], w5482, w5483);
  FullAdder U1635 (w5483, w5406, IN76[4], w5484, w5485);
  FullAdder U1636 (w5485, w5408, IN77[3], w5486, w5487);
  FullAdder U1637 (w5487, w5410, IN78[2], w5488, w5489);
  FullAdder U1638 (w5489, w5412, IN79[1], w5490, w5491);
  FullAdder U1639 (w5491, w5413, IN80[0], w5492, w5493);
  HalfAdder U1640 (w5416, IN42[39], Out1[42], w5495);
  FullAdder U1641 (w5495, w5418, IN43[38], w5496, w5497);
  FullAdder U1642 (w5497, w5420, IN44[37], w5498, w5499);
  FullAdder U1643 (w5499, w5422, IN45[36], w5500, w5501);
  FullAdder U1644 (w5501, w5424, IN46[35], w5502, w5503);
  FullAdder U1645 (w5503, w5426, IN47[34], w5504, w5505);
  FullAdder U1646 (w5505, w5428, IN48[33], w5506, w5507);
  FullAdder U1647 (w5507, w5430, IN49[32], w5508, w5509);
  FullAdder U1648 (w5509, w5432, IN50[31], w5510, w5511);
  FullAdder U1649 (w5511, w5434, IN51[30], w5512, w5513);
  FullAdder U1650 (w5513, w5436, IN52[29], w5514, w5515);
  FullAdder U1651 (w5515, w5438, IN53[28], w5516, w5517);
  FullAdder U1652 (w5517, w5440, IN54[27], w5518, w5519);
  FullAdder U1653 (w5519, w5442, IN55[26], w5520, w5521);
  FullAdder U1654 (w5521, w5444, IN56[25], w5522, w5523);
  FullAdder U1655 (w5523, w5446, IN57[24], w5524, w5525);
  FullAdder U1656 (w5525, w5448, IN58[23], w5526, w5527);
  FullAdder U1657 (w5527, w5450, IN59[22], w5528, w5529);
  FullAdder U1658 (w5529, w5452, IN60[21], w5530, w5531);
  FullAdder U1659 (w5531, w5454, IN61[20], w5532, w5533);
  FullAdder U1660 (w5533, w5456, IN62[19], w5534, w5535);
  FullAdder U1661 (w5535, w5458, IN63[18], w5536, w5537);
  FullAdder U1662 (w5537, w5460, IN64[17], w5538, w5539);
  FullAdder U1663 (w5539, w5462, IN65[16], w5540, w5541);
  FullAdder U1664 (w5541, w5464, IN66[15], w5542, w5543);
  FullAdder U1665 (w5543, w5466, IN67[14], w5544, w5545);
  FullAdder U1666 (w5545, w5468, IN68[13], w5546, w5547);
  FullAdder U1667 (w5547, w5470, IN69[12], w5548, w5549);
  FullAdder U1668 (w5549, w5472, IN70[11], w5550, w5551);
  FullAdder U1669 (w5551, w5474, IN71[10], w5552, w5553);
  FullAdder U1670 (w5553, w5476, IN72[9], w5554, w5555);
  FullAdder U1671 (w5555, w5478, IN73[8], w5556, w5557);
  FullAdder U1672 (w5557, w5480, IN74[7], w5558, w5559);
  FullAdder U1673 (w5559, w5482, IN75[6], w5560, w5561);
  FullAdder U1674 (w5561, w5484, IN76[5], w5562, w5563);
  FullAdder U1675 (w5563, w5486, IN77[4], w5564, w5565);
  FullAdder U1676 (w5565, w5488, IN78[3], w5566, w5567);
  FullAdder U1677 (w5567, w5490, IN79[2], w5568, w5569);
  FullAdder U1678 (w5569, w5492, IN80[1], w5570, w5571);
  FullAdder U1679 (w5571, w5493, IN81[0], w5572, w5573);
  HalfAdder U1680 (w5496, IN43[39], Out1[43], w5575);
  FullAdder U1681 (w5575, w5498, IN44[38], w5576, w5577);
  FullAdder U1682 (w5577, w5500, IN45[37], w5578, w5579);
  FullAdder U1683 (w5579, w5502, IN46[36], w5580, w5581);
  FullAdder U1684 (w5581, w5504, IN47[35], w5582, w5583);
  FullAdder U1685 (w5583, w5506, IN48[34], w5584, w5585);
  FullAdder U1686 (w5585, w5508, IN49[33], w5586, w5587);
  FullAdder U1687 (w5587, w5510, IN50[32], w5588, w5589);
  FullAdder U1688 (w5589, w5512, IN51[31], w5590, w5591);
  FullAdder U1689 (w5591, w5514, IN52[30], w5592, w5593);
  FullAdder U1690 (w5593, w5516, IN53[29], w5594, w5595);
  FullAdder U1691 (w5595, w5518, IN54[28], w5596, w5597);
  FullAdder U1692 (w5597, w5520, IN55[27], w5598, w5599);
  FullAdder U1693 (w5599, w5522, IN56[26], w5600, w5601);
  FullAdder U1694 (w5601, w5524, IN57[25], w5602, w5603);
  FullAdder U1695 (w5603, w5526, IN58[24], w5604, w5605);
  FullAdder U1696 (w5605, w5528, IN59[23], w5606, w5607);
  FullAdder U1697 (w5607, w5530, IN60[22], w5608, w5609);
  FullAdder U1698 (w5609, w5532, IN61[21], w5610, w5611);
  FullAdder U1699 (w5611, w5534, IN62[20], w5612, w5613);
  FullAdder U1700 (w5613, w5536, IN63[19], w5614, w5615);
  FullAdder U1701 (w5615, w5538, IN64[18], w5616, w5617);
  FullAdder U1702 (w5617, w5540, IN65[17], w5618, w5619);
  FullAdder U1703 (w5619, w5542, IN66[16], w5620, w5621);
  FullAdder U1704 (w5621, w5544, IN67[15], w5622, w5623);
  FullAdder U1705 (w5623, w5546, IN68[14], w5624, w5625);
  FullAdder U1706 (w5625, w5548, IN69[13], w5626, w5627);
  FullAdder U1707 (w5627, w5550, IN70[12], w5628, w5629);
  FullAdder U1708 (w5629, w5552, IN71[11], w5630, w5631);
  FullAdder U1709 (w5631, w5554, IN72[10], w5632, w5633);
  FullAdder U1710 (w5633, w5556, IN73[9], w5634, w5635);
  FullAdder U1711 (w5635, w5558, IN74[8], w5636, w5637);
  FullAdder U1712 (w5637, w5560, IN75[7], w5638, w5639);
  FullAdder U1713 (w5639, w5562, IN76[6], w5640, w5641);
  FullAdder U1714 (w5641, w5564, IN77[5], w5642, w5643);
  FullAdder U1715 (w5643, w5566, IN78[4], w5644, w5645);
  FullAdder U1716 (w5645, w5568, IN79[3], w5646, w5647);
  FullAdder U1717 (w5647, w5570, IN80[2], w5648, w5649);
  FullAdder U1718 (w5649, w5572, IN81[1], w5650, w5651);
  FullAdder U1719 (w5651, w5573, IN82[0], w5652, w5653);
  HalfAdder U1720 (w5576, IN44[39], Out1[44], w5655);
  FullAdder U1721 (w5655, w5578, IN45[38], w5656, w5657);
  FullAdder U1722 (w5657, w5580, IN46[37], w5658, w5659);
  FullAdder U1723 (w5659, w5582, IN47[36], w5660, w5661);
  FullAdder U1724 (w5661, w5584, IN48[35], w5662, w5663);
  FullAdder U1725 (w5663, w5586, IN49[34], w5664, w5665);
  FullAdder U1726 (w5665, w5588, IN50[33], w5666, w5667);
  FullAdder U1727 (w5667, w5590, IN51[32], w5668, w5669);
  FullAdder U1728 (w5669, w5592, IN52[31], w5670, w5671);
  FullAdder U1729 (w5671, w5594, IN53[30], w5672, w5673);
  FullAdder U1730 (w5673, w5596, IN54[29], w5674, w5675);
  FullAdder U1731 (w5675, w5598, IN55[28], w5676, w5677);
  FullAdder U1732 (w5677, w5600, IN56[27], w5678, w5679);
  FullAdder U1733 (w5679, w5602, IN57[26], w5680, w5681);
  FullAdder U1734 (w5681, w5604, IN58[25], w5682, w5683);
  FullAdder U1735 (w5683, w5606, IN59[24], w5684, w5685);
  FullAdder U1736 (w5685, w5608, IN60[23], w5686, w5687);
  FullAdder U1737 (w5687, w5610, IN61[22], w5688, w5689);
  FullAdder U1738 (w5689, w5612, IN62[21], w5690, w5691);
  FullAdder U1739 (w5691, w5614, IN63[20], w5692, w5693);
  FullAdder U1740 (w5693, w5616, IN64[19], w5694, w5695);
  FullAdder U1741 (w5695, w5618, IN65[18], w5696, w5697);
  FullAdder U1742 (w5697, w5620, IN66[17], w5698, w5699);
  FullAdder U1743 (w5699, w5622, IN67[16], w5700, w5701);
  FullAdder U1744 (w5701, w5624, IN68[15], w5702, w5703);
  FullAdder U1745 (w5703, w5626, IN69[14], w5704, w5705);
  FullAdder U1746 (w5705, w5628, IN70[13], w5706, w5707);
  FullAdder U1747 (w5707, w5630, IN71[12], w5708, w5709);
  FullAdder U1748 (w5709, w5632, IN72[11], w5710, w5711);
  FullAdder U1749 (w5711, w5634, IN73[10], w5712, w5713);
  FullAdder U1750 (w5713, w5636, IN74[9], w5714, w5715);
  FullAdder U1751 (w5715, w5638, IN75[8], w5716, w5717);
  FullAdder U1752 (w5717, w5640, IN76[7], w5718, w5719);
  FullAdder U1753 (w5719, w5642, IN77[6], w5720, w5721);
  FullAdder U1754 (w5721, w5644, IN78[5], w5722, w5723);
  FullAdder U1755 (w5723, w5646, IN79[4], w5724, w5725);
  FullAdder U1756 (w5725, w5648, IN80[3], w5726, w5727);
  FullAdder U1757 (w5727, w5650, IN81[2], w5728, w5729);
  FullAdder U1758 (w5729, w5652, IN82[1], w5730, w5731);
  FullAdder U1759 (w5731, w5653, IN83[0], w5732, w5733);
  HalfAdder U1760 (w5656, IN45[39], Out1[45], w5735);
  FullAdder U1761 (w5735, w5658, IN46[38], w5736, w5737);
  FullAdder U1762 (w5737, w5660, IN47[37], w5738, w5739);
  FullAdder U1763 (w5739, w5662, IN48[36], w5740, w5741);
  FullAdder U1764 (w5741, w5664, IN49[35], w5742, w5743);
  FullAdder U1765 (w5743, w5666, IN50[34], w5744, w5745);
  FullAdder U1766 (w5745, w5668, IN51[33], w5746, w5747);
  FullAdder U1767 (w5747, w5670, IN52[32], w5748, w5749);
  FullAdder U1768 (w5749, w5672, IN53[31], w5750, w5751);
  FullAdder U1769 (w5751, w5674, IN54[30], w5752, w5753);
  FullAdder U1770 (w5753, w5676, IN55[29], w5754, w5755);
  FullAdder U1771 (w5755, w5678, IN56[28], w5756, w5757);
  FullAdder U1772 (w5757, w5680, IN57[27], w5758, w5759);
  FullAdder U1773 (w5759, w5682, IN58[26], w5760, w5761);
  FullAdder U1774 (w5761, w5684, IN59[25], w5762, w5763);
  FullAdder U1775 (w5763, w5686, IN60[24], w5764, w5765);
  FullAdder U1776 (w5765, w5688, IN61[23], w5766, w5767);
  FullAdder U1777 (w5767, w5690, IN62[22], w5768, w5769);
  FullAdder U1778 (w5769, w5692, IN63[21], w5770, w5771);
  FullAdder U1779 (w5771, w5694, IN64[20], w5772, w5773);
  FullAdder U1780 (w5773, w5696, IN65[19], w5774, w5775);
  FullAdder U1781 (w5775, w5698, IN66[18], w5776, w5777);
  FullAdder U1782 (w5777, w5700, IN67[17], w5778, w5779);
  FullAdder U1783 (w5779, w5702, IN68[16], w5780, w5781);
  FullAdder U1784 (w5781, w5704, IN69[15], w5782, w5783);
  FullAdder U1785 (w5783, w5706, IN70[14], w5784, w5785);
  FullAdder U1786 (w5785, w5708, IN71[13], w5786, w5787);
  FullAdder U1787 (w5787, w5710, IN72[12], w5788, w5789);
  FullAdder U1788 (w5789, w5712, IN73[11], w5790, w5791);
  FullAdder U1789 (w5791, w5714, IN74[10], w5792, w5793);
  FullAdder U1790 (w5793, w5716, IN75[9], w5794, w5795);
  FullAdder U1791 (w5795, w5718, IN76[8], w5796, w5797);
  FullAdder U1792 (w5797, w5720, IN77[7], w5798, w5799);
  FullAdder U1793 (w5799, w5722, IN78[6], w5800, w5801);
  FullAdder U1794 (w5801, w5724, IN79[5], w5802, w5803);
  FullAdder U1795 (w5803, w5726, IN80[4], w5804, w5805);
  FullAdder U1796 (w5805, w5728, IN81[3], w5806, w5807);
  FullAdder U1797 (w5807, w5730, IN82[2], w5808, w5809);
  FullAdder U1798 (w5809, w5732, IN83[1], w5810, w5811);
  FullAdder U1799 (w5811, w5733, IN84[0], w5812, w5813);
  HalfAdder U1800 (w5736, IN46[39], Out1[46], w5815);
  FullAdder U1801 (w5815, w5738, IN47[38], w5816, w5817);
  FullAdder U1802 (w5817, w5740, IN48[37], w5818, w5819);
  FullAdder U1803 (w5819, w5742, IN49[36], w5820, w5821);
  FullAdder U1804 (w5821, w5744, IN50[35], w5822, w5823);
  FullAdder U1805 (w5823, w5746, IN51[34], w5824, w5825);
  FullAdder U1806 (w5825, w5748, IN52[33], w5826, w5827);
  FullAdder U1807 (w5827, w5750, IN53[32], w5828, w5829);
  FullAdder U1808 (w5829, w5752, IN54[31], w5830, w5831);
  FullAdder U1809 (w5831, w5754, IN55[30], w5832, w5833);
  FullAdder U1810 (w5833, w5756, IN56[29], w5834, w5835);
  FullAdder U1811 (w5835, w5758, IN57[28], w5836, w5837);
  FullAdder U1812 (w5837, w5760, IN58[27], w5838, w5839);
  FullAdder U1813 (w5839, w5762, IN59[26], w5840, w5841);
  FullAdder U1814 (w5841, w5764, IN60[25], w5842, w5843);
  FullAdder U1815 (w5843, w5766, IN61[24], w5844, w5845);
  FullAdder U1816 (w5845, w5768, IN62[23], w5846, w5847);
  FullAdder U1817 (w5847, w5770, IN63[22], w5848, w5849);
  FullAdder U1818 (w5849, w5772, IN64[21], w5850, w5851);
  FullAdder U1819 (w5851, w5774, IN65[20], w5852, w5853);
  FullAdder U1820 (w5853, w5776, IN66[19], w5854, w5855);
  FullAdder U1821 (w5855, w5778, IN67[18], w5856, w5857);
  FullAdder U1822 (w5857, w5780, IN68[17], w5858, w5859);
  FullAdder U1823 (w5859, w5782, IN69[16], w5860, w5861);
  FullAdder U1824 (w5861, w5784, IN70[15], w5862, w5863);
  FullAdder U1825 (w5863, w5786, IN71[14], w5864, w5865);
  FullAdder U1826 (w5865, w5788, IN72[13], w5866, w5867);
  FullAdder U1827 (w5867, w5790, IN73[12], w5868, w5869);
  FullAdder U1828 (w5869, w5792, IN74[11], w5870, w5871);
  FullAdder U1829 (w5871, w5794, IN75[10], w5872, w5873);
  FullAdder U1830 (w5873, w5796, IN76[9], w5874, w5875);
  FullAdder U1831 (w5875, w5798, IN77[8], w5876, w5877);
  FullAdder U1832 (w5877, w5800, IN78[7], w5878, w5879);
  FullAdder U1833 (w5879, w5802, IN79[6], w5880, w5881);
  FullAdder U1834 (w5881, w5804, IN80[5], w5882, w5883);
  FullAdder U1835 (w5883, w5806, IN81[4], w5884, w5885);
  FullAdder U1836 (w5885, w5808, IN82[3], w5886, w5887);
  FullAdder U1837 (w5887, w5810, IN83[2], w5888, w5889);
  FullAdder U1838 (w5889, w5812, IN84[1], w5890, w5891);
  FullAdder U1839 (w5891, w5813, IN85[0], w5892, w5893);
  HalfAdder U1840 (w5816, IN47[39], Out1[47], w5895);
  FullAdder U1841 (w5895, w5818, IN48[38], w5896, w5897);
  FullAdder U1842 (w5897, w5820, IN49[37], w5898, w5899);
  FullAdder U1843 (w5899, w5822, IN50[36], w5900, w5901);
  FullAdder U1844 (w5901, w5824, IN51[35], w5902, w5903);
  FullAdder U1845 (w5903, w5826, IN52[34], w5904, w5905);
  FullAdder U1846 (w5905, w5828, IN53[33], w5906, w5907);
  FullAdder U1847 (w5907, w5830, IN54[32], w5908, w5909);
  FullAdder U1848 (w5909, w5832, IN55[31], w5910, w5911);
  FullAdder U1849 (w5911, w5834, IN56[30], w5912, w5913);
  FullAdder U1850 (w5913, w5836, IN57[29], w5914, w5915);
  FullAdder U1851 (w5915, w5838, IN58[28], w5916, w5917);
  FullAdder U1852 (w5917, w5840, IN59[27], w5918, w5919);
  FullAdder U1853 (w5919, w5842, IN60[26], w5920, w5921);
  FullAdder U1854 (w5921, w5844, IN61[25], w5922, w5923);
  FullAdder U1855 (w5923, w5846, IN62[24], w5924, w5925);
  FullAdder U1856 (w5925, w5848, IN63[23], w5926, w5927);
  FullAdder U1857 (w5927, w5850, IN64[22], w5928, w5929);
  FullAdder U1858 (w5929, w5852, IN65[21], w5930, w5931);
  FullAdder U1859 (w5931, w5854, IN66[20], w5932, w5933);
  FullAdder U1860 (w5933, w5856, IN67[19], w5934, w5935);
  FullAdder U1861 (w5935, w5858, IN68[18], w5936, w5937);
  FullAdder U1862 (w5937, w5860, IN69[17], w5938, w5939);
  FullAdder U1863 (w5939, w5862, IN70[16], w5940, w5941);
  FullAdder U1864 (w5941, w5864, IN71[15], w5942, w5943);
  FullAdder U1865 (w5943, w5866, IN72[14], w5944, w5945);
  FullAdder U1866 (w5945, w5868, IN73[13], w5946, w5947);
  FullAdder U1867 (w5947, w5870, IN74[12], w5948, w5949);
  FullAdder U1868 (w5949, w5872, IN75[11], w5950, w5951);
  FullAdder U1869 (w5951, w5874, IN76[10], w5952, w5953);
  FullAdder U1870 (w5953, w5876, IN77[9], w5954, w5955);
  FullAdder U1871 (w5955, w5878, IN78[8], w5956, w5957);
  FullAdder U1872 (w5957, w5880, IN79[7], w5958, w5959);
  FullAdder U1873 (w5959, w5882, IN80[6], w5960, w5961);
  FullAdder U1874 (w5961, w5884, IN81[5], w5962, w5963);
  FullAdder U1875 (w5963, w5886, IN82[4], w5964, w5965);
  FullAdder U1876 (w5965, w5888, IN83[3], w5966, w5967);
  FullAdder U1877 (w5967, w5890, IN84[2], w5968, w5969);
  FullAdder U1878 (w5969, w5892, IN85[1], w5970, w5971);
  FullAdder U1879 (w5971, w5893, IN86[0], w5972, w5973);
  HalfAdder U1880 (w5896, IN48[39], Out1[48], w5975);
  FullAdder U1881 (w5975, w5898, IN49[38], w5976, w5977);
  FullAdder U1882 (w5977, w5900, IN50[37], w5978, w5979);
  FullAdder U1883 (w5979, w5902, IN51[36], w5980, w5981);
  FullAdder U1884 (w5981, w5904, IN52[35], w5982, w5983);
  FullAdder U1885 (w5983, w5906, IN53[34], w5984, w5985);
  FullAdder U1886 (w5985, w5908, IN54[33], w5986, w5987);
  FullAdder U1887 (w5987, w5910, IN55[32], w5988, w5989);
  FullAdder U1888 (w5989, w5912, IN56[31], w5990, w5991);
  FullAdder U1889 (w5991, w5914, IN57[30], w5992, w5993);
  FullAdder U1890 (w5993, w5916, IN58[29], w5994, w5995);
  FullAdder U1891 (w5995, w5918, IN59[28], w5996, w5997);
  FullAdder U1892 (w5997, w5920, IN60[27], w5998, w5999);
  FullAdder U1893 (w5999, w5922, IN61[26], w6000, w6001);
  FullAdder U1894 (w6001, w5924, IN62[25], w6002, w6003);
  FullAdder U1895 (w6003, w5926, IN63[24], w6004, w6005);
  FullAdder U1896 (w6005, w5928, IN64[23], w6006, w6007);
  FullAdder U1897 (w6007, w5930, IN65[22], w6008, w6009);
  FullAdder U1898 (w6009, w5932, IN66[21], w6010, w6011);
  FullAdder U1899 (w6011, w5934, IN67[20], w6012, w6013);
  FullAdder U1900 (w6013, w5936, IN68[19], w6014, w6015);
  FullAdder U1901 (w6015, w5938, IN69[18], w6016, w6017);
  FullAdder U1902 (w6017, w5940, IN70[17], w6018, w6019);
  FullAdder U1903 (w6019, w5942, IN71[16], w6020, w6021);
  FullAdder U1904 (w6021, w5944, IN72[15], w6022, w6023);
  FullAdder U1905 (w6023, w5946, IN73[14], w6024, w6025);
  FullAdder U1906 (w6025, w5948, IN74[13], w6026, w6027);
  FullAdder U1907 (w6027, w5950, IN75[12], w6028, w6029);
  FullAdder U1908 (w6029, w5952, IN76[11], w6030, w6031);
  FullAdder U1909 (w6031, w5954, IN77[10], w6032, w6033);
  FullAdder U1910 (w6033, w5956, IN78[9], w6034, w6035);
  FullAdder U1911 (w6035, w5958, IN79[8], w6036, w6037);
  FullAdder U1912 (w6037, w5960, IN80[7], w6038, w6039);
  FullAdder U1913 (w6039, w5962, IN81[6], w6040, w6041);
  FullAdder U1914 (w6041, w5964, IN82[5], w6042, w6043);
  FullAdder U1915 (w6043, w5966, IN83[4], w6044, w6045);
  FullAdder U1916 (w6045, w5968, IN84[3], w6046, w6047);
  FullAdder U1917 (w6047, w5970, IN85[2], w6048, w6049);
  FullAdder U1918 (w6049, w5972, IN86[1], w6050, w6051);
  FullAdder U1919 (w6051, w5973, IN87[0], w6052, w6053);
  HalfAdder U1920 (w5976, IN49[39], Out1[49], w6055);
  FullAdder U1921 (w6055, w5978, IN50[38], w6056, w6057);
  FullAdder U1922 (w6057, w5980, IN51[37], w6058, w6059);
  FullAdder U1923 (w6059, w5982, IN52[36], w6060, w6061);
  FullAdder U1924 (w6061, w5984, IN53[35], w6062, w6063);
  FullAdder U1925 (w6063, w5986, IN54[34], w6064, w6065);
  FullAdder U1926 (w6065, w5988, IN55[33], w6066, w6067);
  FullAdder U1927 (w6067, w5990, IN56[32], w6068, w6069);
  FullAdder U1928 (w6069, w5992, IN57[31], w6070, w6071);
  FullAdder U1929 (w6071, w5994, IN58[30], w6072, w6073);
  FullAdder U1930 (w6073, w5996, IN59[29], w6074, w6075);
  FullAdder U1931 (w6075, w5998, IN60[28], w6076, w6077);
  FullAdder U1932 (w6077, w6000, IN61[27], w6078, w6079);
  FullAdder U1933 (w6079, w6002, IN62[26], w6080, w6081);
  FullAdder U1934 (w6081, w6004, IN63[25], w6082, w6083);
  FullAdder U1935 (w6083, w6006, IN64[24], w6084, w6085);
  FullAdder U1936 (w6085, w6008, IN65[23], w6086, w6087);
  FullAdder U1937 (w6087, w6010, IN66[22], w6088, w6089);
  FullAdder U1938 (w6089, w6012, IN67[21], w6090, w6091);
  FullAdder U1939 (w6091, w6014, IN68[20], w6092, w6093);
  FullAdder U1940 (w6093, w6016, IN69[19], w6094, w6095);
  FullAdder U1941 (w6095, w6018, IN70[18], w6096, w6097);
  FullAdder U1942 (w6097, w6020, IN71[17], w6098, w6099);
  FullAdder U1943 (w6099, w6022, IN72[16], w6100, w6101);
  FullAdder U1944 (w6101, w6024, IN73[15], w6102, w6103);
  FullAdder U1945 (w6103, w6026, IN74[14], w6104, w6105);
  FullAdder U1946 (w6105, w6028, IN75[13], w6106, w6107);
  FullAdder U1947 (w6107, w6030, IN76[12], w6108, w6109);
  FullAdder U1948 (w6109, w6032, IN77[11], w6110, w6111);
  FullAdder U1949 (w6111, w6034, IN78[10], w6112, w6113);
  FullAdder U1950 (w6113, w6036, IN79[9], w6114, w6115);
  FullAdder U1951 (w6115, w6038, IN80[8], w6116, w6117);
  FullAdder U1952 (w6117, w6040, IN81[7], w6118, w6119);
  FullAdder U1953 (w6119, w6042, IN82[6], w6120, w6121);
  FullAdder U1954 (w6121, w6044, IN83[5], w6122, w6123);
  FullAdder U1955 (w6123, w6046, IN84[4], w6124, w6125);
  FullAdder U1956 (w6125, w6048, IN85[3], w6126, w6127);
  FullAdder U1957 (w6127, w6050, IN86[2], w6128, w6129);
  FullAdder U1958 (w6129, w6052, IN87[1], w6130, w6131);
  FullAdder U1959 (w6131, w6053, IN88[0], w6132, w6133);
  HalfAdder U1960 (w6056, IN50[39], Out1[50], w6135);
  FullAdder U1961 (w6135, w6058, IN51[38], w6136, w6137);
  FullAdder U1962 (w6137, w6060, IN52[37], w6138, w6139);
  FullAdder U1963 (w6139, w6062, IN53[36], w6140, w6141);
  FullAdder U1964 (w6141, w6064, IN54[35], w6142, w6143);
  FullAdder U1965 (w6143, w6066, IN55[34], w6144, w6145);
  FullAdder U1966 (w6145, w6068, IN56[33], w6146, w6147);
  FullAdder U1967 (w6147, w6070, IN57[32], w6148, w6149);
  FullAdder U1968 (w6149, w6072, IN58[31], w6150, w6151);
  FullAdder U1969 (w6151, w6074, IN59[30], w6152, w6153);
  FullAdder U1970 (w6153, w6076, IN60[29], w6154, w6155);
  FullAdder U1971 (w6155, w6078, IN61[28], w6156, w6157);
  FullAdder U1972 (w6157, w6080, IN62[27], w6158, w6159);
  FullAdder U1973 (w6159, w6082, IN63[26], w6160, w6161);
  FullAdder U1974 (w6161, w6084, IN64[25], w6162, w6163);
  FullAdder U1975 (w6163, w6086, IN65[24], w6164, w6165);
  FullAdder U1976 (w6165, w6088, IN66[23], w6166, w6167);
  FullAdder U1977 (w6167, w6090, IN67[22], w6168, w6169);
  FullAdder U1978 (w6169, w6092, IN68[21], w6170, w6171);
  FullAdder U1979 (w6171, w6094, IN69[20], w6172, w6173);
  FullAdder U1980 (w6173, w6096, IN70[19], w6174, w6175);
  FullAdder U1981 (w6175, w6098, IN71[18], w6176, w6177);
  FullAdder U1982 (w6177, w6100, IN72[17], w6178, w6179);
  FullAdder U1983 (w6179, w6102, IN73[16], w6180, w6181);
  FullAdder U1984 (w6181, w6104, IN74[15], w6182, w6183);
  FullAdder U1985 (w6183, w6106, IN75[14], w6184, w6185);
  FullAdder U1986 (w6185, w6108, IN76[13], w6186, w6187);
  FullAdder U1987 (w6187, w6110, IN77[12], w6188, w6189);
  FullAdder U1988 (w6189, w6112, IN78[11], w6190, w6191);
  FullAdder U1989 (w6191, w6114, IN79[10], w6192, w6193);
  FullAdder U1990 (w6193, w6116, IN80[9], w6194, w6195);
  FullAdder U1991 (w6195, w6118, IN81[8], w6196, w6197);
  FullAdder U1992 (w6197, w6120, IN82[7], w6198, w6199);
  FullAdder U1993 (w6199, w6122, IN83[6], w6200, w6201);
  FullAdder U1994 (w6201, w6124, IN84[5], w6202, w6203);
  FullAdder U1995 (w6203, w6126, IN85[4], w6204, w6205);
  FullAdder U1996 (w6205, w6128, IN86[3], w6206, w6207);
  FullAdder U1997 (w6207, w6130, IN87[2], w6208, w6209);
  FullAdder U1998 (w6209, w6132, IN88[1], w6210, w6211);
  FullAdder U1999 (w6211, w6133, IN89[0], w6212, w6213);
  HalfAdder U2000 (w6136, IN51[39], Out1[51], w6215);
  FullAdder U2001 (w6215, w6138, IN52[38], w6216, w6217);
  FullAdder U2002 (w6217, w6140, IN53[37], w6218, w6219);
  FullAdder U2003 (w6219, w6142, IN54[36], w6220, w6221);
  FullAdder U2004 (w6221, w6144, IN55[35], w6222, w6223);
  FullAdder U2005 (w6223, w6146, IN56[34], w6224, w6225);
  FullAdder U2006 (w6225, w6148, IN57[33], w6226, w6227);
  FullAdder U2007 (w6227, w6150, IN58[32], w6228, w6229);
  FullAdder U2008 (w6229, w6152, IN59[31], w6230, w6231);
  FullAdder U2009 (w6231, w6154, IN60[30], w6232, w6233);
  FullAdder U2010 (w6233, w6156, IN61[29], w6234, w6235);
  FullAdder U2011 (w6235, w6158, IN62[28], w6236, w6237);
  FullAdder U2012 (w6237, w6160, IN63[27], w6238, w6239);
  FullAdder U2013 (w6239, w6162, IN64[26], w6240, w6241);
  FullAdder U2014 (w6241, w6164, IN65[25], w6242, w6243);
  FullAdder U2015 (w6243, w6166, IN66[24], w6244, w6245);
  FullAdder U2016 (w6245, w6168, IN67[23], w6246, w6247);
  FullAdder U2017 (w6247, w6170, IN68[22], w6248, w6249);
  FullAdder U2018 (w6249, w6172, IN69[21], w6250, w6251);
  FullAdder U2019 (w6251, w6174, IN70[20], w6252, w6253);
  FullAdder U2020 (w6253, w6176, IN71[19], w6254, w6255);
  FullAdder U2021 (w6255, w6178, IN72[18], w6256, w6257);
  FullAdder U2022 (w6257, w6180, IN73[17], w6258, w6259);
  FullAdder U2023 (w6259, w6182, IN74[16], w6260, w6261);
  FullAdder U2024 (w6261, w6184, IN75[15], w6262, w6263);
  FullAdder U2025 (w6263, w6186, IN76[14], w6264, w6265);
  FullAdder U2026 (w6265, w6188, IN77[13], w6266, w6267);
  FullAdder U2027 (w6267, w6190, IN78[12], w6268, w6269);
  FullAdder U2028 (w6269, w6192, IN79[11], w6270, w6271);
  FullAdder U2029 (w6271, w6194, IN80[10], w6272, w6273);
  FullAdder U2030 (w6273, w6196, IN81[9], w6274, w6275);
  FullAdder U2031 (w6275, w6198, IN82[8], w6276, w6277);
  FullAdder U2032 (w6277, w6200, IN83[7], w6278, w6279);
  FullAdder U2033 (w6279, w6202, IN84[6], w6280, w6281);
  FullAdder U2034 (w6281, w6204, IN85[5], w6282, w6283);
  FullAdder U2035 (w6283, w6206, IN86[4], w6284, w6285);
  FullAdder U2036 (w6285, w6208, IN87[3], w6286, w6287);
  FullAdder U2037 (w6287, w6210, IN88[2], w6288, w6289);
  FullAdder U2038 (w6289, w6212, IN89[1], w6290, w6291);
  FullAdder U2039 (w6291, w6213, IN90[0], w6292, w6293);
  HalfAdder U2040 (w6216, IN52[39], Out1[52], w6295);
  FullAdder U2041 (w6295, w6218, IN53[38], w6296, w6297);
  FullAdder U2042 (w6297, w6220, IN54[37], w6298, w6299);
  FullAdder U2043 (w6299, w6222, IN55[36], w6300, w6301);
  FullAdder U2044 (w6301, w6224, IN56[35], w6302, w6303);
  FullAdder U2045 (w6303, w6226, IN57[34], w6304, w6305);
  FullAdder U2046 (w6305, w6228, IN58[33], w6306, w6307);
  FullAdder U2047 (w6307, w6230, IN59[32], w6308, w6309);
  FullAdder U2048 (w6309, w6232, IN60[31], w6310, w6311);
  FullAdder U2049 (w6311, w6234, IN61[30], w6312, w6313);
  FullAdder U2050 (w6313, w6236, IN62[29], w6314, w6315);
  FullAdder U2051 (w6315, w6238, IN63[28], w6316, w6317);
  FullAdder U2052 (w6317, w6240, IN64[27], w6318, w6319);
  FullAdder U2053 (w6319, w6242, IN65[26], w6320, w6321);
  FullAdder U2054 (w6321, w6244, IN66[25], w6322, w6323);
  FullAdder U2055 (w6323, w6246, IN67[24], w6324, w6325);
  FullAdder U2056 (w6325, w6248, IN68[23], w6326, w6327);
  FullAdder U2057 (w6327, w6250, IN69[22], w6328, w6329);
  FullAdder U2058 (w6329, w6252, IN70[21], w6330, w6331);
  FullAdder U2059 (w6331, w6254, IN71[20], w6332, w6333);
  FullAdder U2060 (w6333, w6256, IN72[19], w6334, w6335);
  FullAdder U2061 (w6335, w6258, IN73[18], w6336, w6337);
  FullAdder U2062 (w6337, w6260, IN74[17], w6338, w6339);
  FullAdder U2063 (w6339, w6262, IN75[16], w6340, w6341);
  FullAdder U2064 (w6341, w6264, IN76[15], w6342, w6343);
  FullAdder U2065 (w6343, w6266, IN77[14], w6344, w6345);
  FullAdder U2066 (w6345, w6268, IN78[13], w6346, w6347);
  FullAdder U2067 (w6347, w6270, IN79[12], w6348, w6349);
  FullAdder U2068 (w6349, w6272, IN80[11], w6350, w6351);
  FullAdder U2069 (w6351, w6274, IN81[10], w6352, w6353);
  FullAdder U2070 (w6353, w6276, IN82[9], w6354, w6355);
  FullAdder U2071 (w6355, w6278, IN83[8], w6356, w6357);
  FullAdder U2072 (w6357, w6280, IN84[7], w6358, w6359);
  FullAdder U2073 (w6359, w6282, IN85[6], w6360, w6361);
  FullAdder U2074 (w6361, w6284, IN86[5], w6362, w6363);
  FullAdder U2075 (w6363, w6286, IN87[4], w6364, w6365);
  FullAdder U2076 (w6365, w6288, IN88[3], w6366, w6367);
  FullAdder U2077 (w6367, w6290, IN89[2], w6368, w6369);
  FullAdder U2078 (w6369, w6292, IN90[1], w6370, w6371);
  FullAdder U2079 (w6371, w6293, IN91[0], w6372, w6373);
  HalfAdder U2080 (w6296, IN53[39], Out1[53], w6375);
  FullAdder U2081 (w6375, w6298, IN54[38], Out1[54], w6377);
  FullAdder U2082 (w6377, w6300, IN55[37], Out1[55], w6379);
  FullAdder U2083 (w6379, w6302, IN56[36], Out1[56], w6381);
  FullAdder U2084 (w6381, w6304, IN57[35], Out1[57], w6383);
  FullAdder U2085 (w6383, w6306, IN58[34], Out1[58], w6385);
  FullAdder U2086 (w6385, w6308, IN59[33], Out1[59], w6387);
  FullAdder U2087 (w6387, w6310, IN60[32], Out1[60], w6389);
  FullAdder U2088 (w6389, w6312, IN61[31], Out1[61], w6391);
  FullAdder U2089 (w6391, w6314, IN62[30], Out1[62], w6393);
  FullAdder U2090 (w6393, w6316, IN63[29], Out1[63], w6395);
  FullAdder U2091 (w6395, w6318, IN64[28], Out1[64], w6397);
  FullAdder U2092 (w6397, w6320, IN65[27], Out1[65], w6399);
  FullAdder U2093 (w6399, w6322, IN66[26], Out1[66], w6401);
  FullAdder U2094 (w6401, w6324, IN67[25], Out1[67], w6403);
  FullAdder U2095 (w6403, w6326, IN68[24], Out1[68], w6405);
  FullAdder U2096 (w6405, w6328, IN69[23], Out1[69], w6407);
  FullAdder U2097 (w6407, w6330, IN70[22], Out1[70], w6409);
  FullAdder U2098 (w6409, w6332, IN71[21], Out1[71], w6411);
  FullAdder U2099 (w6411, w6334, IN72[20], Out1[72], w6413);
  FullAdder U2100 (w6413, w6336, IN73[19], Out1[73], w6415);
  FullAdder U2101 (w6415, w6338, IN74[18], Out1[74], w6417);
  FullAdder U2102 (w6417, w6340, IN75[17], Out1[75], w6419);
  FullAdder U2103 (w6419, w6342, IN76[16], Out1[76], w6421);
  FullAdder U2104 (w6421, w6344, IN77[15], Out1[77], w6423);
  FullAdder U2105 (w6423, w6346, IN78[14], Out1[78], w6425);
  FullAdder U2106 (w6425, w6348, IN79[13], Out1[79], w6427);
  FullAdder U2107 (w6427, w6350, IN80[12], Out1[80], w6429);
  FullAdder U2108 (w6429, w6352, IN81[11], Out1[81], w6431);
  FullAdder U2109 (w6431, w6354, IN82[10], Out1[82], w6433);
  FullAdder U2110 (w6433, w6356, IN83[9], Out1[83], w6435);
  FullAdder U2111 (w6435, w6358, IN84[8], Out1[84], w6437);
  FullAdder U2112 (w6437, w6360, IN85[7], Out1[85], w6439);
  FullAdder U2113 (w6439, w6362, IN86[6], Out1[86], w6441);
  FullAdder U2114 (w6441, w6364, IN87[5], Out1[87], w6443);
  FullAdder U2115 (w6443, w6366, IN88[4], Out1[88], w6445);
  FullAdder U2116 (w6445, w6368, IN89[3], Out1[89], w6447);
  FullAdder U2117 (w6447, w6370, IN90[2], Out1[90], w6449);
  FullAdder U2118 (w6449, w6372, IN91[1], Out1[91], w6451);
  FullAdder U2119 (w6451, w6373, IN92[0], Out1[92], Out1[93]);
  assign Out1[0] = IN0[0];
  assign Out2[0] = IN41[40];
  assign Out2[1] = IN42[40];
  assign Out2[2] = IN43[40];
  assign Out2[3] = IN44[40];
  assign Out2[4] = IN45[40];
  assign Out2[5] = IN46[40];
  assign Out2[6] = IN47[40];
  assign Out2[7] = IN48[40];
  assign Out2[8] = IN49[40];
  assign Out2[9] = IN50[40];
  assign Out2[10] = IN51[40];
  assign Out2[11] = IN52[40];
  assign Out2[12] = IN53[40];
  assign Out2[13] = IN54[39];
  assign Out2[14] = IN55[38];
  assign Out2[15] = IN56[37];
  assign Out2[16] = IN57[36];
  assign Out2[17] = IN58[35];
  assign Out2[18] = IN59[34];
  assign Out2[19] = IN60[33];
  assign Out2[20] = IN61[32];
  assign Out2[21] = IN62[31];
  assign Out2[22] = IN63[30];
  assign Out2[23] = IN64[29];
  assign Out2[24] = IN65[28];
  assign Out2[25] = IN66[27];
  assign Out2[26] = IN67[26];
  assign Out2[27] = IN68[25];
  assign Out2[28] = IN69[24];
  assign Out2[29] = IN70[23];
  assign Out2[30] = IN71[22];
  assign Out2[31] = IN72[21];
  assign Out2[32] = IN73[20];
  assign Out2[33] = IN74[19];
  assign Out2[34] = IN75[18];
  assign Out2[35] = IN76[17];
  assign Out2[36] = IN77[16];
  assign Out2[37] = IN78[15];
  assign Out2[38] = IN79[14];
  assign Out2[39] = IN80[13];
  assign Out2[40] = IN81[12];
  assign Out2[41] = IN82[11];
  assign Out2[42] = IN83[10];
  assign Out2[43] = IN84[9];
  assign Out2[44] = IN85[8];
  assign Out2[45] = IN86[7];
  assign Out2[46] = IN87[6];
  assign Out2[47] = IN88[5];
  assign Out2[48] = IN89[4];
  assign Out2[49] = IN90[3];
  assign Out2[50] = IN91[2];
  assign Out2[51] = IN92[1];
  assign Out2[52] = IN93[0];

endmodule
module RC_53_53(IN1, IN2, Out);
  input [52:0] IN1;
  input [52:0] IN2;
  output [53:0] Out;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  wire w119;
  wire w121;
  wire w123;
  wire w125;
  wire w127;
  wire w129;
  wire w131;
  wire w133;
  wire w135;
  wire w137;
  wire w139;
  wire w141;
  wire w143;
  wire w145;
  wire w147;
  wire w149;
  wire w151;
  wire w153;
  wire w155;
  wire w157;
  wire w159;
  wire w161;
  wire w163;
  wire w165;
  wire w167;
  wire w169;
  wire w171;
  wire w173;
  wire w175;
  wire w177;
  wire w179;
  wire w181;
  wire w183;
  wire w185;
  wire w187;
  wire w189;
  wire w191;
  wire w193;
  wire w195;
  wire w197;
  wire w199;
  wire w201;
  wire w203;
  wire w205;
  wire w207;
  wire w209;
  HalfAdder U0 (IN1[0], IN2[0], Out[0], w107);
  FullAdder U1 (IN1[1], IN2[1], w107, Out[1], w109);
  FullAdder U2 (IN1[2], IN2[2], w109, Out[2], w111);
  FullAdder U3 (IN1[3], IN2[3], w111, Out[3], w113);
  FullAdder U4 (IN1[4], IN2[4], w113, Out[4], w115);
  FullAdder U5 (IN1[5], IN2[5], w115, Out[5], w117);
  FullAdder U6 (IN1[6], IN2[6], w117, Out[6], w119);
  FullAdder U7 (IN1[7], IN2[7], w119, Out[7], w121);
  FullAdder U8 (IN1[8], IN2[8], w121, Out[8], w123);
  FullAdder U9 (IN1[9], IN2[9], w123, Out[9], w125);
  FullAdder U10 (IN1[10], IN2[10], w125, Out[10], w127);
  FullAdder U11 (IN1[11], IN2[11], w127, Out[11], w129);
  FullAdder U12 (IN1[12], IN2[12], w129, Out[12], w131);
  FullAdder U13 (IN1[13], IN2[13], w131, Out[13], w133);
  FullAdder U14 (IN1[14], IN2[14], w133, Out[14], w135);
  FullAdder U15 (IN1[15], IN2[15], w135, Out[15], w137);
  FullAdder U16 (IN1[16], IN2[16], w137, Out[16], w139);
  FullAdder U17 (IN1[17], IN2[17], w139, Out[17], w141);
  FullAdder U18 (IN1[18], IN2[18], w141, Out[18], w143);
  FullAdder U19 (IN1[19], IN2[19], w143, Out[19], w145);
  FullAdder U20 (IN1[20], IN2[20], w145, Out[20], w147);
  FullAdder U21 (IN1[21], IN2[21], w147, Out[21], w149);
  FullAdder U22 (IN1[22], IN2[22], w149, Out[22], w151);
  FullAdder U23 (IN1[23], IN2[23], w151, Out[23], w153);
  FullAdder U24 (IN1[24], IN2[24], w153, Out[24], w155);
  FullAdder U25 (IN1[25], IN2[25], w155, Out[25], w157);
  FullAdder U26 (IN1[26], IN2[26], w157, Out[26], w159);
  FullAdder U27 (IN1[27], IN2[27], w159, Out[27], w161);
  FullAdder U28 (IN1[28], IN2[28], w161, Out[28], w163);
  FullAdder U29 (IN1[29], IN2[29], w163, Out[29], w165);
  FullAdder U30 (IN1[30], IN2[30], w165, Out[30], w167);
  FullAdder U31 (IN1[31], IN2[31], w167, Out[31], w169);
  FullAdder U32 (IN1[32], IN2[32], w169, Out[32], w171);
  FullAdder U33 (IN1[33], IN2[33], w171, Out[33], w173);
  FullAdder U34 (IN1[34], IN2[34], w173, Out[34], w175);
  FullAdder U35 (IN1[35], IN2[35], w175, Out[35], w177);
  FullAdder U36 (IN1[36], IN2[36], w177, Out[36], w179);
  FullAdder U37 (IN1[37], IN2[37], w179, Out[37], w181);
  FullAdder U38 (IN1[38], IN2[38], w181, Out[38], w183);
  FullAdder U39 (IN1[39], IN2[39], w183, Out[39], w185);
  FullAdder U40 (IN1[40], IN2[40], w185, Out[40], w187);
  FullAdder U41 (IN1[41], IN2[41], w187, Out[41], w189);
  FullAdder U42 (IN1[42], IN2[42], w189, Out[42], w191);
  FullAdder U43 (IN1[43], IN2[43], w191, Out[43], w193);
  FullAdder U44 (IN1[44], IN2[44], w193, Out[44], w195);
  FullAdder U45 (IN1[45], IN2[45], w195, Out[45], w197);
  FullAdder U46 (IN1[46], IN2[46], w197, Out[46], w199);
  FullAdder U47 (IN1[47], IN2[47], w199, Out[47], w201);
  FullAdder U48 (IN1[48], IN2[48], w201, Out[48], w203);
  FullAdder U49 (IN1[49], IN2[49], w203, Out[49], w205);
  FullAdder U50 (IN1[50], IN2[50], w205, Out[50], w207);
  FullAdder U51 (IN1[51], IN2[51], w207, Out[51], w209);
  FullAdder U52 (IN1[52], IN2[52], w209, Out[52], Out[53]);

endmodule
module NR_41_54(IN1, IN2, Out);
  input [40:0] IN1;
  input [53:0] IN2;
  output [94:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [16:0] P16;
  wire [17:0] P17;
  wire [18:0] P18;
  wire [19:0] P19;
  wire [20:0] P20;
  wire [21:0] P21;
  wire [22:0] P22;
  wire [23:0] P23;
  wire [24:0] P24;
  wire [25:0] P25;
  wire [26:0] P26;
  wire [27:0] P27;
  wire [28:0] P28;
  wire [29:0] P29;
  wire [30:0] P30;
  wire [31:0] P31;
  wire [32:0] P32;
  wire [33:0] P33;
  wire [34:0] P34;
  wire [35:0] P35;
  wire [36:0] P36;
  wire [37:0] P37;
  wire [38:0] P38;
  wire [39:0] P39;
  wire [40:0] P40;
  wire [40:0] P41;
  wire [40:0] P42;
  wire [40:0] P43;
  wire [40:0] P44;
  wire [40:0] P45;
  wire [40:0] P46;
  wire [40:0] P47;
  wire [40:0] P48;
  wire [40:0] P49;
  wire [40:0] P50;
  wire [40:0] P51;
  wire [40:0] P52;
  wire [40:0] P53;
  wire [39:0] P54;
  wire [38:0] P55;
  wire [37:0] P56;
  wire [36:0] P57;
  wire [35:0] P58;
  wire [34:0] P59;
  wire [33:0] P60;
  wire [32:0] P61;
  wire [31:0] P62;
  wire [30:0] P63;
  wire [29:0] P64;
  wire [28:0] P65;
  wire [27:0] P66;
  wire [26:0] P67;
  wire [25:0] P68;
  wire [24:0] P69;
  wire [23:0] P70;
  wire [22:0] P71;
  wire [21:0] P72;
  wire [20:0] P73;
  wire [19:0] P74;
  wire [18:0] P75;
  wire [17:0] P76;
  wire [16:0] P77;
  wire [15:0] P78;
  wire [14:0] P79;
  wire [13:0] P80;
  wire [12:0] P81;
  wire [11:0] P82;
  wire [10:0] P83;
  wire [9:0] P84;
  wire [8:0] P85;
  wire [7:0] P86;
  wire [6:0] P87;
  wire [5:0] P88;
  wire [4:0] P89;
  wire [3:0] P90;
  wire [2:0] P91;
  wire [1:0] P92;
  wire [0:0] P93;
  wire [93:0] R1;
  wire [52:0] R2;
  wire [94:0] aOut;
  U_SP_41_54 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93);
  AR S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, R1, R2);
  RC_53_53 S2 (R1[93:41], R2, aOut[94:41]);
  assign aOut[0] = R1[0];
  assign aOut[1] = R1[1];
  assign aOut[2] = R1[2];
  assign aOut[3] = R1[3];
  assign aOut[4] = R1[4];
  assign aOut[5] = R1[5];
  assign aOut[6] = R1[6];
  assign aOut[7] = R1[7];
  assign aOut[8] = R1[8];
  assign aOut[9] = R1[9];
  assign aOut[10] = R1[10];
  assign aOut[11] = R1[11];
  assign aOut[12] = R1[12];
  assign aOut[13] = R1[13];
  assign aOut[14] = R1[14];
  assign aOut[15] = R1[15];
  assign aOut[16] = R1[16];
  assign aOut[17] = R1[17];
  assign aOut[18] = R1[18];
  assign aOut[19] = R1[19];
  assign aOut[20] = R1[20];
  assign aOut[21] = R1[21];
  assign aOut[22] = R1[22];
  assign aOut[23] = R1[23];
  assign aOut[24] = R1[24];
  assign aOut[25] = R1[25];
  assign aOut[26] = R1[26];
  assign aOut[27] = R1[27];
  assign aOut[28] = R1[28];
  assign aOut[29] = R1[29];
  assign aOut[30] = R1[30];
  assign aOut[31] = R1[31];
  assign aOut[32] = R1[32];
  assign aOut[33] = R1[33];
  assign aOut[34] = R1[34];
  assign aOut[35] = R1[35];
  assign aOut[36] = R1[36];
  assign aOut[37] = R1[37];
  assign aOut[38] = R1[38];
  assign aOut[39] = R1[39];
  assign aOut[40] = R1[40];
  assign Out = aOut[94:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/
